PK   T�(Uf��8s:  D    cirkitFile.json�}]o%7��_h^���Yoۻc�fژ^�>؅��lS�jU�v���K�Օ�M~E����[7x�d�d�I2�y��6?�ǧ����������oo~꟦_��ۛ������_���?�|���w����s3<��4<�69O���7�]X��VM;��3V���A؁�|����������������
������������-��:4,��Q�@��p,B%>Vr|�DC8�p��p,��X�C&±�M4�c��h�8��>t�!��
;��>v�!��&>v
|�DC8�؉�p,��X�c'±��N4�c���h�;�Ϗ��O�S�	��>?~������{�����!�7����Ϗ���A�\Om�5�r0J����$ۛV��x��I��]OE���Q���8m��b��g)E#�V4ʘ��g��vуZ��F���Ʈf��1A�c���H�qZv� i}'i}GʎӲcE�;E�;Rv��;hZ�iZߑ����������.`��vS?�f��(޹A�g����S7���oȘP��Һ�Һ���]݋�y;��noi�NʎӲc���w��H�qZv��q"@���������b�QgR��81?�����y-?N�Ͽa"�qn���i&:+��ͺQ��ͰLs3�]�A�q��T�81�ę'N�h�����Rb�Wĉ'άh�qb~�-(����+Z~���K�?�4��'���<��8ߡ��#�b���.x��4z�.t�vlZ�v��àG%G->tgK�8]��ǉ����ux℉����IwVz;)�a�T���A�Y��w����� εq��>�ԋ��fԲmT��M?�a��v��ӂ.
��v5�{+�W�o�~�"���y�l3�vj�le���4�d'��5n�D�qr(��CA��������b�gx��x��Տ:jgx�8��E�rL��ٙ7\(����b��C�>�$�*N|k~��뉓Ð_������m��f�e����6�ȅ4n�2����JA�W
⼒�'��W���8����#��~��8��y%-?�w� p���R��uMt�*����3�T�n�=�������Xc9#�J6�nn�	�n����\8
�/�:��4G]Z$.|�~~i��d��LfA�H��M����Z�>x�;�����dˌ�6�K�D�m�ҠR�v����ۍ;�owX�#�t�-iƩ �B8*��J�O ���"`U�#8$� �>tT2�J��
,� �D�"4,)FRQ���{i�'䝀�=��IȀ9$���J:�k�;ѐ�.�@T��Jک����h�P� �S�=�F��t��	se��r��@�%�x*M]Ya��0W֘+k̕��Lw6����|��sg��̽�Hzl��ό����@��èl7����Iv+�Fe�{o{�#�7��=��x�_�@l�H�`�F>P�a
{�#��� ������>-]6OL�rn�\\���S�0��{��˅�L�j��}P�t烚���<�����5Ow<�9����<�`�����������������̀	k�T_f���G�/8�ho{l�C�/3���#���`��Îz��4{�#�'���H�I���ԟD�O"�'���H�I��$R
�?�ԟB�Oag~H�)��R
�?�ԟB�O#�����H�i��46�@�O#�����MHw?�y��A�ӝj��{P�t�Öu���;����j��:0�`e��]&넵G*/�u��#���:a���d���H�e�NX{l�C�/�u��#���:a���d���H�e�N����_&넵��H�e�NX{��2Y'�=R�����L�	k��_&넵������d���H�e�NX{��2Y'l��_&넵G�/�u��cS��֬3��si��tjm��H�k��R��z�ڻ܇��tjap����g�d��V�j��l�$�j��Q�ć��N��ϭ�5��9�y&�A�g��y����H�gYH��i�	6��X�VvH��*,��H��*,��H��*,��H��*,��H��*,��ظ��_��j��_��j��_��j��_������UX@�/R�
�=R�
�=R�
�=R�
�=R�
�=v��_��j��_��j��_���:#������#������cS��2��a����:@�����01�[�~T.k�K�w�i׳f����g�^P��@���5Ok�<-=P��@���5O��<-;Ps��2Y/�=Rw�����L�k��^&녵G�/����#���za�q��L�k��_&녵G�/�����<��	܄���'���}��#]���>Hm��gG\9���q��fx���+'��\y}h[����ǧ�������{�o������^ĩ���h�'��0"b���aD�| �aD�|��aD�|�aD�|@�aD�|ZEÈ��L��[�?�I���6Y��d��
���/'���ɂ7[t"Nd�p*$��8��pNĩ��Z� �D�Y�Bbka�����nN�Y�BbkQ��Ydq�
���3"Ndq\��q*$�.m!�D�YO!�����q��(P���wߑ��r�����h�����_C�~�q��u��6�n?�F��\y����9*�_kp�U�����l䨄~���W���o�����W^�+�~���Я!W�q�Wv�~-��Я5��Y"�l��F����h<P�+���H#G%�k��
W���NbP'��a�����m���[^��UǷu2�*ly�,�,MXJ߆lI�u�/^'�~@�ʷuR�([�W�$���ª��u����u|['��a��;��m�l�
[^�-��(�o�ddU؆D���u�2^'+��a�.>K�b�N^V�m��\�w6u��we��P�uX�-�o+���F,dK��:y�����:yY��[v��bJ���˪�?�L��e�N^aK��eۯUW���m�WdU��udu|['/��a�.>mN��:yY���ݩ�m��l�	x*'��ˢl���}���.�"Pֵ��қe���>��JwB���e]	>L�Y�8
��`��S����0�m�Z����i�h]�vlZ�v��àG%G톓���(�U�;Q��w�Ȓ^f��ѹ��I5J��iW��"�̸{�Fi˪����H��yiF-[�-c�O�m�ꭝ�h�� ��R|@(��4�~���63o�F�V��H�f��$z޷����P��4�xG�u��.��f���86.�M?r!���`���P�wB)ޑ�\D�3o�Pnd�t��z1�h��W[6�� J�	 ���_\\`���q�.2�7�2��4�v�)�A��R�#J1ցP��x��:N�$F{�(+�4�@)�x<�a{e[�@y���g^�u��z(5g �$��DI��ى�ؗ�%��f�ꊁS�S �r��$v��Q���I��C#�Ԏ�04"N����X)���Ш8��u/��S�J��Ш8�ys/LQŠ���+�$(E���M�R���$(E��Ph�Rz �b̃��H�4�Mֲ�F��#Q���(�<r�`h4\�a04*N���(Ө�<r�`hT\�a04*&�S�셡Q��Q��Q�$�JШXҨXҨXҨXҨXҨXҨXѨXѨXѨX͈iT�hT�hT�hT�hT�hT�iT�iT�iT�iT��;k뢊A_�,��RT��$(E����L�RT�k�$(4z)=J1��TG$^��k0��k0�k0�k0�k0�L��r- C��r- C��r- C��r- 6�Ҩ�\��M%hT\��`hT\��`hT\��`hT\��`hT\��`�f�4*.�`04*.�`04*.�`Y��˵ ��˵ QbG��c- ����8��C�bM�bC�bC�b��8�-���	��MYŐ�ږ;
�R�'�7�IPʱ��i�>*���h	A)�J9ʀTG$^�jH �jH jH jH jH �L�b@	C�b@	C�b@	C�b@	4�ҨPC�M%hT�!�`hT�!�`hT�!�`hT�!�`hT�!�`�f�4*Ԑ@04*Ԑ@04*Ԑ@Y��5$��5$QbG���z��5$LQ�v&fu�`Fը�.M�-�Q\Ϛ-j�s_�L�P��%B)*�R0��_JQ� ��zA(E�Ph�[�L�`h�[�L�`h�[�L�`h\�L�`h4\�L�`hT\�L�`�b0��˕	��˕	��˕�N�q�R4rjE���~�i=��*n�P>u�R<]�RܞB)�.B)�.B)�.B1G�O �������x���?�7~}���W������S������#aDt<���[�FD@l}�H���%aD��X@��q��[�FD@l�TH�c�C"�6]�&�ۜ,pS!�crGÉ,vs��M�Ďi''����8;&�4��b8'�TH옪�p"��,�S!�c�����nN�Y�Bb�Z	'�8.��8;Vqh8��qAǩ��q�'�8.��x
i�������Q�����*\y�n̮���U$���W�ꞡ*~>XE�\y��|���Я5��*\�!�R5*�_kp�U��C�*jTB���ʫpe��UԨ�~���W���ש�Q	�Z�+��/SQ���W^�+;_��F%�k��
W���NbP'��a�����m���R�U'��u/^'��a�߫��m��
[^��?XǷu2�*ly��=g���ª��u����u|['��a��;��m�l�
[^��^Ƿu2�*ly�~@���ʪ��u���u^,��˪��u��uu|['/��a�ח��m�7b�^����D��L��˪��u���>u|['/��a��-��m���
[^��_UǷu�*ly�~Y���˪��u���pu|['/��a�����m���
[c��uTc�:��V	ݨ��fPm���h��]r_�N��Z�7�e������7�w]���5�`�y��q2�ͦ;Qh�$V��m�M�I17\��QF�Cj�8g}'�2���R���*��d=Z�G��ֶ]��0�Q�Q����Bå�]Jbe�ʬ�0:�6�0�F	>9��Y��wO�(m�/ ��_�1/ͨe랣el�i�S���-�@APh��h��<��mf�N���tϑ0�<�I��ox�R~�!(�;��լu�m6C�Ʊ��m��i�;���R�#J���"��yÅr#K���׋iF3�Z��2@����R�#��h�����ͰLs3�]�A�qЀQ�R�#
�c�������M�TC�9�7�7��I��4�����v!(4~I�gډ�؁�%�gh'Jb��N�ľ��(��4{UG$^���|�ojc�^��/�pj��^����!��4*N�Q�C���Nн04*N�|�}��(JQ5 ��h`�'A)J�%`��`@(4z)=J1��TG$^��Gn�~�#7�F��C������Qqy���`�Gn���#7�F�D#w�p��04*�4*�4*�DS	KKKKKK++++�1������������5��5��5��5��5QbG�bM�b]T1蛣EـP���E��8	JQ2�oB��K1�P�1�:"�Ҩ�\����\���(�\���h�\��Ш�\���`�k0�k0�k0�k�Q�F��Z �h*A��r- C��r- C��r- C��r- C��r- C4#�Qq� ��Qq� ��Qq� �:hT\��`hT\��`�;�k0kk���!_�-w��O�r7��=N�R�$зwIPʁ�R�3�r�����HuD�Q/�����/����Q0�����0����Q1���!��4*Ԑ@04*Ԑ@04*Ԑ@04*Ԑ@�.��5$�T�Fŀ�Fŀ�Fŀ�Fŀ�Fŀ�hFL�b@	C�b@	C�b@	�uШPC�ШPC�%v4*Ԑ@04*Ԑ@0E�e��խ�U�:�4}��Fq=k���΀=� ���A(E	�P�
�B)��R�/��^JQ� �+0��+0��+0�+0�+0�+0�L��reC��reC��re��z����Z�(c���k�Ej��أ
B)��R>�	�R��(JQ1 ��`@(�z�����ߟ��ǧ�����R���r�49|�ԏ�t�8<>M��͇~�^v�V|n:��ԍ1]�(�OM�U�t�C�t7t�낏��_�#�,SWf��Բ�o�m���\[�7��m3.��R*5
��g�al�_Y�����_��G�\_�	��&��Ɂ*IE��x��J�
�</S-�4AG�A
�A�C�pT`ax���W���0X�Ns�[��,���h�{��th��Vnky��l{)��PT$E�$kac:�	L(�y����;1Gr�:�Ҙ����1���nQ��LJG�1w-D���3��O?�ʘ�'��Zs��7��s�ǁ�#.��5�D_��c<T��+'�(� jD,K�Q�y��K'c�c��,*#@]:Y� ���tR���qs[�<x�0�
,%���x�C*�hg��!zh���Y��9u�U���R��32DUw��x0�N����R�஖赁3Rԥ>pJ��]Rݷ�r����vT�=�	2&�j���Q�B��D��s	|_��r"����\9�pߋb:� ::�Klя
����H��˾w���O/���6O��a�����qv������xȗ�Y��=� ���J��E�n�O"$z?���>����X�@�	���#�.+���6d���<#�eya��j<#�EYF��ψz	D�ѻ�����=Dd�Ǻ<!������$���K��f� �t� ��� ��?!Ů��2��*���+���"
ص����?�#W^�	 `�	`�a�?�r|n�]���\��3�yv�F>(��R<#�xF؅x���%F�Y5��I�w�}�!M ;��	����o3��|�@�c�mR-4tf�Nx���&:@�����$� �Q(�ތ��y�(��S@'��~�&����M���=�C!��
�ƀ�@j�l��ē ]��'�X|]������	Q�a)�e�&���׭0"^�^o�t{��_����b�X�N� ��=>�e�O.���:(��Y�{ �}�خ55�# O�xc �v ~Bn�@��@n�� �w S������s���.x�8���%NeK��2s�3��9Ge��;b�?����Ǽ�� \B�������?<�<���͇��~\���Ϗ����͇_߮=<��4<:[ص�zR���^��`�I�Hh��Ԋd��`�I�Hh���d��`�I�Hh��T�d��`�I�Hh��q�d��`��Hhv<c�(�'E�$��� ��1��3X1�Q<;~� ˃ �r�@��`�O%`y�RNL����,�x*�)�?��A1����SAO����,�x*�)�����AOA<�c���H�<� ��!�޺�V^(�|��T�>ܰ�OG�l���'�.'�n�os�i�j/PE:�-���+��Kˏ�c�A�x$����7B߯"��"�-��e�~5��4��h�qb~l����������*FK��/�!q�%v'-�`iP�=�7V����%v'-?N̏:b�u����ǉ���;��:�!fȩ���>$�`hrj������b���!�����0`��� �Jf�i\J��3��� =@��pꌆ�!�f���Q��:�!fȩ�w��>�Ne�rj���<BR�/��#�j0*_����]J��3������45o꤆�axVi Kd�b{^,ޥ�9N�p��i���4�l{j1���oj��ZXK�O�"A�3������4>�΀���u:G��e���x�Rg@!Í�y:1aBO
H���{K�O�R��HP�G�95Cv�R�G��T:G��u~������Q�p��Ķm��D�"�x����:�_��>�!�z}�A8\���a+���с��p�����?7B�}x'�}��zg{Y(��<�/�Y	eL���7\��XR~&��>�0yw�
�s՝p�羋��L��N���N��ݥNŀ}:^�M:�E�|2��h��;��G(&�x8/�}$%�D�`5s�;��E8ԡ=)���	�$� ��;\b�����;\��eg�`W����n���] {����0�\�B��y�/�H��<��N��x�N�� X��{Q�`e����'4)��ae����i�Sq��\H �0�M}o l��j����TU��'�}��YR�'>�9&�}F����g4 j�� �}F����c�?�@�3a	�� �
�����`x�^ �
s$ ��� 	�*1<�`/ :b��a X%�FD V��1ܟ� �D�U��*Q��e�%V��D�U��*Qb�(�JTX%*�V�
=C�*Qa���JTX%*�V��D�U��*Qc����
V��D�Q"���gT j��}F��	�>��l� �=��3��>�`�A��\�
�j0��� �*��0 �s�* ��\�
@�B�s�* ��\�
�*1��� �J�嫰1��\�
@�X%��U V��|�Ub._�`���Wa X%��U z��Ub._�`���Wa X%��U�<��\�
�*1��� ��
V�k��Y��X��x"t�,�S�թ���`uj"kB�0����\��aUlr*n����4\wc�Z-��3����Y�)���u�������H�\���u �=�����>7�A���}.F�� V�ٚ ��l��Ua����0[� `���y� б��l��Ub���*1[� `���y��4��5 zX�*1[� `���y� �J��<@ X%fk  ��5 z��Ub���*1[� `���y���X%fk  ��5 :Y�*1���Ub���(�.�Ĭn��\�m����(�g�5۹�e̠���gdj�Q!�}F�����g$j�Q �}F���X��2f V�����`.c�`U�˘a X�2f V������X%�2f V����Ub.c~�=�y��p���ϻ�n��߀��o�����R{�ApG��v{���~:<?�����@�����Í�@~���rd�[���AN���
䬗˫��H�r�� ��9?$h9�#h9�"h9"�=�.հ����?/S�6ֿ��o�|@ZO�YτY��Y��Y7���Yח��ۼ����H�F��!_���Z�[���B(�����-�o!}�[ȕ�o!}��4���[H�B�ʷP���-�z���-�o�|�[(�B�ڷо��-�zӾ��-��@����v`ʁ�|�[���Ʒ0���-�^H����eG;WBfW�W�!0<��~tC����0?�����w����F&	����&��Cv�u�yx�m��$���±kK��v�����lCvm��6;Qb�a�a{Vz��;�I~8v��;�1찾�%߉;ࡎ8v��N�|;��n�咀�LEc�Ix8v��;������p�J�,K=��C���<��Pg���Z9�I��T\Ժ��Mj܄�:�����I���5�׳���'�f�3fK�X*x�~F�+�wD�s��$1EАL�S�s(1%ԐL2��b�)��d��V�����Iͤ�������K2�����A.6��Dty*%���S�T:|e����"Sjf|cCEn��oE����χO�0򵋍�����������'��2/?��'��j_~jß������ſ�i�m~��x��8�&����7�&O�-�������?��<A��� y�O��3�ə<��ӭ�w�Nw޸xm6�f"��$!jH��\�w.N�'��c����r<�?Ɉ�:��q�➍�ӧ��4������������g�++̢̲���5�m�Fl�܎�ꙛ���?}�����O��싇�gU�ז��S��?���_��Śۚ�|a_�W�쫺���������|?��/������[��_������������z{���W�_v}R�>�;�7�߾���˟��ü��������/��_����׿=������<�|xv�������ҏ�_�������X���_���?�������<+G������?-��Z�JSߺ1S�qiO�n��'�G�p3L�sI��t�w#�4��k�ǖ�˴�����×��a<��8��yt7����ݼHu�?�/���Q��1��}���y�:�X�򧏫��?����t���������;�8ae��C�yg��@��?��w_�!,������V0}'5�:W���]�qO�"����~�a�-��c�n� Z�U���_
� �pR�W����wa������eĬ�n�]�{��d�E<�̅i?�	���޹ ��)��sMjZv^��k��O�]��r��?z�B@�5[}���3y�$���.'�\PԎ�aq��iח��zq�-n�y|N�mc����$�U#�n��=��ajY��}3φ��E��5�Հ�mU3=��覑zՍ�*��돚D1�Kp?,s��N�nz��)���:w���0�m�{$\�u�yЭr�Y.�f�X�`�VQA,ޮ>j��,�Y�'�n�R�nu۝S�m�i��J�Ј�"�}kF�D$������H7x9�4��j��̹
�Z7����ŏz�����/����9�`��8��hK�&.����.^w��_�TQ���>.b�x����M%��tbh��#�m?w��
 K�@Aݍ7�)B{����"���|��?���1�'��/kn��Nln�r�ҥ�&>σe���ﮤn�tr�N:��[�����R��Γ�[#�{:��r/o��߯�s�r����ir&/��e�:3;�Vy��?����L~������{-�FƬ��d�T@i�<�(�N�vI���E�e����m�n���S׏.O��8+��m�Vl�o�Ɍˣ\߬�;�߂��32ō�����dǏ�Oe��o��]m~�j9�����	�p?8�\,�9=Ri�e��ě�s:��h]�ss�Q��=彜� @��B������k�:f�5D
�R�8���h���_b�5��}[�^|	�d�~�I�~��7�5+�<l}�r��pLk/��.R-fqs��,n��h�/w��0u�Л I�����Jl*v��^&�̜��ް�/�2eh�����vܮ=J�e�[���y<7"�vn��"蔡\��d��ur�ҝ�q�۩�g�vv�sy��Nv+���hv�kq�c/.lSvr����'��'��O�|���!�����%n�9nt[�,PA�,TU�.�i�.�}�,|��f�C7�]5B�ꃉ���K���Z���q���m����Y����y��g�|�4vn����t���:!G���i;��6�@F�5@�6*$������o/)�Z	> �N���-��`���I��.�wN��s�KF��/q��g����SyK�Lp�Ydd�{a�RW��/1t]s�V ���(b��7�X���l�H��O��т�C��݆v�[����8�p���$�vq��]�a�0��8��Ĺ�0��3�#�q���eG/�&E1b�1L��Y�Y�s�m���]�ch��1�2�]�*��x�O��4���-{5��J�.z+�����b���v��]�ah�`1�3�ǩ1�y9D��C�Èa����?bg�%F���Vda�����v	�Ðᷘ�������ŔF�v��\TUZ�MK'n���\O�b���vjЪW���A{�!�_?#��G����iҳZ��٘��9b�^n	u��5�MY�Ӡ�J_F8͋�i�.]�ǅźS�ǼUض�yL]�1i�c�*��ΐ�<����,?Z�H&/5� ��9!j�k�0�UQ�X�Gc���45��{�"��Dc�c��½gRv�ܱ=F{��{�V�L��K)�uǿ�p;޾Ŀ��!��]苨]̹q�Hw��{>nQ�0"˸aD�q�ȣ5�=�q���7<�q�HЉ�����d�@�V��w�$⃄eĭq�XO%,#�����)a�h��\�	�ȣ���<�qK͍�#m�W��;&uk͋�=�7򫙎�䤡��8G�V�דw�B浒�2�흰Zꓟ���O��U����g���͕�_��V�^�6�u��HZJ�A�z�� ]�
��&~Y�=�2�3��?O� /��s�]�&���
=L�if������4����Q/.��<\-:^(�����P�}��|���[���\M��ƶ+��]<O؄(���p��b���~Y,ࢽ��/�8�$������.�0�KQ4���d�e3�7�8��,EOY��.�Ֆ�f)z���͘�Z�E`�̸!w����/���E`��@�"0K�:9�K�  ��������.Y� ��R�,�{�]��R����i���\��H/0K�S@�v��ҙ�����"0K݅ :9��յ�w���"0��~)��q�U�Y�o�Tw���i���� e�n�bh&6-���5�hyc���R���*n�1�в���:�ʽs��4.�|��34wF*����e�vy�KwX{�ʼ���)�v�~�����`ޚ�S��܈�<�U)��u�:�Z��.^77��=U���T�2	���92��gc���w�]�t�.�'[�����Lw�����Y$7��f�L;�a���Zu'�<�h=�AТ�Ӛ�嵫��Ɖ���^q71��IZ0}ǙKl^Kqq;�WA�1)�Pk	�@k	�Pl	C�g-��;q^��0�vo�N��3���w��B�3C}':�FlR��|)0���s�۝ӆQZe��k�*ݱ4�w�4�ՈčH��e��^� P�κ�ht��j�\�c����.���$����v��Ǻ�i��o���Ã���`��xT�F���W�����0�`�ݺ����5����L)O�ŭ�.ص����{��%H#\������z�]�w'����s{|~��s�����r]y'����F0��츋i�Q�����qϟ{�;�O����6<~}������g�Kӱ��ԯ;���Z��Z�躿�r?=��_�]���~�W���΢{m��m�\^��8ߏ?��^O���i~~��_��_���Ӽn���G'�O�O?�|���_�q�Ǜ�o�P�������t���+��0E���ܮ�O�/������"�Ϗ�����?�����7�(�?-�������~������[��=G���m̪�Z�M�@+-����o?����v)��['������!����҉��+��-i9�l���:a�&���[�V����ڲ��pW�/M+�����+�#twʰ�37�u��ʊxl�YU�`���i�c��`;�RJ'Bw�t:��֪�Ɠ�_F0��U���]a�`�d;�V��J��J)�ݝ2\�98�I���̥�QY�+���3�iţ��vp�O��n�\̻��R@4�1��I����������/)�j�_�vp��X��^�]�X�ܶfV��G"f��̬��L\��AVU��դ�+���ZI�׆��3��R�4Kj�¤�1���t6���VaT�
;w	�%Z��+��+�`#t�
�]δ���Q�n�.�ο�]aUE=�/ݐ��_[����P=1�{�#ԥzD��;n�v�^cVe���~�3�\)���{�ԗ�H|��4�,j&�V�L�h����`���ص����#H?�N�=y:@L_
�҈�;���ko^X��fuy,���.&_@+7Y�Z]�V��9L�Y�{-�7�2���I��vpKj�*z;%{vzӪ��*0����dv�w���^���s�U(�Ԇ�GO�G�@R�}�.�=� R�Ao��.�K��J�Kuv.���v�Ձ�E2�S�y��䇌]\JnDQ'�������!��NJ�{�X^J[��D.�1���W�C)v�9]�(K)%������#��Law��Rz݂(�]��������V����p�]T"f����I\H�қe&R�Z��#��B*Tg������ق@�v�����1�f]tjv�=�=fPY�{e
�<+i�j�}c
�J��F�����7U$2ÍU�
�s���}��T	;��GH�`c��Y�����^�VP&�������=xv����A���c������g�ՍY�m��l�S��K�ּ�
�ܝ�f��6fo;X�,5"�'�R��N��X��T�꺂���:�ȭY�c��Of�����D��K�h��2+��u?L�ȷ-/�De�Y�A5�"5�"5�"�u�|=q>�ȍYJj��o���(\J��P3���Kl�.�jE�R����*�n<�"�"�E��v�ڗ5�䨽�c_y�+�����lT�R�c(5�Kv�Ҏz�jT�����
����,5�Ӱ�ߥ���?V�;�cU�2;��z�ȷ-�3�Z��i4^�<lW��<��;<ّxc�Yb�e�
����!����v`��ZG<WV7�>��x3R���u"���]��T)�I�㕱ד�w�%*h�`>�Ch�k��ZG;W�Y'kގ�Ȋh�X��Nb��b�������������惗ӗ�?���<�{����ǟ��<�������n~��PK   T�(U��c#��. ��. /   images/46b9f12b-d0df-46aa-ac71-73c8a35b8753.png4�{<����6�d�6�e�i�b��6jl(ws�Hh�I�~+���\s��+*s��%��B�$D!կ����������z?_��N�ěr��@  ��5" �  �㿞�{� � gd`Map\2�p6����^F3z���yN,����S�Kb܊ґ���l�t+�2�S��>�������NƢp�����ޑد���[���~.�����]�㕨�?��z���/=
=ݬx<k���ϯ������w��e���tG�l�;A�����'��y�����c�~�;"]�N��9��|Y��C�;�N��?��w�������������_�:\_}m]Ը��2���}���?�t��r
�3�Mޜo\�sO�ݪ,��<9�>���=��@E�������}D��K����ⓒ;S�����\pg�3�����9ˢ�D�_��>7�yE�q���W{]l�+��L�����WV�������X�er����V�Q�$֏�U�X�A��T���;���	�b����ʅ��;�`�d���ɗU�\�U��j�1%�{�Rbx�)��l�QS���4[4�7]�\c��(&�ӎOB׌�ƻ�	�d֋� �|o)������������,ϪQ�~�����Om��0p;�����N�Sʥ��G�N��aR�]����V������fM�ݢ�j�&����}�]�xF�8~T%�XV�΋7{�~�'���#\�ۏI�)�<	��lI������1�X��wK7s(��uq�2�q�4	�yw���(���w�%р=uf>��r��<V"_�x��Dw77	nyNà��<$�wx��������b\�=$�Ms6 0g�S_��t���On ���sa�J��<(w���` [�V}O��U�K�������M����	�eQ��L�r=$f�k{����Ԟc����X�#�����,��C���{����q�g$������7��nѓ8�=�7�}��'�<,1�@�L}9�����"@��+���N#A�E[�%��l��9��%�TE�
'V�z��4�`�ZhW�w"]5v����Gf�&n�{H�2E�m�����3�f�Kb��G��V����{���Ŷ�+�d��7=^�P�SK����t����X�K���|�_l�SbU̜��L���wR�r�6��8��'�}���ɦ����{��b�<j�}9��MV<ù�l��!GW_�+%˚���V�@��U�u�"�8�����0S��|�b�.z�ܐx4��:c�_�!W�T�;u��iޤ,��%"��n��kF��%���q�Y����]S�g߫m�ԣ�.B��k���!o�;R���b,���ئ��Y�[W��S�Ě��8.��cL�LdKƈ֒�%J/ ��A�5��Y��0C�?��#��F�d0;�ק��Ě!���ܹi)F�Ke�r~�O]��c�1���	b���Ng�y�@v��tr T��ь���O���z�����Y13<V�_㥷�v쎀�Ht쓪f�J��jix^�m�������΃Pm3�/�{:w�hN�e,l����@
U@�+1��C�}p)����K�&��1��������u��Z�>�{)9Ev�pT�z�u�������9)�
��>}�f�:�<�f�j=y=A$J ^�W��0u���B~�ү>a�����~(5m`�����VǠ�
�HZ*L�0j�C���E�v{��԰�����	��{P/T"�E�s�F\���N7�&��.*���x�@?��Ċ��3x��+R�����X���Ő�׭�j!��jr2V���#�R�vp�Ch�Yh}�����1�4���S^���˧���k���B�n�1`�9�c��RWM�co��܂ʕ�W&Y���d�_z���۲�˦	M�,9?|�Aӎl����ފAGA���|��������D��w�g��q�ѱ��û-N�u�����6�t�e��M��mvU�5�\<rQ(��3�M�̂�5�D��g;'.�n���5��jm�q�DL�씤���^�����rP����_ƴ�_��L�8"	�kg{]Ԅ�z��=.=hSS@�{��#Y��*ږ����/߮k?Wx|����N���U|zgk�g�f��j���ݶ�e�kG��ޘ#q]Y&|�x�w�v�@�|�>�G ����p��!�,';f���$f���+��z4�g6��Ԍ/��@~Roo]����]��D���n�D�����@2��r�Ӌa�v��ma?�OF�~��n?ӹ�v�����H
�+ ?V���.�Ͱ�����bw��Ӎ{����罱9����Y���a��%�R���`g���T�cS-�@?�r��@y+q[��%,�ex��}(t�n�3e���r��ܦ��V���4�P}��2�Ъ|�8�ms�!���P_�K��� '/�}{\6vM����b�������5@3�o�)cIG�s�-&[j���.B�k���5��5BI��#�Cb:FL����Pv�F���D&fxΈ����Jd��d^������F��z"9;�;��Y-:"a��WѺnXҜ,e����\��]Ai&���\���=τ+�CI�:��$�\R�ώ�	)�d=����Yq�L9Pz8j����.�kly�:{�^����t���?w��N���ܬJ|�!a��ژ�B%%^��&۩�vV� @���<W�5~T����Z�Kv=��ѐ³��3!�a9�<'���܏qi��_2�\=�aD�+*m|$���?�ڮ��b������<�j� �{���I7��ByٵT��.��Y��.��	Y�q+2H~�����s���^N�PwNK!���mѰ�"�+�ǹ��[����x8��e�	K�R�ڛ�Lb�� E�i��2�@��W�E|vb�pi;k�����ˍ�����{�m���7���dOrk��ӝ'�fؠΕ���M��ԍ�6�]�V
�SC���_�4y.4��+o�fd�>�7��7�Bj�L�����&�# SY{Z��w�e
�2�>@$}*���U|i���/��˜�ޡm_jύ�r{���p�����59�i����`����E"#��Q�>�]ޱ^w�٫:�8�^�t�ͬ��!��b��f8rԽ��-*�02���u���DB������M��� E�k۵qݟ"`TUj��\�[��+��7V@��F��R��m�mᝅ6@�hI�����/�@о���[5ϴ��y�,O�E�O/L(	�m���=v fJZ��\����<}��2�MT6mZ�����IF�����vǃ������k�[�ż3d���*5E��*��.}K]�=�nT�(���c�����|���S��XV8��v	,F�OjD�R��U����+
��&��AC+��f��N�W:c�w��&�2��\�];z��9�a���S��!���<�x|^�� K3����X���H�j��RP�nA�Յr֎?����2+g�4������y�I�i�Wv��������Oϭp߬��(�$�v��"��B�%��J��@)F�g$v2��E�Ø�U*rY�,�Xm�zR�4�������=uvƨ���(��L�
�m(�p�α ������~��T�v\��-mi�Dg�Ǵ�"�H�[�K�٫��"��.	��C"S�e��t0;W���A�R�s	���'��n�_{�G���T�"�ω�,�v�8{�Q����őt01䙚F������P����_q�fJAR�F�	H���}�-g�R#���\{D��g�l;���y��mm���Ƨ��Ӻ��f>��{j���SY<���n�&'[���U�kȀV}�5�i�V�
�BP��j�{)��G�Z�SB
u`;�JkF��c ZB�)�V۽f��\�&�v�4�}O�Gxj�����{�><����8y , TC��64ƻ�ߧ1a2���d�����G�NT;��L:0f�&EF}U0C����ܕ���[EH@1�*>{y���
o��nT�L�k�cY���dN�* �B�+Ŷ��4�c����]�NУ��b	��(LS-�g�_�e �w	[�
�d2"J+����ʡ��i-��d����=n?x9N����p�xt�]�%+'�
y�6	��
�_��^��F�~hc�k�W5�3��:�)}�J��M/;T����D���.�u�*�Rf_�\�3��O�x���[)c%�]�Z>�ؿ'&7���B	n5f.�!��v�B�U�,f���+���:���S�h$�*���B�;�Pǜ�7�z��ݕ�`D��Н+��3����q��@w���z�*_*a���7i?�A�EV{��mNrߞ^�׹�����눫q��6��$���5h3g��7C���Vq&>,B�ja1W����p�l�KiT�?�h��I�8�:g� [���GB=9MDO���(0A���U�&�0�C)�+�i{D1g�����Ey�F��g�y���ͰStR��-=���b�-�qS�!O�����^i�3��I�N���KĹ�>������@bA#"�~Udܯ �x�j��UTu*6n�K}~�~_.~��J^-�]�ֽrI�]zj�YLŔu��b9H8e�v���>�q�L�^����Ԑ��ǁ�w��&�/�HtD0���)Hz/,l˖�m~�a���x�i�XV;�R�]�MT;�l������?X4y\ ���R�n5<�0o�D��8�"
�ى�^�	���~ľ�N��P����qx�Ֆ�)YK��
�W<�+�O�:��u�"�0�a�����~��w23��\-�y܊U_\�s�hH���j�$�{V�'��q�m�l�K���7�����p3>y/]<�����B~r���KS��Yb�2���555DJ��������!����r�n�"d��N�o��j��	�La���[q~��Cˇ�/l}��l��Ʀ���=�oX�51�\�|՚WY>���j�;kM�Y��5R�#�R�3Cq�����#Awd�`m��HA�4��P@�����Q_??N��i��-t�x�QW����ƙ���:����ӜX�-$�k=�zw���>.r%���}�+�
�ց��M��%~��^�(���<��r�`k�/Q��0Y3c����s{wӴ���<]~axZ^!}�L��R��{ŷ;����v���K���.�[WH��*޸n�a�lg��rI�����ݵoU�\������HXM�/6����3����ސj��T��`~�U6-%Ǩś_=���#�׋k��c�_hP"<Mk��tۅ�Vư�����9�2H��0�p0K��y	�ʟ�����.f��A=���3m��ZѣTe�V/��g�N����8��|W�H���)���3ķ�D��v�,4�b9vfCɺnu�W����!6�l��#��h��ƣ�Ѹ�oc�(��-�o�
�NS1��
������YU�J�R�W�ĒI��,��W��[�DlT->��S�L,|H�U�p�'I[Y��=�Z�~S18���bL��9ߖM���KD^�ߢ�܌1\C2�7�:%=f%m�v�g���l��+�gh�Յ�)�{W��FT��͘W�N��6ܡa�^i��9�0=yKR�Ѩ�S�w������|g��+�c�vY�|h����3�sԛܝ��..���JU�2��L��V��@�j�����hp���������t;��h��z��ōR��[�����`?��o �j����/O������$C�&�e@�ܪi�Н�m����f�2��9�;�o;�%�<O�
�m�n^���i�>u��y{��fK�V}�&n��}��.�p����Ku$`�u�݊=��0���t�w�@�@_�y����st����Y�Ȧ��@DW��)_�����{�K^ٞ�����%ƕ̧�)W%���?8,�^-�}�U����	{Νrc�/�(WH*ی����ϼcd%B�u�)|<�)��3v��K���� O\zSD�Di�8���Lu٪�ܹ�noP�h��������ddY�2Ug����� �h[�^jG��/���)�\�|~\����{%q'��Es��tF�ɪ�������g����^Ro��3b�����ɦV�X$s�k��rX��������C����i�0ӄ�(��)��J��
�n� 2��J�t:b_��g��v����!/iA�ӯ�;�P���ew�
2�� ��m����G�h�����������K�C"̍���E����`��h�-��us�zw>���Α;auF`��a��`q�@9���e��B���O2q4��/�9A�m0g��w����Aq(�.�n��p����Yk�CMƑ�k�°��u���k�0���2���_�2}�A�;��Q�ÄmY;�[Ǌ��kQ;aY�b�x�|t{�~"~��" ,��уC3�I8B�E)=�E����JZ&�1��"�o.��-�;V�"��c5�V܇%`��J(�|��J�F
�tU�F܍�f�u� @�3�b�֊j?�7O��(s���ɩt�$�r��.Oꮭ�VVW�rv
P�����#��,s����>r�gM���K��^}V�?��Gό��L�]�!	UM!8����;��#�0�Ո��!�����>*nj�
_�����b��S�F����Ό�;_�����;�;E�v���4�^����@��V=o' ��B.��G�ӳ	�b'9K�}ic�NK�bek'r����bM�����[~�d{���@�9�E~@xs����('<8S��s�R�-�'�������.;���`Xo\K���'9��D�J(V���úF�ɚ6�v�d+@_Y՜{����˚'�$]�>��1�=}{������i �2N�R�o�34Ax��@�� �Ry�
-5�����z��
����D#$����y���:�M)]�܌4�`hϬB:ň�����<��`�+��cחr,�D8P[1�["j݇N�P��J�{���q��S��C��\Ƿ'j�O�끫�S�7���7�lo��5y�q=�2��_�>��h3���ύAF�K�[�޲��G:��>�ECW{& �>���E���RS8�� �3�v��qKl�B�)�hݻ�6���"]{*�T�����U�g�<��y�S���ޏ�}$Ӎ��Àzp�zq�
S����(�R��)#��GD#@L��c�giM���?#f*{T�*nu���-��s�a�A�՟����X�,Gd���#NJÜR��$��Km3��}��AD3�#z�+R�8�������U���j����\�~�w��.�;%�m�2`�mC��J�B�����B���s�9C=��iI�،�m`c5PR\����tf�G����p�ѐ`	�2��u�W���f��f���A��U����[�Y*�;aR,��8��!&�8K��6]�\�Y�,v���SIH��ii4�cF,���%�[��7�b4�~���yb����g�߼g�����T�f��De-��H��Z�|�*C��gC��8i[5Tu/�F��:��^Si���a��h�V����l��^s堋�E@Q�H���}m :F��ݴb�)��{��),ڡ�!d��0�p�36����5ZB�^oL�|솾����*+g�����`(v5�;�5�#`a�w�
cR:o�\��"�(ճ@�~<І��@E_���T�ԅ�5���l�R�E`�;!k�g2BH�UT����b�X���>|�������DLKe[�LIM*���n+=���(�J~���+��OE-������,-D�py�}����e�\1��Iȟ��mx�y�ћ7މA;��Q���V7���Vg��U@a�j</.䢔���HA���Vս��ޏ3�oV2�l]\�}OW��+en,7o2�4�p_G��P+�f5�s��\Z�����t��Md��l@=Z�Y�b���,��<��a���@|��UETԝ$ѕ���HG�
JD�L5L�C�������|F=[)�H��S�<�XL �_t2@�p���'�{�:�!?�-!Xb���<�v:і�����@,���I&t��PDo$���ko��4-�Ũ&�H�޻ȏ��EI����}	B1�O�t�u�`sZK
_��tnX�%�e�k�z��Dd�oܸqF���P]ͽ���an�C�uX�_}W'����5�o��}�C�>Q����A�S�e�-���)��_0�3{��;==��@1��K���J�Gl�<�95\�c^V_��m����?(dD��<����|���j]]����ly�p͘���R���`����{j�j��^E�xVN|��济[��Ї�w=���)j˿��H�{8�~|it��Mq�4M<�H\�s�-�vҞ���:?��� �u٦�
{3�l�c1A�2&Z+8�S�Q�=Ql�xQ ��RX6��V�ȭ�'	����k���rf�D�T��?��������!3��z�׳��[/﷭Z\pn�?�����G����ɏ�O�Sn\ƥ�&Q;mn]V����=2���e��gQ&1q�J۸/K�u$o���:������G|�z.�%��;�2*��m����
�Z~�ҷ����Vj�3OH{�A�rvOok��Z�El�����owiff���evY=��Yr[��\%��L�7{��Rڭ�Nۋ� �$3��9�/Tn����vg]��^9 Pww����K|�N	m]S�r�j�L�s�^�R�g��5[h�+J�2k�LH�I��)�����R@ҥ�&,�UL��#5?v�'�ښF������dϏK6#oi���5�3�-V<����W�X��o��{���� m�u����2�KJ���uS9*a��{}�ESm�(o����C�.P�	N�ʳ�m��ٛ��M�� ���3�rE&:��-]�I�ߞZ�0��������tTv;�p�FxQ��'UJ5����.�s���h(�7W�i�^��������ٴC����3�o������gM(�Ժ�\ˍl��1XW狀����x:Sj�.i>][w�v�2���hwhrg�Yl�^Gl�>�uM�Ʒ����M���<�%�~���*�)��N1�(ȧ-�A��(�Iy^��t��B��1�ƍ3�I�Y0��&S�0u���Ed5��{�8����daR=�)��D�5mh������~
"�ؿ7�b/^}�l�0U�-����y�)�����O��3�4P@ۃ�����4d�<VE��\%q" �LIծ%c� y�V�q���f" r{���'�J�r'vm*�ܸ����l=�Q&@T�����(�1�$��g�0C�ݎ줴��o�8�F�	R�u���iq"�;��^kS9����B��yXP�h��3=UF/1�x�-�_������*:�G��j���M��:����,b�=��*��nkn=I=��>N�,t"1*vR��o!����^�IHݍp��ܣ4���ڙ)�!n�1~>�ı��:�LFx�pU������;[~!��>�a��1�Qe�����n\�!�-9
b�{���.o��D��dA"r*��4J-�:�b��#5���|��,y~ƽ\�SL�w����KD�;�k���n!8�xQ���[�"��#��z����Ys/�g�(-ظ�A�7UPL�.��)D�Y�a���͕�_!�̠�,K.���z�I��n3b������K!??�/����?5�_ӟ;�(��$��Z�.Uf�W�Q`�a��{��L�i��=t�|�%9����zV���x�6�y����j����!���-�i�TfS��y�i�d��+\ЗkR�(�����=E�5	zc�I��W�3��䧒��bh��|�ح�|�;��f�t۸34��NO��w�\�R�b�>%������g�0�z��KfY����s�%`�8o�X�a�v�m�Ә����KG;&�3��@ɣ\�jERҺ�F��xZ���:ď ���a]{� I�+��[n�G$Fj��q&�(v� '����`�p m�j��cw�f��&�ш���COX�J�`�[�P�-!�w����<�b���) 1�Y��[�����qw@���<���`�j���\i�x��|��M��\dK92����iw���c�9�`$S��:�9��c*�;G7v��'�B\,#g�(r<'�9�w+���ȱj-�14YEQ�׼$z$����LL���FS$����f��ذ��/"=�Q�����=L�@Lx'1 I_"la��`�����e~�P�����ؤ_jt)���Q9�w+��_���\�k�a�K���3�gu�L��Fn	^sn��=� J�B&<�J,�]a���mj��K���r�l�>�%�m�{l4KqW�R>��$��VGM��6�����w����(�BW����-��2E�t�Ln.;_�I����9�܌'����� !�d���5���L�=��_�v��'։D���%\o�ɡ��l@�y�v%��E��ύ��'��fƃ	�{��lo��� 0'�,���ڪs1AO�eH��^�J���ѵb��Ie/�y΍�YTO�W�f�� �Re3_�U��t/�ŎI��<S^x��<g3
�]#L�W�\Nt��L�]�K孋���c3�渭>虱�>~&+�YB�i�Ӌ9�c!��5����e�N0$�#qg(fԟ�M/��Ihh�3(�S�bolX��(�u�n��vi�TA��O�L�[(����i�T�B�R�H�VA�L�;�b��-��Ǭt@ʫX�|���#�%[G(�T��2\���b��iX5��}�s����z��K�^�5�>H���F����2��ӗ:�,��z끽v!x���b6Oj��`-�|�b��ŰwxeQ)�Tu��p���|�y��T>@�2-WBbzc�z}:}�7���ؖ��w���66�i�&����aD�h�.��d�����$�yT65a�}b��Y|E�++]�}`�z�C��D���`��ۊ�4gN�o��}53��Aq%��D��$�*^p�`�*��,?���~��4yT�p��ɦ�*�(�K%ؙ9�����k3�j���.�$4�c�[���ʺ�,�c���X�o��h\>��8(H��c�!'�pP�d@x�:�K�I|w�����@�OP�l�z��$i"l��}Z�6��1��������r,*�wN�: �:D�!�WJ���^�����C�=M�v��נ�E�j����K_&��U8���BQXh����(���M.Ÿn��hT��ّ�����2Î�YV_�\	zL����_rUnKS�	�o�����/ �G'{[z^s��JM��Pu�k��e�\��_/ꒋ��Y�b噐(wV����mI2��I�#;�j���@���fu~���h{��:�L�Ǝ�@��$��mJ&pZH�+2b$�ZJT�d�n��h�YF�R;sfO5�h� ��S�/���܃�R�gm	���~G�9iO��2��8B��G9!S���<w�x��{�|)�g��*�'e�I�H�"f�`S&��.K�}v�9�z�aV��w(��n[�R�iJ�����/���+�������|�J�o�ӽ�^YW�w�3γ"����Bݻs�	/��G��,�Wx�1����5.���UzO߱���z�f�+�cb4���䴴"�r��2�y���❯���hJ�K����*y������\���7�W*�u������������=����V����|P�ww�o������߆%�����T�:�!�c~ķ��c��
��O5Cm�9�m%R�B��c`��1�S��Z@��e�N4�I���[�u�R��܋�+��|,d
�l�J�Q@�4`�-XN�Xv�Ko���,_�b�6��\{��t�%s0[����{y8�j�Ψ�z��.�b�V���D��HTO�4Yb��wr��K3����+��5ߘ}�!!��B��9��NMP���t�|A5�G%T[1�m���W�,�a��VT��$�(�|-)u4XZ~�\��h��Vu]�E]�N�5����~���=�@*��2H��;] ��q����N�Q�f��F(�i�1�}�O��A3ڽ[lbJ߭�ZBo~���,}����r�-���!*7}%~�#�h�mV�w�uG�b��# ����:���Д��4T71K����؍�P�{$<Rg���g�X%Ѽ82�I�D��4����@>�)�'3y.�́��;���]MZ�2�����I�q��io�'� �5�Ɓ
?P�$s/�O|a�u��|����+I��^���a}�dB[�7�R
�����A���ϗگe"�1ssk6��{��ҋ��}�k7_��G�;^�����vM}�pOѶ���&���f���^�wE�i]���[	֥����oJerJ���5^�<���>-ҚQۗ#a��t�	··��}���u�	r���pW �g���xv����y�	��˩RI�S�r���X�ؕ�M��'�^�[:��o�(�Ϯ�d���h�M�^N����
.�uF%��iX1+Fia`K��꽖�
�����6���*<��9���9��6
F�562-��h���_&��(���$*5�9Y�v�Q�n��U�rv���+ɇT�v����"�tf�n(MSf��w��C�]�F��N���`���ޜ���iV�ׇ�#�5SC�uઘb�>j��s˧S�7�t;�%C�,�/�/�a0�,���w��})�I�&dL��.Z�����f�����L)T0},H�K�L��Ӄq�U��I�,��oƝ�z��g��0�1��҂��F�ͫ���l��I�9i0�ڽ��ɨ�.z�0��������I�_�i�y
=rp��5� 
���)�G�	��=�s��@��H�]UA2�� ����K1�E_uc�;m�)*G�H���FdzI�,�Ӈ�:����q�ɒx�3 ��B*�E�c����t���hl/�⇧fż(��kM&��R[���Z^@��'hU�K��-�;&ؔL.\�!�g�h�'�|�����g�t�Q	��4.��&d�^oܫ�_� �"Ū�Q�?^e �`)8 ����{�a�Sb��q:�������v�%�)^6kO=͐
��l�E�n�yu�̨�ez'��X��'��y��	WJY��*d�"iTM��|�Y�=��ә?a�ooFAM�b�J ��.�`���oc��Ѐ��F���*'|(?�l������Vì�^'�nH�ſԗ��޼�ZY��	�M�ܖt3�Fȹ
�JL.(�N����ځ�;V�!��� .��n`�'�Y���qC5@"GY��ϳ��G�sĂJ����cOµO�#�E2�}�v��H�z8��Ґ���ޏj���,�a��K#h���l)����E=O����e�6�(Ը�eXJ.k�����.����	���S��е�3��vs��f���~+C�eR���H�Z�C�+r�B�RQ��s�cxCU�3�s�Ⱥh���m�M��D� WcdG�ۜ�L�ӱ��2���WO̊[��`n�-ۿ�Y��\����P���<u9
�C7��k1�ئW��cL�G���4,���*�L���T��!�tw�`I+��y��<�«�WN|��.y��AӓF��k$�b�<GC�@�W�'��J��r�o��6���d�̅};�M�y�t�y��`p����8���5#�ӝ͵�RvhBy���Je��#�F{ -��W/.՘]=������S3�Y3��lU���Y�w��0ɛ���&�g ڝ�_�.`n�#e t$e�56(}�{+Ѧ0�.[���%Spo��,·�Q�=s����>�S�����Awo��$�JH�	��1��+ @���9@��vŐi&�d�b�͹^������6zR��x�+�RhБ�\���E�/��������C�n7�0'�gS�_�+��:,F���W9嗼��W+j�#����v� 0��$��:0J3j^*aw�L?��c�	�p�m5l$��X"c
kG'ʛ����ϊ�nk�Z���}-�`}c`����aPÅm�KT���1ry���|���$��,b^����?�ڂڠy+��`�R5;���Z4�hι�b���'�/�"��(�~���x�y�Y�R�RL���
�ggԽ�;�,}:�S�>�R*�B��k�D䛖�}���"b�����Io�/��l�����˰���'��h�����B��'N�<�vRG7�җ�/�-y��F�S'wr��4h�;�!��vH����'�c@v�*l��[�v6�~?_�<�x��j~_D+@?�W�I*�x���w7���f�O��!�����(�V��|����������C���Rgfso�;������Q��~��hvN3��j����؊̴�����2Ppkr�[�g���o�(L��v>08l�!:y���m�s}���=�ń�Z{h�4����~�Mn�^�3��^
D-�ܗeΈ<�������eZ������z�[�_.�2���w9����"����+���� ��eȀ���-S�����[���f+��22X�,'n����L��dC~%&[q�w��\�S�jf~rIR@/��T��T�"��_�躅��4�!7�.@��>^�E��1�	���qT���ռ�yo�܌�]�K2�y�A��\c�b�+�ׇF�Ƨ�ޗ�{h>o��ֿ��	+i�AB{��2��#���H��+j�:��֏� r��L�%����!G�p�t�{��\�� ��z�c��6
��>ɠ`�U-�2�UlB<�#Y#�)�~��<� �����k��ȴl�1��)��:ɥc�?�϶f})Eg���+�rw�T�5�*ؤ��ȉ��70'O���х�&p~Ԭ��G��P�;�	�Q�%��K����1���#���a�<d�חfN����q�3������G��*�ON?��L@K�����\S���*^��7a�2�Ožw�t�G3���U��4��ȇ�7�1�x	oJ�*R�'�| �b51�{cӭ4�99�$�p�}�J�<�?�Fa��v5/���#�_)��R�7/7e���� �t�M���{���c➦҃�p���I� ^����],������ȁ�G7��<�h�kO=�w+h|�G]�ڭ��&.�RY4#g�I�:�x���)|�||�|np|�����OsqOA*j+T'�5�jFd��!m�>z�xv�I�a*3��4{4]W�7r�[3l������(����׳4��j�TSb�g;�;1���)9���K�3lQWo��ե��H���)���bl�khgX�����e�9���h�%�wu�K�<�]V�3Q�L��eK��=1�"Eyy	�;}��фdz+S�a��@�Q��%vV���ϵ�!���K��(�eh��[�g�r�[nkk�:����+{lvf��������Y�_�������Җ��`:쐖�J�Ap��h���� ��gk���yt:^sh�DYe������������g�K��8���#8.�����a�C)E����r�MV��1}��Je�څ��OY8�� oENB�/���j��>71}�_�OdbH� |J�yĶnԤ�49��*/Ô+$�f-Y(Ѵ��Rb>Xݼ?��m&�G��	��C'��Ŷ��:x:%����_�̀�Q�Wu����_��G��fTf�GM���N��Sj�0��|����YQ)�7*Ѳ����+7ap��黪�&��,�&�E`���O�<��)�̎2$h"��y,gZ����/��y����"ا\��?�q��	3 �����$k�y��jH�!��~]N^#�gf
O�jeN����"m��S!S+̪�V��������nC��f�>�@�5�t4v�sq�c�7$y�}��g�5�%>oQ���y	�{��VҀ��B$���c�៼�S+,u�N���I%���=hw%!1:0�
@ORf����{��2	�pR\�.��[����NU�Ɂl}��f:(:�#����nwTۉ�����"`��P-ܚ�ݛ{ H6ƻ8QMF��Z)�맛��(C�y]�t�@o������Q��BEB��$ܚv��j� 7wVz�P?�,����M�����K$��0(�.P���B	��8��au�y�q�l�'��$�c��L�,���O�'�ٿM�?Wo׎5
v
��)��i�XK��ԟ���I�Gh��#�z���bsxVx��|����X��H�l���T05:Xd�_hd`�[z�������勹�,��d�ve��_K����M�;�ؔc(�p��"�- ��HyF��<���:<'.v��r�"����������.�k]�q��kt	Y�k]#qm׸ffE�*����,����H�k��Hq�H	-I�}~����y<�y�6�P��{4�Y��$����A�P۾W������Ey�:��9x��:����}U{$�~�)���M����0��Ğ-��~=����,��:�,=�@7,f]ž4�Ox���g8ڨ�i��F��N��N��e-:�!B� !ަ�r� ���@�y�/�P��������j�[�;��!�I>J�Q��5
�b�X$G��	&s�rQ?�6��q�ѳMx����-D�[&�q��v*�2������-����������n�Q HC��{�?1cr����g%]��>*�aK���g�F6v�zo�����`^Fg���������� ���+8�V��1&��ɭ�/�
��}�:�ɩ��y���/��R-���L��w��l��=0/N��iZS#����@_:\��mE�����Iy;����PUU5<l���������V�'��#+�x��%l0i����_�
m��|	�nV��Į��+qKt�^{qt{�Z���lM�Qz��$��.͚��\�Vh^�,�������j��4����g�/�r~�r��w��(�c���}��#����|u�*�RS��Y�8C:���w�@8���a%��M}�u�$��3��GO)��c���AL�����P��xf��.L̘�|���u7��xtq�$F%+��?^��9�7�6�ː��B�}�jژaY%�jt8�X�����q�<�7+H�*R���ŭ�:�j^��I"5\ۨO�O�+8T`V���P�	&@��\�S�!���!K�]p�0�3���~	�h�U��!2O�?�4A�(�8^�\���|.�؆S9�@b5��{�xIJ�^�O���w�d,XS�V=�LR�G���*�e���]'�Ǽ��̗gG(�9�F��6���^.y���x1m����["�?t\�7b15}wTP?�'�����0n�����29���#��Z�.�]��Ҷ��f�3�E���	k��	�V�w8���5�P��(�I_�) h#�Gߊ�TTJ ��y�b��M.ԅ��k5������Y}��Q]t�k`�P��z�h�,�9�4�� �/����J)trE�0,� �Y�:)ʫGk�q�[�q�F��2�"Q�W��3e�s=�&���P0c�䴆��f&l�dqbV8���:�jHp�4�4�t.v�W�w���7#�b��<å".+壶ۼ�������V��ծ�;�	��
�nїZ�+�ҿ	��W���~;R��B�ǆo�+�ֿ���	�
{Ny�N���Q�*3!]~!�.D���h�k/)@�EnRj6=�^jJ��_���:J������.�ub*O�{��#�2�i��k����w}��)��i����G⎠��]Y������D˺�m�iw��{��רH!��M�v�����.�����F� � �Yi�D�#�7F�����L?c�!d+�!���,�!q�J�X�'c������J���ȁ�\�@���V�4���0ܷ)���w�m3M1�����,k�m�X]&���Oض�9��~��V(�2�|��ч�#�='x?Od��� (�e�/~�L7c�|����k����m�zJ%������;�P�ͳ�ex�����k?��B�-^x�0����Y�><���Z�nt��us0)�=�f�h�ݦfڂ�3����_�ׁź~H|Ͻ����l��3�B�s�e�*���":����k��< +�(qz�E_eK��j5%(���)�����/Px(~����4��U�ϷM+���R�������2^~ua�����U��{u�8a����;z��}̂u�jw1' ��+�~�4ʏ��6��� ���`R�8�D����פ��+
�������B����B��?G�f0?y�9y���3���մ𾨑!��Wqms��CD�B��:v?C�̤�څ�!�̧8�ـ�ui}�C*��*ulv�|sԐ����%1�H��Bv�'.7����3��e���4� �K��n��*	ir�+R���5��9�7&-د1 uq�q�U�$j%?=+O������1}�b@~BqSV%1Q�O�3B�\�@��)���iא��?����=`4��e����?����A6�,���`!:�rР���A7�̘�"�:PH� @�bU�}/���bg��S�H������K�ˊ���7��}§[}'�t�[1Rm�ٱ'R�w�vW����Av��\�,aPG.�오O�M��k(Jr�ehlG��2R� �'��B�x&���	2^/lX(AW��v���hxo��o]Կ�H?H���WW�OU|�OB�ݪ���<�EP/��fN�펀z�c�����(#����+ۢV��%�!a�lVQkֶ_C��ϟj�M&}X�Կ	qǡ�z���[hS��8`�l�>/��],��9zA�i/�)�v��v�`�����I9y��D�c,_����wf}[t%�_�W�n�ِ�uQD�%����;h ���(����Q`�i�����@�ۖa#�l'���
��=X��,[��j%�:D�),�I,n�2	bM�A��Q�Tn�ˡ��>�T�+��ӄ��$k������ �a~���������&AY)���ϐ��K~QH�X� !D�F�n��9�̬"�L��k�U�LZX�B���7�s ��A�k��&G8��Oba4#|�
��4X+w,�'*�ŧ�Ǭ�AYY�~��8t�v���-��;�-�ƹ.qOk~�2n��o ��K�ҁ1��J�A���[���Q���������A-���c��,�����kS�	$�������/S|p8�/)�L���r�D�¿��6�P�,��*H^>�0B�f�;� `��J5Nit�"�w<�K�XSI�{�ʏ�����Im"���4���3�ԅkv�]۽ �;>�{����� ����/]�"�iK�767���W��u��%��]z|��~���Zt8���/�����?��:c}---ϟ�
��V�;�8�u�4�j����j�?b#_�*�f�p!mNT�_��4��� �Z]-�F�ܪ>������n%�c,�[K�/�i?� �Hs��K��w�R����C���7�qf��2�n=���{h����|����[5�Ӆ��o`����"+�	f��HN������Ϙ�b���o7x!�����$}�V���߽|�E
5~C��Nbp�(��`P�1'o�Đ6��v�Ŀk������;,l.�x�����(X���3��*��y��ӯ�պ:�'��u��&��ݓ�%���Z�rJŬ���'�,��N �8�Ǯ ��\��DsN/(�\��~�H�ǜk����y�Ƴ��.��t?�7
C�Xxm��ʃ��.���c+��7���w��ڃbXs��N��ԕ�6ٌ�/���#�J�����S
��8븵Ѫly�B"9�*^�X�	�6�X���4@��3�2k�++EP\L~.x4���{��f��G*-�4�7j�u��TkDEo�Ii.�j�wTQrw��)Ci� bbԏ|W�M�=[$E���9VE�ו�n�0��m�^cM~F�Y��@����-��J��u*Lb�w╎�ʟhJ���eI`d'�%�skԐ J�<q���*����C=��%�c�U_+�J��J��3�ɅAW���[ͮ�@8⌫vP[\�t�Jk����a6�<� ��p�*�.	���s�F�C����*�{7����މ��8�d�Y8��$]6,�nw;�q�����D-�ʢԥE��zN
�S���:\�gmC&��5�\�4�d�}Pf���Wc��0IV���u��e�����#�b���j�4"4N�v��ؠIY���e�i�k��$t4�~?���3�%n�er�V�����/�S�1�?��. ��D�|)���W���P�����u��;�@���9�By����ct{���'^�r�f���ʾ�G�2Ѳ������!@Μe�6�����D4��t��1�t�X��!�'_)u'I)�MN@p���P���X��ۋt	�F�.`����Z��k���G}�k��Q�mu���a	�v��@�̜t���"Q��k�K�Bk>�����P��Ќ}�7x-��~k-!р"C4Ԟ>��������˵�q�K��A1���W�=T��j��^G-r��ީ����M�)���a���"�&�~��@E���W˙
��s�qx/��ǟm��y^��=�/.�L�(����s%y��#Sx��4.�� #��U�T����?���6�5���Ơ����m��D4๐K�޳ث�T*(�g���_W�)�X�+�T]�6���/!��'����b����l���B�t���S��ȵ�j�ׂ#���@��\�񻠄o{޼���t��~_1$��N�M��D���ϭ��A�yۇ��� 7��7��G�~8M���O�����,����R���9߽�=y�_�Ե�<����O
��`�,��~O/��w�*5s\�[X�n,*ʼػ�_T�d��mt����E�՞��m"�#�� U?Mrv?�W"5N~c�����b���:&\w���b�,��.�3<�e���w�F6w���}��ŏ����w�s�g�Q =��6~z��}ہ�����QS�6��׀�o��Z�U}p�<�#9��7�Z@=i)�M"���/����۴����;a��D��w�gU#���9�l�\iy��M(G�Q[FZy��&��pAy�a���O�-����v�}��|�|�.�u�o�o�� 8Ս{P�;EF�Ǡ�������G4�����Ĥ���]˫I��B	w���xE��Ⰽ���8�C<v�Tܯ��/���m����Co��^6�����U�l=s����͞zm(�]��R�xQI��c3���X:X�l�� ;�u��5Me7c$@����-k�|�Q>]��~�����b�c�D�m0����9S<Q���X�����>N67���ޕ7�����1�,N�s���D�E�)�b�����B�ezq/�it#�C��IO�L����@f�i�}e�z�<�H��-t���{��	������/�E���v'&α<7o�FN��L�섢��wf>�Yv�J�1�5�������+�������y����{��\�\S$���M�
@<�a �;�J:�FYjH8w=
 �1�4r����Έ.?L����Q�=���6 p	a�'=�45U \��B���X��>I[Q�v�kS�04���_����}�0͊i�KH�Y#ppј��e���Io����W�ˑ6�6��(9:�(H�C+���B݅�)

��:A^�jr���W�����?g�mӔ�y.���f�{�yr�F-�j.0��4���	�i�R�W�s++V�zr�k��N$GSB׆�8)��Ŧ�q�D�}w?��M1؃I�
����d͟(��8����u1!?*��~4B�˜�܍U,-����[Y���,%����s��%�jŮ�|\�e�	Kv�m|�v�G%$^��v/�5L��	�o�롹OQ��0Q�$�+����!�m�8~�����z;���F��+�ΰ{p��EoU���?�����u1�����?��?O�8"DÙ�on-ܸ�8q��w�1�ѧ��a��?������� v��W/�ۇ�,^�R��~��C� �7���y�:�tQO��t5F��p�J�נ?���>;��ZG4��}�]����]�{��
MM��J�п�0`ET���wϿE�::a6��ܵ�VK���IQ�_����u���gͩ������Q}<���p�`�P��ŗ?V����_ߥ�C;ݷ���՚��O�~)��jZW
m<��4�嵸qcz���Mz�{HPJ���E3+ hX��8�����M\���b 3��TB'"+a����(��H:]�d�3�Om$�f1b!��˱�1@�N=NEH���s)\S�u��ez�@��H�
g�)�^K��.M��$P�c�Uf���^1t�|���Я��2�8XCE��`�H�aO�)9{�$��֤���;g���#.���D�>:SK��'G��@Gm>ۡ��@��/��z��	�Vf�N��En����y��
�W�u)A��b�z�wN ��]"��i@�4Yfs� �N4.~�m.�X�3�r�62��:C�k���}3�x3��y�dIo햑[��K�NP�p\�{K,���-�����8�P`��͊2Ge��K��G��F>}�хF�[li�#Q»3!w�(��w> �����X�y�T�o;\W�ni��?�s��j��X"�	��v�їL����1q�-6�ы�+�m�;k$V���6���~c!��pĜ!c^�B�:82��k]K���/0�m�4�va^�(ק;����&w�O����ۨ��o;��q�������T!���CKz����5�����m����#�.xR��>]vD��-���c#OiN�\�T�;(:�㠅��;[*Ɉ�QRH� ���A��|;�0]�H��ޫ�����<JkCf;��SF�X+��#�z09zJ�־��Ȋ���Û��эhL�J�J6��`�Qo�q�ĕ����:5}�Q�0ZK�*�4oZ��F��pc,�ˉ�aEt)����FKvo�=� 0�ݩ��$6�\��%�}o#X�.��ea{����7�=Hӳe8q��b��6� ��:����2����,w�r�we��*��Ŭ8�^�Deu݉�e��u�#⼞��k��	W����/�;\�̽A`$9��	��ڃ��
�N&	�Ju�.�`�%�'�E`�J����Z�#'�bӪ��뚚�Rc�Y:Z����Q��?}��<m��m4�J� I�-������i��,�1*�f1j��� �?p���-{8�1;�����AS/D���
>�zY�U��9|���t��I�";$X�w�o����	3c���E�9^!��/|����9g����+��׾@�{�}'���b���ޝe �_!�t�����K����%�86�5�9���䟊e�wk�C�Q�wU��.>�KP��+��@��pUv�q�=��`+����em� d�����G׵mL��e�W��V,2؅#`�q��z�h��P����tWs��}r�ۼ���'?��է^N�q"��|��vЧжƌW1�e��1�r���9���ѩ�p�nC�����D��=ns�˔�[ǒ:]��3ӟm3f�^' �툝*�e��~�	�;c��)�GiZ;~n���2�ܖ�X�k`�b�+f׌"�D��*�3#�x-���G���e~�r���ձ�l5�m��]���8���^�bSjE�����죌/K�zr$�o���
dyw��3�m��4��DK������Ʋ��K^��:Y�7u�c�/�g��O����:Y�P:�y�o��7�+�DV��^�Rԅ��SgM����j%DG��Ts���z��;K��t�����B��ic��������
SF�����|?vT{s3\�e��2פ#��O~�F?������n>.�c�,c����`�L'�df�$�Xy���Ö����9�y!
?k�X&�%^o3�65�*��%p�Β�Y�8<Xu#�I��m�*�K��`�t�G�к��>R��ͯR%**2c1��|�Ve.55��Hꔾ��\��� k��*]��~�ba��7 ��c�����ٔv$T���y�� ���خ���a0Vt6�����%�@�c9����;H#��6���_��o�[�q����Þ4Y�$2p�3�!��j��ܠ_3�e���;^�8���Wss^͉V�CuĄX�.�ݙ�4;S������|&[�.�rQ���%���p\��p [�bw$<������[0�Lc�S^��?����9+���;�~fޭ�#�o��~is��jhו��P�t�U`j�����j�/PҼ�y�*�	Y�*���] S���&�RÖV_Ҭ?�[��;K�M���oH�枨,�������P}�E��`�rC$���*%`�l��Ku���x��8�t,�W�g�`��?����y���!;ӊ�!��=f��Q'>~�����R��Gy?�������-�I��/���3{���R#�K��/��x���"�pF ��������b{*���؇�J�9u��RkM����J�����n"��׫r��ߏ�^}�һ��)W?�6%��������||��G�Jz�G�	,H���"���4�_�ޘ� �r�7g�k����_?�"��ڼE8�C!=:���gg�[��>%�m׮{E�,L�k}�O�\B�H�0by�'�w���)ߚN=3NTT�0��1�<]��q.*zaa��5b����ub8}�Y�߰~q�+>t7'��~�!q�Ű1�Ƨ2�8ZIu�k�6��B	u9��������.a,���ި>���ˏX�[����zZ.$s��^ ����c�8�	0l�(� ۶���H�I��2�i�vSB#�x�q�-r?oQ�~��>��w��n�Q�怚�2$5��e��y�w{:&|��|�kن\}^ȋj|9%γ@W����d�����R��-1o���/��.vZS�1�lK�J��/~�X�g��ZF��ˎO���Iܩ�ϑ�o�9X.���mTJff�<6mߺkL��|�~U����HPx�bi,�2�Ӏ�2��{-���]����"�/ܓ₃Xd'��ik=H��x�9�a��#��q��e�����?�}�ַv�S�6�:��0C�����q�NA�be�c9�v�|Q�rL2�������߿'׶�j�_ �H��6��3Y�w�<�vZ�R��.qy�9[-�l.�mo`��;�'.�4��mȗ�.?ءӉ�!�f�����.��+��I<��B/{�lgh���J����@Qw�����> d�U����Xh��*���8��6�|ܿ([��A���'�9zWg�m��J�n��%����M|��Kg�QJ��8�-R΂�[�6,��Z�.@�s�1�n-1�T���x��O��p�RX(�j�k�.,��b����e�����G������qrbڀ��z7�9v�t�f�+��[ţ{"ՉF|��]/��r
f81L9u�__ﰻoS�Փ�9fJ0x'�y;�i#\�Y�c���SX���i�L��)���V(\f&�Rf�oʹ�M�䙷{;!0t�@޿y��p��5s��F%���;0���7�+�muy����l��w|��ʗ��pM�B�9_
����t��7Y�	��io�i�b�V9��v)׶l3�v��z騖�'lb醘TI��'K>��F��b��or��6X�s	|���$3%���@\x|�ֽ7���X��}x�=,��W��A���W��e_w���Lipr�V҇uI/���%I�Fw"16G�#�{�Y	�7�(Ex��ak�acXµ���6<�����P>F�\gX��p�h{�m������}�\�@]��qii��*͞���%Ӽ�e���5���U�o,e�<Z۽���Ѭ��{�$�B:A��u����v�;Z�,��/��I]�KU:��Q���L�iHK�R��9�ʧ���?+aW~@S����/>�/Q���}-ݾh8T�A>Ŏ�ܶ���������(0��&"8Z���֎�=o�^�̰)GY\����#MCM��6|��(�N�r�/-ؿ-��R|)��o�!o������-����%ٛslS��Ł7�՛/�p����;vSl|٦N�{�k�:�v$9��\̫S�� 
�ALZ�%��K;�)qa&��h��� ���C?���-�iύx�s;�s�HܥDoux75�"H���٥L�S�$S� �	��N=�X*
j��q��#}�m ��G��;�Z�u�6l�0-�Y϶h���e[I��t�J=��V�l]���E}�o�u�O?2J��4�gD��<M��<7�~h�;6��_n�e-�!�X	S����ac�׏oUj(������T.Ȅ����%Q��h�N+�%4TD9�F>n��lA&1Z�]������gv�r�&'�EX�M~��q�Y����9{dā�֓vPy�R�0v��/,��|�jCGI\b��]K��%�Yv�hW�Nj��`\ ���K����6�Y:�^dlٯe�c)@cw"q�h� �� �V�����; e�7l�G�NXy�����v�%kpL�+w�xL��1�'��S�{���R���C�i�7�M����D�o�N����������+�$��4�ON�0}}��7eLSRC��������g#J��~��3B$Z0E�k�����@7r���B�k$~�--��,�R3�����Q���ō���Ҝ~�!�Ub�ם35�U�0|�.3 I �����j�-Nw)�w�5dL.G�,$���sR�~*ix�E�a���>�H'�7S��1�����q{��EPY%B[J�����ꋳ���6J'���~[��Bjj�E�.vT�i_�M0��P�����z���	�{��l�m�4[�c��T�v�6�f��g�a����~3���u��˕_5���g��cnL\���H::��zi�v���T�U��'#�nM����e�3�u��cI��������5�fg����p��n�m��g{cXPz���;��75o��N�sn����_mL�I:�h��Kyý^��k
y��_�!�ƈ�[$����O���_3��Ǽ�-�45l����F���L#���k���o���=<��f.gn�P}�O��SG���}�3��0İs�l�#
����9�"��/�K��0$��:of�
�:f���l:b��S�	��k�Q��K�J���>�~���q��s��<+�g@ʻX�t���5�`�������3 ��¸�r������rC�J43/������MK �pka +�+�`�G�҃�3�z�
d	��ŵe=1Q��V ?7�k"Bs�X�i)ǩ��զ�CA>
�e��\�6bDf��$v|�~�R�Rp�aI0�g�
��^A0��T4�Hr;�?�}#m281u֦�3�C�� ;)����l���]�FC��p[4ލ�{�I������>������n)��PHP��-јF�&<'1,ь��b/�=�IV�Y���s2����y	������X�};UeC��{fǖ!g���&r,o���6w�Lcܐ�B5���^j�*���'y�@�4o��*u��8�#{4�~��*i�����aXC�����U��"h':�)�	KQ'`���L����b#5T<�	�D�Z3�tA:�|���X'�^+3�T�^�԰��A�@NV����ўG=7��'02L�O��R���0`���N�!`��P� �Hn ֟M,��:<c��ۥ��n,�#�J���1�6�E"���C!	���v���m֐��bKcFui1���8�u��X�1)��f��������+z�9��7``��o�Kҕ�8�k����7�;�� 3�yy��Y~)m���^d�&��U��hR�bA�}��W%l�2:�۶/v�^6�F�O��>\5�Y_��: �d�JI����\e[GyXAT}Pcq$�����Kv����1	l�4���v����T��G��Kwh	Q@uv�[�1p��"G�\&�Ss��H������#2~BFי0X�8�d�C9�2�t"c'��k���,����5b	��	�N$��,��bЂ�%�r���$�(�3��h�w*��Sd:�_g'|�Ի{���=r�UЫ�gX�X��$�������� �Y�qk����]'t�:�.�޻m��rז�N�
�e�R9i�J!J��R?��A5Fz�NX$g��UC�ɟ2qA}������xW?��V��8��/yȥ"G�=�[k��u�&�\�n6�<���6ȳI��Y�*��� W���e���^{̵w��sv3�T� U�c�������`��Ģ� �����g����A86S��;�J�~b���	�9�I�f{�B�c��_����#ۺ���i���j̦VY����{`�A�noQO�f<����}hM��X�\�C�jG���|?[l���=m��*$q���MW�w���ٲy�[�٧As�t�w��p���KC�� �@N�_Fl�a	���B�C��k�&��_؍�d�qwpta�o����M��j��z^(&v�뱯��f^._wDF���	ڞ����ĉR�x�j+6G�f�N�B�Q����?�>--��9{!,y���0P�==��KEI99�@ѕl4sP�������hx~N�ac�c��=��� �4P�>IU�~��Oξ�o��"y��*�+Q#]4�K;Y*���D��@�s�M��N�N3ğ%��`�
֩����y�X��Ew�YPq���ue������!�����J��o�;S���������o��?���'�F@K��+Z �� ^t񩔣T�z췻��o���Aݛ�LX��<�w
�k.tX��#/���O���d)*+�:ݘ��0x��펛�ov���3��Ё�|y�;1��������LL������Kg�����9P��!r��ߊ�@�7'��O�S���CsK�ݩzV�G�?B�J�,q��0S�)���W��P�d�^&�8��mjN��W	8MW]�?�f�e���u)��u#�\|ƞ4����,�%��ٷ˗��d�.A�
[&��s9�����
��^���["+u����@[n�����`!l��-_��U�*�BAv�N���Y�b!��$��]��AkJY�b/������*�X��&�����=G?k4%ji��~�Є��ůzoS�����륫�����l�@��
�4�E���J�O�p���NkQ���~��S�?�W�jK��F�.�S�e�����ׅ���t�Y�߿�Q��mׇ�FS���<Չ<�=w?o��YB�m~�)vu��M��?���K��ǜ�W��������j�@�IJ_�����d������Ճ���/��X#�W�.ܸF��9�'�C��S1���YfU
��n'!\���_�ް�p�y��t̘[OYeqo����5毛A�W�?7_L��Y`,el�m/̨P�@˛=]��nij��N"E�_��lLŊ� a*�6 �N��6f�pq~R��P�_�/>-hB�~��4}�Y}gk����:�Ϡ�����J����Cq�8�Ut�c;��ڿt�.�ө�t�$��O���N��t��l�A;v�h��{�#p�bt�$Ӗ?k�2�:�%�V�J	$,7_��M�&a P�Q�d���K�6���6�'��V)�|�*)N���O:H	��}���.:PÜ-�w�";(KXT 'ds̔w�n9mg9������ ȥI�#/�Zu<��)K��"Ec2��;Gy]�7I �G�<}����ɺ����'sE{�ۖ�GjGf�O>6�#�F�L�6�����y�p�ӁH4�	 ���v��Ӌf^'��5�V����e��X� oQ��ϚkbY*r�����U�Ua8(c��Q^s�s ���y��(���4^�/�1����8�q^�"%׍�拭��UE��v �.C����(5����1r��6�\��u5c��@�ދ�}J�1�E�k院����?Dg�e�=�!���]��淑,)=�_"��S*�J���M:�O�wT���c�Kv-9?�����Cޓ�EZ��!�3ۀ��S��V��7�2���Ek�|̗�z�(��$u��J����)���2�5�����r����kf���g%�O �`ɶ��#��v{!�-�%)E�-&@��8��̏�{c��@�����L��E2Ь@��)k�Kh�eTp��CK��xi�y@��o��
�2l힨�v@c��3���X0� �0��$���6��*)hǋDڑ�� �+/��_Ӹb�
U�~ݔ��bb�x�q��c�sC�J&g�����Ի�F�y�BV�Gaa�{s�8H�#�sW=qn�֤��Ĝf��"3ܣ���۬�.��(�8z%e�V�0c�D�Y ����a��Ay/��%�Yh�I��)����igwp�"]���e�K_jc��ooL��ď��3Ɍ���WK�ڗ��r��liT!n��@��(��JڪL��p����|��������\�3�&��.���C�$�cǝ�����x�w�k��F^�4�����V\ʰ9�^]x}bKg��$��S���qB �A�/��~/��"���K8966r{l�H/����>�E�&_r���am��1��S���$�U�k�h�ԇׂ���O����:i�sc��)�a�1�j���c���{�	c�G��}c�ל^���@�����-a�	F�[rM���C_�ѧ�!��� ^r�����?>�|3�)j	�Y�,'���%���@�����g�؇�q/sxEP4)Δ͞�!U�;�Go��� ����1���_��t�/
p�m����o}�/ޫ6�^����xil��[ײ4Q6���iR�%	<2�8�E y��N ]9_o����ZX��Q�-ʮLZX�T�Mj ��yS5_�"
v���I��&&���Iz�T��������X��"�	�Fӂp:RB��dqܦ��e�$;R����v;�~����!���mX4�m�=�q��&�[�`�E81��c�W�6e}���к%g&y�ǝ�>`A7A�S��IeZbhGt:�����i+}X�rI�����ӧ)�����h@ir��*�6��J����SVj�flp͝�W��c��"�8c��UM~%�L�ڢ�Q������5����!�F����Z�}6�}����������^aq�gS���4g���TT�><)6nl�q��6�@DO��=d��g�i�d�ɰ# 뎭�Y��V�����P*�_K~�N���fP�M�4Bm��$
�O�^���]�D:>�����~>�����S�����e�㕦���|����g��?>���o��g���(��S�,"�����v�Fy:/�U���9���L��B�i"�7��'m���-���-#Nl���><��y����:e���1�~��Όu�&K`uQA�R���5=0��n��`���k1��W��zy�֋�<y�ײn1��n���q�ʧ�G�zy_^�v��m+
����JVx"�_rH�~kC���)l!��D��r��K���뀚�wO��۲���,4�g��>$~n�̯Wg!�<�Ѱ9�`����Zu���=�}�jU�S���F�}=�h�P�)Tl��sf�*�f�$~*�\�i	�;�i�MOѯ��b����O��7�/��bE�'�&G/���+z"�V�١<F{~[�6_���_�t+�_�|#�+4��G��K�Ғ_[���d���W�Ө�UۣZgJ�eO�}��4���O-�3�0q/A�;�`o��gt����Ѧ�K�>�v*��4�o籛��ҧ�3k�7[��4��C����p׎��(��?������\����[f�������*Үw���|3��Z�I�\2�.*�}R�*Q�۔��������̇�J���%��=@� �&��(�k��b���>�[W��답�[�ǆsud��kTA�R��qx��zr�j�^�"h|�;�(���ךW��@�-˦M:͑S���Dd��N rk�^m��Q��'�LFћ/Sm�GKX�bcM�0�o���y�?����O�]�����T�Ė�i�����,�L\�@�y��l�r�bR��yC@yՍ�{)zFP����ve2�-�J(qb�wz<���V��d�j�P	������5���K�J�b�
Y�(O�S�!;,1A�`�x�=s��|p�WJ�ˬk멷��vlɄDP#���� cK"�^Ae� :��	��b"��%���P���1j�{pW7̑�'��+R���ƍ�������m9>���$�����kCժ��/g�~�n�>�[��;p[�)�[A�jÙ[��u�q݈�*Y+K��c���̸��i
$ٔh�4zW���� �1*����� bpvu"�%��wl�ɔ�a�FuCH���R���R�n��JW�>:��/gnW\��4�U\���G�ب��B9J)�;����薒�F	*)� �8F�HK*�" 
(���_����8�{���"pO��X�XHګ��Ҳ��\�WӚL�
�"*�q�(�#ہ҄��`e����9T\le-z�-rg)g5�bq{v/X��o�-�U��OZI���:+D����~T�%�G
�)�0k�Lkhո̈́���*�r���N����1���6�Uw�ǯ�������p.��b�vg����/��,�T��xGm_�݌��̲���x�s�q �6�u�~���$��"[)������$���~�5�~�;(O��dY�"F���rj��k�1~h��=;x�\:$8�d ����ě+3a$��*d�_���P��s���}e�;�6���6�)Ȼv@:o�4\����;7��դ?�]0�1]mQ\�+� ��&�"h>�	<jOt��Qq[QL����W$
���R�!v	�T9�񰀀Yb�Ye��iR���1�cE�yO�1l
��Z��Eʃ�5hTiߪ}�^��z�\�n��%.�\a[�(U���|��A�Xq���pE��|��<ghuf�і�nX��L=l՛��d�e���^���Ŗ�����)�3X�!��=�&���_��Ҳ�W���h�ڹ�'�Vf�
��{䜚�`��U5M���h&�"s�p�G�hO�VM�fCu��� ��
�O�T^ԌVj�.��k��4�紦��>��ir �:�GT�(�J��*G�� -�{�OrY8f~�l�M3�4���Ԫ@��{�C՚I�-�,e�Ts�O�Z�(�T�L�)��f
pUp$�6�� ���$Q��q�2�[�vК���j#*�W���N̄R��x+����:�h��@���ٹpM�2/��<��4v����t��@7��8����H��ݱ������:�l�����1���I�Ą�*��J,�K�X�Y�P��b�{Or���-�BFxQ~����[Nǆ�1��
��@m����[OOm��U~���m�M\#W����ܝ����ԝ�S
�����9C�{����{n�v뻷�^~�kt���S��ٻ�Q#�~=�{�B���x�R�V����:�F���1�5��1w��ďXfRUy3ӈ�Md��
�ک3�0Up�q��IK������J�ˏN���+����r�s����K�}h��M����<��e6��1k 􊹨<�?���H۬�ZLi��x#�rͫ�x|lq���*�9���<͘���Q�D��ѳѱY�� �@�Υ�־J��l����;��!�18K�\���nq����;�6y�7��\{>�h���>�Y��!x���:���	����£~�n��%�wN�$�Y�X��䮨ڜ,�`�~5��������E�K<Zq��q���DC�YwbP�)�*��%����:�kN�S����p��z��Qf�����-F��k�� l&_�z�_3���M��L.�m){�|�7ƹ(�wٹ(�����l�'�� �k�Y��%W�BT���+䉏�Pj�\��Ӭ���-��._���4�q���+�f�rTu�0�e`�w3��A�m̑zX�㘙0��-���b+'�|r�G2�!1�z�BFk\v��ͿDakך�/}/�-�#IU���'cӯG2�-1iW��p7"@䥒��L��"����x/��������ɑ���O�[n9��|�Wƾ	�,z�c�J.z����O,�	�m���;�T�m����b���*v��W��M6���m�S�%M �Ǥ��g��U>����lq����$L��ށ�$d�;Ug�Z���(*�Q �335%趽�����w�s2��|�p��"������������*���b���o�4�P�L�Es�i�6���?
=����/>B߷x'�B}d\T�Fz�sY��ްwMsƺk��0|�g�/�L�E{�Yð���]��:�����kl����Z����Z�>	:�`�K���٦�5q��ױ�q�]��tu��vR�x�}�(�P�>�rs�޺EE�6��.�3��;���<J[���WNU�"a���o��w(���� ��=m ܈����*p��'�� ��a�]���yM׳!!��4��='�On�[�������	�Wb���Fw@1@�h�z�-���z:4�Oh��ټ��;Kc��0#�/֎�( �Y߷�ؐH����vBY�[�z��D%G�Х�����:�2�Bߩ>Q��t,�a��f��h��ѻ�&xԄ��b
���ELP5�ؾ��x/ƚ���m�b>�G�]��'�hi����W_eWKK֧����+������z��(�3�󳟴1l}���gr�����C7�z(B͗��2C�T*����@��uf�(�voml��ަ�Ȅ�؄T�]�6k��m=j�w5k�M4W
�~��"�*�[�������]Gԟ����e��&F�{�e�g��b\�����56��U5��.=L�py��l�'�L��*����RA[%0/fQX7̱F�cϪ����a���]ٵ��or�I�i��4tR(2�^��GZ,����{i�{j�|�-��w�m����9&'j�9�{�S��M��ܔl��y�9������/��kL_C�*��P�/�aj?#����=͆.ۓ�i�4�7ŷ"��B���^ߩ�.�_#�^���Y�Ə�������"؆Hڥ�V�bQfɥ�$�--�{�/x�z�V��B���6G�!�	�@y���IV)��U|Zz��-�:�� �~�U�>��y?�_��;s��Nؙ�!p��R�(�=>Vu��냉!en�}�� �A]T|:71WB�wm�X3�w�A(�B���Dx ��pQ]Ab_�[|��+\^���Eӄ=���>8z#C��ly��Ig����%�ճ��s����7�Cd_�b>0ה L�n�S�oLǣ�z�� �����7ŻA7�|]��z��S�Ug+SĽ&��%��l8��Ί�=���ݤp�N�Þ��.i�&<*j9����7���E뻩��ͣlTR��L���ٿ��B��}�)&ܒ}���a����W��ǟ�U�Ù�?(ޙ!�J,�X��>p�������	����'4�[ W���_(��7�d-C|F�i4F��[�_Y�/Y}̉��up�s��A�ص�W�(<�C��O�Ӹ�Kԇ!�ٿ��'��.���\hIb��冸/w��ߨ,�x3�Ov����UP^فN"�ݟ��zy�nu�א����W��6=���>��~`�w�o��:���$�׺;vO os��c��Hj�Au~m����Z#��q7宕����qKQ'��������f�׫����>>6��~h�mZO���@��pk�X��رV�Q�p��RtT�7Y�I���Ax��L@w`w������K|��S�*	�=��,����&+]��+q�Ԭ��kj߇��|�>��R�;O�� ߥ�g�3X�����Ce�w ���z_��c诿Ǉ����Py����<���h�RB��í��m�o)Tj��\x�6�
���-`����o����q?u����܀��ح���:Ί.[�����#��ƂAQB�.��ͻ�������[��5bPk���b/�9�w9�~|N����7��
)��������,rމN�rE.iP��м���'�y��/-&I�f~4�㻜�s�����iZL~+�Z�c�$^�o?��W�v�~ʗ���I	�Q��ѵX�8��;���2�F�ߧUp6Tl�z!V����!ߏ�.�_`N��Y�{����<d���e��s�(Z	R�S����t���ĕT�:R��|���t�Ƈ�M���$��P��{��"))9*����zd�b�K���;5U�P��j�պ��_v��x|3E�⎍�+XKBC �`�٬��t�:|��`^��AWַ��l$�k7`���iz�TE�i5'r��w�9�(I��gy���8f���3,��/��|;[L��v����S4拢h"'3����-����[�����f}�s����p�Bw��.~�����l��u\�0t.���_�?��7�(z��:r?m���z���3119i�0Ȣ���+�P^���4��f����Ld�4�^�:��+�~��=K���u���gUYh�y��&&@��Cn!���j���������.�.5�a��7bY^1�����������>�&?}��.ۜ�"�|ޤ����{�o�T��5A�SF���?��y��ס�����8�w��s�{y���f��Z=rbI%�aZ<bAw*����Fݫ�k��d����U�	`������D���Z���z��@�O��O����@LF�!4���ZH7��ſ��J/0yS]�����Dl��71�ب���H��c���"f�&W<H�lɴ]��e�sY���i0Ҋ������h������������T�q���A�P��ַ�ʣ<IΫ����w34�����=]X�=�D&1B�_H��H)�Ͼ�:�6�X��p[�n�q$e�����]E띬�58$s^�Z��FGū��1�|��>a�־��M�����>X�,�L��zX���h���'�����7���|�2�BQm0"
�b�v���l�"���V>�_3?�}섨�<e��7���?�W��X�ϝܦ!}�Ui�eV>
^5ń1���P�257h�j�w�?�#aAwh�=r�^��K�a���r(� 9�������j6V3I7��9���I��T��8ol��ଭ�ԒU�7�}�,NL�I����б���Ⱥt<kЖ/�:���^�2����%>�y05"(ɸ�5��֗F�CG���B�{v_grHZds HI�9ڟ¸���a�*��ǒ����Q�0G��f�������:����O@��A&����Й�M��vHG�k�gǊ���d��J{��L`r{�C��Bkgf�*�	���
`4��pf�l��U��X��<78�msk����m��;��s�8`��FwY=��p5�nv�:�B�&���$�&�8����%�诱q�F�x#�C������T��'TU���b� 2'������^��&�˴\��?�=G_�>�Z~q� �2y�s~c�tp�-v��Vq��w�/zT�>D���QZ+s=�nL	R7�%.�_���1ߡ��O�&��H��cr��:�¦WDi��]x���`N|��?��ZD�� c�D�Nv�Aư�����U��`1&J�(r'D�٬����Xk	{B�"���R����YL�Ӡ��+�\�xucb���H���A�r̀l�O��8��$o��R�Ge�V����;jE�I5G1�y��Lvx��*�T)G�,������>3����20�%������������	sy�и���B�L��
�z�1�Ϣ'����ߌ����F�$@�l���e�b��^�֨^�����zQ�pAHi��.=�i��F���/XpZ34<o�I֚}n�|Zi��I������M����Ԭ�bL��jK�щ��cA317��L��`�3��:H`8� w4Y���<N������R�W�vT����7	8F�QƓE� �	���굘Q���Ѹ�-������%���Z��\0�d��A���0���֒	����T�z�-���b
�#�<A�@ x��^�*�_�x�>��!)4bˣ��Ի����0�e3��A	Y~� ޺.s����7��T�@�#�~l�p�x��s
�G�h�N%���������^r�=o~��j�F����<'b<���+�u�?� @G�I�Ez�eђ�x~ᝮ_ƣW|��qS�<����ԟfW�W�ώ�HMe���5�g"ϓ��Z����G���j�D��el�]Gh8*�;�' u��o�a(}ԥ9ĂM��繧�(p���Z���aLn�ѐ��|ۯ8|���x���`n�ְ�;7=0Gт�S|2�f�.Cq�h���*�U�V��?�M+�;�~_�38y\Hѻ��}��{�>��������7�oZ��h�1T� ���s��sW�fG�"���a�xˊ�e˽��������m�
%fD��a/q��V^DfL?�س(��G��%�\���ř������B�P�Ӿ��@I
6�O� y?l�7�?���t�������N�G��=+P��/M��/���=|�1��y�1,��=���O�v}g��� ��;��������q#�Jeo���$]W[��d\9��G	x;b���e&b������9�5CH����!���5�D:^m'��{NIq��fԊ?�r�G�rп��V.
��q��)k��'�X:����^􃶚�2O�����h? �&���|����}d��kI�K�ՙަL�`�~]pn�b�r)Ǟ�)����;q��6C����yb���Bk���K��2��<66v��&�����{2:{���
	��m�����gm�1��ǻ��Gl��ݲ���|���E �:�i�#TW1eN��-�|d/Ցr�L�=�E&��"����<� xc_hv_R�g����^�(���]&��kU�c*3��go<������}���xo�+f���Wz�)�"�̤�A�;����r�xvPZ$��m�3��,.o�H�{r�o��o�?�7�[�٬�����ґ�Z>U�5��q��p���$��r�h	>IO+��M�C�l�]������	��D��g�ixd�?��Q�����NL��0h�0D簰�Y(�z/�H{�@���F�\-��׳��
`���'3��>����^Y��p�"W�C��@���U�5�y��Uhp�J<}�ݫ��Y�����D�p�n=�β��[l"QM�(��unt�=��¾�>bm=Iv�K�EpG#�r9F>����F�g�=5wM<)�塁h�E��=+�����ϼd�,�'�Z;��R����[L+H�"�ȢzNV�槔$V)5_j Z�Cf���RX����y�#r�����%�+��'QF��,�|ok	���46$�i�(?��]	鞂���%m:�\M�^�LX�\����[״3|�����H�NE����#�#\5Y�[NZ`�X<��6��D���O(�\�X,t~��	ퟆ�Ϯ�idq #�G ������-��"X2=�k�b�~�A�-���)��m (���<�n/{��syxs(H�kb�m6�L�V�l���w`��O��w��;����h�#�����ܝRǺd�!�^�qU�R� �*�R�w��>��)�m?��@�QW3���� ������˄w0_�����ADS�c�|�^�#M�k�bTtRuY��������%���L�ou��0�[}��7{㴰Yƍ�|]��q1ay<c����d���C��lK>sHpՐ�Q4:�
����y@�)�fp�9xi��7�)���=ν:��D+��LO�͔�$��`�	l�Fp}e6�pm�؞u��E=����9aO�)]�dk�-�pϪ׬�{*���e��>���#������W.��q�ZȀ�c�',7��K+��w�/�fI�J�Y��H�#���dq���������g=����$�ڍ43���U��bBw덖�t�H�=q�Vc��3�:�R�e�ƧZ�7[9�{�pz��\+늕�mp.X<�|<��H1z&be��C̳������u��SL�W �1��e�T������3�k����D-�{����vƏn�$AM���g�/VA�|l)��!�ݼ�܊��:y��ڈ^�t6���dByf�߉�%�Y3���J�4H�
���'e�����s�q�F���в#�aD���_ؘ_���Bu��#ޚ��ZEe'�mK-k�������b��̰�qRG:`���.aOp��Ɩ!UF9��8������>]\�Ã��s�+��5N���g���bv��v�$MWb���N�סM�[tb�:�{K��K��@5�O�Q�Q�����o<��(V�A��������쓛H6Ӕ����|+�:	x�(U�b��X}��M�D��v�|񀕈�+U���M(1Bv�h�	�.��Y]���-$Ds��=��~`�ER��D{����F�'�~���G�~Y�i�S��0uG:�4ʠ6" .���T���@ږ�_?�&�Y���G�O�v�,5NjD~�X�c��i+nN)���g���v#P��7��]�(���q��8�bK�V-�o��X�噼��5c	�$�V�L5���Q!���2$�8tO~m<88cKꤘ˄R��v������0�lj[���K����:Zf�����V[�}_�s��~'�4�_�l�Iט��}��l��MRf���ܵ4�Q���B��4�D��$x����t�"�v:��>�#�C"ԃ�e)���_�ܴE����pO��ƍ���S�/�j�_�-�v#���W&�>�TMidY�'UU���>߶��Iy�*]a�S+���j�v���kM�
n�Ճ���{�B������]��;���,�?�c_*��3!C��8�p�̨M����6T��H��T����ӛG~�p�us��EF�1%�a�v���cJl�W�ږՃ�r�=ל'���FY0*t|���������}�o�\Nog@Zk{��e�@���ພ��I�2��8�Ue�Z��L}Ҹ���"���٦�?��w���(D���g�;�������8/�*��6�v1�+��¯,��0��6 Vb"�#$�����y9(�qH��v{��iTG�3��2���7�]��z�S�C{�$36	AQ'N��4���Vӕ	�X�c��h�R���D�EjrڴhYk9ZJp��]�§����B�XX���ưiͬ��"bw0�@�҄(ŕ�Cq���^a+_%[Tޞ�����u={���0��\�M���(��������,��Cn'���:�?_���|v���"�`���T�1������.��wmO�l��`S	{-��*����S["��7.I�q���跠Z��^�]���㿊C��2VA�&��D�Pç�s?�r`y3�m�̇U�n���`�)p׾n%��&�R�I�>������W�U����'�G�w����+�l��=`�A�:��,�G4يf?�Ǘ����p��(�xh�S� �Z��׺iN�8��v+�� e�J6۬���F\B�M$��酠�f6�}O�1���o�*�7�G��`��yڐM�>H�%�T��6;oG (p\�y�Ҳ$V��O� 8 ���b��ҶE;A�uTk!4=��^(f�ꆁn(� ��q�N��6�D�Q��iQ��CoXc�����:�L�؊��<�T��m��-�V��#zy23H��eeyY�x���;v�{��p�����CT^�u����ؐЍ0� ;<S.#a� �I�1��%�1u��a���m�jAI�M��u}��O;w�y�(R�R���~���Ũ�I���*�^��_��ĻfAfn��9Ц�C`������B����;i�ɖb#&�#�����QJO��Bּ�;!G�͹��1���y-]�F�d8M��V��C����dۖn����N�N]�����r������-x���%��н�m�f�����Ya���N:�-9bS���nd9</�]̨7�E�}ױ���(�,W�;�2 Пz�x�[8��1��K����~�I����k��-�3�_	��.��Ϋ²Ϲ}���KI��D��-c&�@,��H��M��������>���
$r���J=#v� �ΌZ���sY^5�l��U: PWۓ)A�F��1A^��u�c.3��"4�EF�DϮ��7�[�3+��)�}qK�F��F� �[5r��,���HK�ɡD��\��?��3���{:��GӚ:Ω	w,'��q�	��"zp7{h�FF�6Ryt��0쟁�W���A���J��bc�� �aM���m{U#}cqIEL�)(d�k�ٯM�{�`��jZHO����W�e���t3&�gH��z*/ó�-�[o>6���i�iYY-T�*Q�	�y�Zr�]��1NCJ����u2���qn���|�_���D�c�d�sN/���E�pCA2�2W2�_f͗ô�KK�,t-��1�L���٤�1/8�}�H	� t���!�K+p=AN1��$ըUף��G)��ʦ�Z�n�wa�$-��
��=t.�UʡU��@��)U����M�b��b!�ŕ���<��b2L�  ��I�z��������2�f$0<$�
bF�h���:��T��vt���V�9��p����;�6�/��Z�����=t�&���u��L"J<��`ԳD2	���:�.�������iq��%���(�[=��u�1�bu�1�-q��M�-�?�ᤄ&֥=7���;���;�t�:;<��ֵ+�L&^gR�vSa���ٴ-k�hÝy�4�� 񼸣]�d��W����M��wS��|������jĳN�t�|�ORӳ�IK��-�Z�"�t�j�P����mF�<��T�
Dݎ)��ϖ ��R��蠐0GDq/�[O��.-�8́��ᣰ�V$�p�14��7*���W����"r��Vf��&z lhxc�s�3�D/Ϋ��3A�L<䮻ctwfx�s�S�vA�����\|�3���[�L���+�Ii�D3+�wZO������0������G;/��#p�����[;���_�4��:�w�9�5<�)B�,jC|�����~R�,R������öwkq2zG�yF��eX��h](��6�)��RC����H˳������*��}�g���Mh��l��C� ֖�6�si���x�@������Y&�e����ه�bҏ���j�<�w+��K�v��Ւ��C����*S���}.JWp;5K+�aV���1��`�;�`3T�Ba+�����{��T,�M/&L�$��`X�!�D�o�j��[6z��>Ԛʹw�m5. i���s�A�k�B��]����&�dBs�&gMt���9�����!B��v�xr2�JF$#V�d����cث�>��%��`Q
#t�_?�x�u����+����-a�s���1���;C��m|RY�ᮞ_7���c��n�{M�Ujʄv�WXԭW���F{h�)��4��r9+w)�V8i7����3�4����,5D��)�e���S��LP��uo%xq�k9���[*n9��h���A��J������]�ɣzY�W5*�,j� ��*^�kI|C"�1�4I��Գ�!pE���Q��0��G�@7�rؑG�����1?�E�
gC�����+�d֌��~�:��7�vV�I~y���e�U�������U[��
Wp��"���c�xߣ�2'��;�W��[2!��c_Խ��=~�R��[��c.z Jb�
#e������~[���t�5=���~Z�T%yZ�Rr�2gZh�{6rg���++���W�?T���o��_�V�����i���u�aַ9FB�T��d�~��/"3R喚H�R�~�z���(!l>�Y^���\?>�b���C��nգ�j.�cO���ӣ��{5Z�O���������b#̠N�i�<�ՃZ����� p�2�H�)|��O4I�X�:X�,_D0��]$�$�P6l�3Yr���Q�;�{�����fq��~���<���DAZ!��H��ᩴ�(����&���RC�'�xiwߺP�fnܫ�����7�d����FDo�d��X�q~<=� ���.].�#��n�g2ʬ����Oe1[Z��f6c`�0P(c���r��s^k@˵�A��l?���J��;�R�Z�8y�ʕ\Fx�0��q�I�U^�(�b�
7����$�Pv�W���#iN�+Q���ͦ�8�qy�<4���Pc�CEc��=<���Ԭҝ���p��&��L�#���3:{!��T"��"^O|,���L;JC�Įz̃��2\[�\q��Va��J�6$���J��X 5@�TWo��¹ f�{�
:1U�/u�v�`$�~��Ay�P7MÔ�0�\%K\M�y�����O��>�.=E#���hmJ>N��uA��-f?�o2F�#f^HgH,�*w�	�D� ��+:��.v�r�\B�霳��p��d#���iFd�L�Hƹ�L���uڌ^���# �Ӟ�`�ꛮ�;��_�Rш:ʵ��v'��4'm�C�����fطuE:H��	;	���'�ʏϹ�o��BBG>|�S��X�TP��5��3�tcG�.Ű�n�~�ό��Ҽ��^����<���Y��2S���_I6N�n\�"�'�e�<V`X��L_@��p�g�����jS�!0&)P�S��|-k&������*ɮ�l�d���Ѿk�3��r�mi�\5%�}^�8�Ia�6��'}D]uq�P�gd*�xʁ�䅐�Pmvq��+�<�_��=S�������>�]���;�m�:2�籕lj[��;�^�sڱ��T�p֩o�<���:e���]⤶Pj�x	��3ˤKyq���D6��k��N֮�"���V�hl�D�u�L�9Cc��[�K�%��K>8����dIS���`��R}2��i�9u���w��3R$?h�}�PU��wn3�yP�*a�Cxt"B��s��"�ͪ1�*��7�H�׵�$�u-q�d&���8��b��J�QL`�Xٚ��榚�q�5�n' >��������3��KW*�z�m)�������dI� + �����-�:���}�\�,^-���S� ���V;�L�\!Ki���}�W���.��AnJ|��	`�n�e�c[�u9���1R+L��Fxj�ObH��ɧ/!PVI��V��i\�����OfDS�0�z"u�i��(U��KP��P�%&������	w��{�����c���������QK��5+@�x�
3!����[�f�III�#��xẝ"�� �`M_��I�}5 %��f��bT��{ʬ��-��eCW�����|��>׎�����`�{��DiT;���P�A����y7�^w+�������;�@H3��&{p�0e0����q2J����<�N||�YϺ�����w��m�2��
W{N3��/�X8u:�p�T���g� �����l���<c�K�#h����J��;_��j0�t\[g�r�M��
/�[���v�p �Ŷ��=�"d�1]��*	k[��-�^�s��B3�.��X������r�r�&�[Hd�L�-h���n*��������J{�-�r�[?O�Uq#S��g�om��R_Gʶ�����l��2���cX鏜��]�� ���7��$`91X7���p���P.����i��� �,2�3S���x�'�ٞs!_�v&|��L�Z9x�|W���@�")`��v�t�fZ�L����ޢ����UH1V����7����m��V+����N�D�G���}�_���2��)f�'�k	+*a��K���L�V�`�wX[�kYB�)W����Q[�ߩ�둇o����WL"Y�a�Y���4��
)!ң�`����
�;��7�Xa�;\�@ X����JL�+pb
��Z�)��3r�A(0��n������"sf���l��n��n�u��t�>qf׉v@V���lDe��n�.\�������\�ʁZ��}�?ctYR���Rv���Ͻ%���a�-]
��wʥ$j�`����,L��^��<��L��b�/���w��+�����֟T�^��y~��kOk	<�z[#�ݔd�-%�ǧ�٣_5�C�IM":�)P6g��$`/O���������X���Ӷ�{4:�k��L6�}x%�S�P�UT��9�'�wK�>�s���]�B�͹���Չ���P�E,������>+b��`��@-Rn�j˭�!��ړ�D��?-^�`�#Ѻt��������Ѩ�;���BW��U��P���RW/������ɶ�u�;m����~�$���#���CG�ǐT,E0m�D3��R�M�6���K�ֳ����4U-�&�	=A�:;#P�7d|%z�:�m����e�tt�es�K�!´/CY����0w��ii	vͲn�JBl����s�D&�G��i8_wz(�Oq�	��v�� ���R&٢ vɦ*qph�d��d�����mr�ɔG�(o�[PJ�`�*�at�i����G�@L�QǯQ�&�cuQP��[~�4W]U�&M�rPά�H+�eMM׺�b��&\� ��t ��}�As/�DK���ie�@u�b��ܩ94�N��b5�C���|3�}}�bt�i����3vl~��=Ѻ���!����e�Vȯ.��_��&f]�4���{U���5[�鳠',{!�x�:�HQ7�.����^P>Y�̓W	��E��	�USb�SL��7�C(IS�cfy�؟1:@,�!;� q�g�,K30���1CL���k;FR�
f�q��'F]ή�L��v��J��K���$7�z��Z��u�X�(��� ��^WC`�����A�Ŕ���M�t�d�HfȎR<Y�@qC��5Lg��Dd�\3ڔ�r�D`#4�����$D��\ek��娡���L_��|e�'Rd��<\+�6�!Do^�1�]��%��L�ּ��k?�37��M�X��>�����ؤ�O�t4��1v���v��0�Hﹻ��MY�H� ������D�`����V1�(�����ÌzT�{M�����_�T5�z����yW��Q��(.C��v�c�� H��P?:�9yWH���X�|	��Mb�CB�vͯ�C ����(# fxHO`Dޞ����[g4�e�h�m�����҇�#�uW|�N�������vL�9�L������Th�Zq�6�U�Ӛ���	�<���$:�c˺�[�])<�sR0�N`�04Z��ٱ/��0��H��F�>s�-�+��<�8 wB�?m��wr�ã���^�ۛ>I3����U����g���1�A�Wr�=n4��ޜ��δc�p�m�ǋ0���)�	���P[<��RX�e1�̽w�L;L�ijt��[��U����������ӝq�:�q��2���$v�Mf_ךK�ˢ :T�H�2�f���s<"��DLa~b@E���Pùx�m�M��"2��M��4����Fd���K���\��:(���T�j@����n��0�:��%�_\��7��޲S`4��bī��"�����H�\�(��	L�=2��9��)v�4�Q��hΚ�-qiY��K�E��e�ؼ����A��ÿϸ�zM�*7���)�g�z����P<�E����	s�M�mSW�=���8\�L����g(�)��2�+����U��C�_�P�h���{��(C���k��fZ�o�Ak^���:����q�ٕ_ ���ul�KP��6�z��-�5������(4X�n��R�OY��O���G��B���$.a醘J��ИB	�/D�z�O�ɉ��{}�Y�ѵ@�Vdf�nƳ�x$.�0�0�w���dc��:�]�&��ҩF�^�R�_ݝeq�����f�]���4�����r�W�τA�8.�J`]G�-<��T��㢉�LE9so�����ʌo3[S^�[Sdt��4���n!s�(\�
��P:�bvG˰(� �l.������b���Qi��KD�CsAa~�y�u���7���4�IL�/�����,�3T��ѱՕ�i�_%�'����h�z�Y$�l�Sy�D|���N�h���lH��XЋ�QƆ�kߜ;�?Q���=��	�4��I�L�}zJ�6Ck)�QƦR�����n?w�����$�g�vT�v��ʷ�G��鮦IJI����7F'Xs�t��b�Ų!)������?�P{]���	.������&.q�?��&S���j�W<m$=)��pf4���(��G��,�i4҃.�Ό'u*�=�r%~~;B�S6(��	�����9TKS0��9D�EAv\��L�ً��9�0��[��~�u�!��Z�0����#�T�Y��z^���o��[l8�R���|ᜥ�qp�7ׄ�!ȓ�W���Ǚ:���r�Ήq��u&_*pq\Yd�?�*��3�ket9�1������T9"�2�� /@п���xlWb�������'�؊xȧ�~�|�����������%�6��L% ���(J�t7ڐ�;zЈD3Yl�����Pq�ӟz��\����J�3T�}��������ײR��}��r�Qh�$&=���l������˿�B��k	�0H�g��-�z���Ať$e�嗚Ȏ���(��uH����g.@�^���N;�D���L����i�'K�i��˱v��&u�ܞ�Z�TΞh���.IE(�X��X�Dao	�*iXrxJɑf�Fq��M:/��nd+mS�U�0�d���Xb���,��R#�MWu��f*�Ԅ6��o�ȉUcvK��*�.g	[�[tz��0J��=��b`��,�y�(1���vm��(�e���]D�Vˁ�*]z0F�|��0�s���bco	�%c��b��Y�%lJ�V��dg�p�R�e�%AB�G�5��pVKψ��R&0���j��:#_`� ��g�>@
#Ζ�1���������z��N$,`
���c`L�D�4/c�H����"P�F^V��H�'?�Uv�O��|��e�1wU�g��HX�)r�K����1S,�K�����zb�B�ݡ DQ}LE�����#<f,���*\�������`��n�bCH��{���+�p14*��1\�1[��F���2-wJz=A��(�ʅ����锧s)��o�Q;;��J.I:��,�C�C��ʴ�+�#e� ��@ ��4�9� �,0R�Q����V�Yt�Xi�%'_:��U�k1���X
ɑXeŭ��P6�u���R�F���l�^e�N!�K ��W���eIؑ��˴�ZN,�X*͔���O��M �)��΅�U#���@��s;���8�s�?^�F�����fw3? �<�ڹ���ߟ�� 7��nݦR���Zq~u���*GV|e�w喾�5�)���yUQ�%ӑ�d��
v����`�P"�jZ����p����)w ����Z�vZ^���Ei��I�V��:�p^��'m���R傰'�8��)=��翍��m�:/�=LOPz;*��8J@D�m�"Y�e�@��TB�ƪ�; #��K�V������V��`ieB!��#=%��!E, ������ږ �#89>:���T�9�����6ܹ��p�O������/�6�WgW�;�[_u��/���{� <��t6��5�b��H�a9PD6V;�ШXH�,��c���)��H�XT	��I�1 X%\�[�O��K�
�\�%��×}�= LJþRB�ɼ,�5��Db��`��88���nu9� ˾p�}RzFbږ� "}F��(��@o�3�Y����q��+^2�#*̔�S��q��$E 1�[*7�zN��F�1f�dl��E�"=q%O�>?^�tc��R��^��7W~�P���ڂg�;/hF�FFו�q��m�ȑ�,�YdE!P1��5�i�,������.G�^�6	
<�� �F�W�	�Tu�x���^�����LL���H0��*�(+��싖EhY� �-��q���U<�F�œo;��-��c�1f�ҳڕ?���V��tF^Vc5��H˓c;ʪ�Π��4#� ��n���@<��?[��$��Qt�J�!.���>�ƿ6N)�KPq�n�k/��R�wp4����W�,uDP�EL��bER��j��a�3_�Bb�,Y5��!�-J#m�/XM%o���'#�b	R8#�|��YV\�JOKaZ�CS���G]��Y#�ʁ �Rmd'��dd3ax�J�����v��0�if�|0�`�Id�}-#|F`"m��#��ޑ���C}�ު��:^�F=�;*"����ι�ﱹ����S*�� �R���wTt�( �P�5��MK@>�	Q�qm��08�~:{H���S�����z�I�W
�@h#BBg�)[����3�Y ��Nad�KmE�U��<;d%O�FP�g��)k����21&�<-���H r0A��ޒ� �
�r�K����/S��L�q�\Ez���{iv]+�J!Z�H�QՋa�e���{��Vٹ���(�a�Y��|��\t��t07�{f��^�U�Q^$�RzQ�a�[�Qv�����4]<�.(��苆�� V�qқVWM�^�xN�aۗ_~�����#t��o���ZL)D�] cK�k��;�;�óØ��d�0*�o�k���}�sI�gd�'tG������ߛ�=��9��MK�G�FS?����!w��g>�ט��������8
��l���,<\(�@>|�EV�z��o߾�����!�
t!�K9\�;ߔ-���ЫΔ�&�W�%��0-I��E��,��ȍVY����e_����枛�h��ٍ��DQ]�3���,��Ő#���,�1rSz�u��(�=V�0�+P��v��Ȝxn��3�K�:lu�L
����F)V##�B:p���M&8)���Y�Rj��Oo*y��N�t"xc�UJ��u�H���b1x���8_8bp��a�q 0���2��B>����?��S�F9 ��2=���q�_��_��"|����~��$~����a�0�|\��U-`�'��w��\]����l��}�����>X[H-�+g������W���G}$=�[�ɞ���f¤`Ih�cO�-��R����tMT�
)�0�T�>�IS�F
�G*���������U�2�Y  ��Q=~-+"w�u��$�����K�ci8N� uT�M&%#;ZK�X0#�X 7�
��c��Ɉ!���:�F�I���%c	P$`��CU c��0x4���*�m
I�����i�)b9@!㌇#
Ř2�>Z��u	�zQQ���L) 89���)�;�X^����6�-�(}P>���x	g�%���x���0� [�I����K�@�U-FHK�Ppˑ�U�y��f�Ka'uƔ{G��ml�ގ�!�+" �*.E[�Љ(�1����a�&`vxK��A�ˈ�;����D�(�jd�alՔ����_ �����rT# G#*I�	Ƒ}q>*�h��3J��ȅc�.�`�;�YJ�ղʈ����r��b�I��i.S���RqUa��	�UyZ��^��S2�����;GƕU�$)��N�ƫ>й$Y�\�˭�<��`�o��(��RW0/%.�r�o\(0�j�2G����i����0���Q��tx�'zUr�X�JY� �E!u���@	c��ё�2]m�',V)�ڨ+�V�g�`�F�U��f
�9X"eb�4�yx%ʋ#dW	!�ԱY���@�,)H������p,m#Z@��\���do	��FF����}.��J le�Rn�!�t�F��x�Ed�3a1�����d���>p|����G��Ϯ���-�C���x�{���j�|^���Z����m{d��5���OϿ}暈��ý����՞��Z�S�ë�d��e�Q�PzUD' �jU�]&�'HL��L��m����B��)*J.t��Y�R
d�,��@������a�,�]6�QL1��Vɟ������(��%9��������O���;V�.�>�2^\^y�9`����Qh�+:LF�BH�sG!V�W� �r���b�ت%
�
a/��K͑@��R�s/$`	�،�F03%�%b���犸����p�`o�����vn�}�����1oo�(y�3v��9w�7v�������ë���]\:�蠝_��_��;�#'Y͠r�.ѱI�Ԫ�P�<1ӭV>;���H��x �)H��m�*�����U]�j���Νй,�tx�ؕ�RP�e�U���C�f���� ��V�⅑�@��{��7��#�[��r�C�y!�Vċ@�R"4�n����] Q��X�����E�T,{���ưʧ������ZBH�2M�TJ��n��i.�@
�(b:%{���U-�Yxy����w>Ws��|_&{��[`4�CC������F��{�Os{�*�b�	�%qKI	Q�	�՘��j�#,F
�'� E�Uu��(���<�ew��Y�q���(4K:@1Y%�k
�@�ޞ���hZi�-A
Ԓ�J{Y�YJҔ���p�������J M��%4_٢*#r��` Y�Hb�����sȊe�ĝ蒩��U���F^��b,�r��!6��K��Z��jQ!��8*p-%�AKG��� J�5�B�}�K)�U�C����]Ԡ�;���K$�n����nov�~���}w:>Y��\ ���R�hcU�3ҥS'C���8����` ���9
Ge		L����%��j/rF9`��O0��sg�����-L� #�$R�|�����J(�4�Q`��,�T�e���N(�V���Q�%iu)��
@1Z=�]��H�v�
̅��$=# <Z.t͉���v#���Ht���{�`�������2�lL�ƥ)]��^-�(Ev۶c���ݷ�?���B����*��cG�el���R�+MBC�$���R�� �=vD��0[V܅�/�R�Î�#�bQ�Y�:LT�A��bȅ=��CS�7 �|��?���^�x�"`Ɂ����"T,���5�!^	;�|,I��M���S�eYUp�0JzF�s$���߼y��>���BH@gʁ/Ū$1X��T�MCZ��Qy%�`A�x�u��/�˗��=����9�n�m���#�p,�L�!z=�=����b��.���4
}~6����-+G�<a���7kd"�U?"�n*.w�0�C�^V	*��tM�����ן|�I��ȥ��z��{�qL[*������UF�]m�C��������O�$�<=����b�yI�`/�x8����+¾�<���o���1}V���C���r�*w}~q���g�}��<��@:_W}&ڹ�����z�9x^fz���U�*li�������]L���K{@[��S���h��2r|x���n�s�-����uCܵ8b��%.�ڞŔ�%�[2�a [�td��)A��T�`)Y��˜K�����eb$,!9���M�`�T��)ekT���[e��pE�ti�wi�gTf��Ħ�Qq'�9´jdq���&+-傁�V�0��U��l ����`�r65"�^���W̦	f/�|�m*?�������Hp��V��a�K�����}((Oּv�'�]� -!|�����j��AS'�&��#O���?��U��a�7T���O?�T�ڣS�M��ۿ����S<�=su�;_t���>��B�~�����*��<������������/���k��CW,,���S���Q$�Bec�`�(�kЫW��������:�?�r��VPpo$������_��:^��8T؊�;8��x��_���j�`,}/P�a�ܒ��U'풷ʱ�X4���vY��;iw<�Z,�-�����Ȣ
F�� J����gW����`��0���)�O�����|����pQ��m�j��_p[]YYB���)��¾2)tKUo	�������n,
fb��h5Y�08m0�l{�q�Ql��P?Y�?KⲘ�V�D���/�����,/0�VELK�F:/�8��9�D���8��d/�)�L���	:f`b	mF���fZ����%N��)�!ˡ�4Ŕp�kD��3@�� ��8��EX��d��oH����LkȒ)m�9�X*�r�10cq�m`�21�v��g!���5��O���YI��JΥ��Ё�w�d�ŒZ*�W'������)63*z �a,$8-��B\My�K�Һ��h��%ʫL� 1���O��a�Z��C�W�v+Gm����v|c��|�׶.�]�x�m�m߽�#g˓��;~�[�S��q~�+�S)�чMg�s���Q�ܴ�n����
FQ�]F�]Ī*��a貍d���Oa�Y��g��{�!	��Xє�=YE�-����"Uⵘ/�!)%l|��Y���09���4�I�)��S9��L�EJ(mk��͌�4���`j��F�lJ�G��|:Ju`�mK��i_xlvt|����f{u|t�Gh'�Y��v��ɡ�=��w������=9:���:>�{txs���b<_���ہ��uy�ծ�����x&qvq��w�Όw����g���[?�8���:��z�X���f�K�^v��#I���R�d��߇�}�pݨ|���FzS2;:�_�M;���tL)�"��ԑ�fK�E��Ʊs0��j�[��|�dW�7A6/�$]a��6�>ԏף]7]`uiw��������|�����o��{���.|����:��=����滋�;��|_�狺���-_=����e�\f��d8������lu�(��R ��Q�v򚪠f�󚋓W7��) �u����0��o����I` �9�U�;w�i����`\[<1>��<9�;���=��$����}�ϫ����vs����;^v�|���z{�x�����w����y^����ړ�wgW�|w��޹����ڱ�������Ӯ��f�3¸���$sF����fT��8�!��Z��졥��QZ�Sl3#�.�0���ҵ+�Q���{x���GW�9IM�1 #���>~S'�с���:.���g��?�/|c'�Wv����v��h�q��S9�}��v�@�K�w������fg����O�w��w~5;^b���q0�_��3w3v��Ji[Q���9`9_&R,��O;��JU�V�������`�FR���Xj,;�<��3��X� 3�;��5u�7\��Pn���|]�w������<�h���h����������_�E��g���>��ty�����չ��m��M���>���w��N�=���	�u��q�\��n̛���Q���n�Zl�BUUA�@�M��՛L7ҽ�TS��+�h�v=���3"=��(��**7�<6T,���#� ccvziP0��D�./��8�j�@G��sЕ��E�K�,k\��h'��Ͻ�y�f�{�|�};��g�|SE:�z��{�k���Ƿ���{���i-�O��f,�Ny����M��M���ZbA�%�z�š�2�C�g3��l�,�<�� �0�܍a��;薜k�wF�O�bi���\���S7���w^3���}'��j��R�7w�Zks:co�u��������������ߜ�����������n叫�=�Bd��?71�P�3w�2^���?~��>/�jI���(�����f��PQ�'��4���Xhuϖ��*`XК�7�y6m���N���US:w�
QVHH�Ԏu�9�����ǔ����0-6__��o����������vo��K/��t��}�Jo�N��8�獍�32�s��q��J)%,yK��F�Z�,q�"t�8N���,����Pǥs^�L��gә丌;"�/�^��=�����9��&[�FS#G)���s/Q�n��g�j�8���o����m��s�*l�+#�����r�3�<���ց�r��==9���d�n��?�"�j�}̳c�72�X*Wi��wVd8=^��y�Wi�o����������_�v���d�		Y-��)z2��T�`��z =���2/:i5w����B��S�b�<�m��w�mF�����m����q�P>|w
����!�3ڈ�E�#9=?󊇍>.�h}�����?U�($ϙؾ���f��֥~���,���C8�mq*c{�ʏ55���/����&�M@�@�>\HM	��%z����s�1�X%�X�,�B�$���aՉ��8k^�x��~r4���8�q7b���w_.,�f�������0�½W�w���ޝ�D8�7���d������1ՙ�>����]��=�3_�?���� ���붻�ch��ԣ4_g1���K��m;w��jP�8ܷ�͵�    IDATn�{�y�S��+�K�8����!ڨ(�tl$���\�:�a��aH����Q�$TJ�ƒ'(6���#�ޒɷ���G��[���\팿C���]�2���n�!�;�%F�w�׾����w�=�<=����+L^PO��[a�8m8�?8tQ�Igk��o���l�h�_~�3��i��jFv=��@�]C�|�|@bh�z�|HʹD��F�!M��|���v���F0	h��$Pn�|��--���2�[����Y/`b*t�%Д��	�)��3BZ���h���'sY�s4�)��L���c̒QFQ(�N1��C2�ҳ�x�a�A�\ڐ�+�0x꒔�f7���2�J\��C$��E����H۔`�O	#y�*�����G��E���g�BC{���Tto�S6O�� '8+!<6�#��k/B�@9wO����?		~���<#�*_;'��իW�v;_x�T��ْ睟|�Q9����|}��wٚ:4NA�¸��_�B	�W"D�.m�:��^2�hܖ� GNDo߾�c�����ABV��NH��)?�ݳ��E<�$�B� �k�רf���2����BDi�Km
������*(*#w�TU,� ��8�U�2w�eJG%�t.D:(Fћ
�b
�%1UlH$�)�m���L�[�|�a�o�p�FQ���\������d�E #;������b$����TbF���� C���,��p�y����LJ%���&�e1%0���Ud*(;0;}Q醄���ՙ��|����Y(����Α��!��u�����L"��v�Q!q�Da���FXzV����Lv�TP�d�H�%i	'6� �.CS^�P ����x�QJ)����ii1�0�7��9/�(���n �ܪ��Y��q2� �9���y�r��F0nj_�0��ˇ@�c����,�pw��#�	)I!�0����\J/Z �̴c
F�Rv�,�)ME�cK����t.�B�L�n�n���<���X%vu�F.2g�S8�kW���xHץ�X>���&�!q�V[�Y'T/���B���Y�`�|�$lJ,��>��l#OF.������=�����o��V�9?���v�Sn���ᆦ��W�zt}w�~���<6�i��w�v��򄗬��N��j����B[2J���­�뛜UJ'|�b�"��1K�P S�F]�L�2:;����k�6���i�� \i��1~!(�F�\�)u>��|�fDh���[⒘��h��H�(�{y��� �y��P�	:��V!	��+��u����.��mj$L Κc�s�5:�)}���S�I�v�۽;�>������{ϟ>{z��'� �?r���౅��ys{ხܮ��x&����'��g���y���o<Ѽ�<=|vq�q����s��/.}B�����P��m3nZ��[�n���6����IO�f�
X�PiGD-dVw��Vx�� #��SF���q��uV5ْ�g�c��CJ�'����WzH�'G�o���%����Sg|�bn`w̏���|������k#�N��x�<N/g����w��}��������O�s�`l���g�;}���w�/n�5��)�����۫wW��{u�J��Y�վ6�:���������婾�r�B�m��:U��&�U 
����(G�!�5PK���h����9�)/K�1t0�th�����cˌk����/�w�nww�yr��ٸ�����xo��������]�̚//{�<6�_m��J\{�����̏&�ߍ�qyq��Ľ��뭟�^�c˛ӓ;�n�����7�7�����#��h���}|���q�wӔ ��1�T؁�]��*@�J�d��cZCP��|�[jʅB-1��%i���+�̡����gg�[��m�kGϟ=>�w=L�ҟqwl������=_��PA�]��������}EH��������g'�矝����~{�su{6^���R�ɼ`�?��^�f�nv�rk{0>�!Q,�Hu)U�1�&+�ޒ3�E^jbo�1LO��=�U�u��UF�B�����V!�A3�����_����vo��p��{��gǇ�N�8��&�6����./��ѝ�5������vǫ���6��؀�5Z}���{r>�ӿ���+��o.�]���r�*����r����d<`�z��G>���Ui�Q��j1(�]颒�\�� �L S,qOg�%##��Ύ�n�D�1;_ ���1w�ܵ�n	�;ד��Gz����WC_(�V���s��]������G���mwn/��ɱm.��:������7�q��h�O�z�9?<q��<��88��][�N��9.�G�^
�*��n8�K�҃��2WCXj]Ū�BxY�euD��_�x��DE�غ�E��?^��__`�
6v�j$�k��2�3�a�o�jj�G�.27*��~�>�{���d\K���Ã��=O�������A��xw鱎�2��/ky�a���'㙰�~}5�:qs������ͷ�/�_m�>���(�������&�ى���p�'u)�g8��(V�қ������ �)��e1�*{�j� N�������Q�ДC-�(/��A���q�g��8�R�4��]]���v?�a��G�ώN��>�m7���1������vs(��q֍����w�1r��m��\�߾�ն���#GA��R��ȁ���8MP�[	W/��jK�Ȝ�Q3���zp��~�ӣ�i\F~�g�#(�,|�8D��Fb�^�ۑ?��Oܑ���O �@���<]�	��qE�؋"�v������;�7ܾ��o.�Nu֮���W�%����c��v���7�\��������������#L�4������7�{*�'�'�����;�����ȧBg�ϖ�F�f�_�
���?���d�$Ei;�ƾ,���S�(�:��t���8��&=|IGR+,�p|�������k7H%�1�����=��١����~��7_}��܀�l=�;��8ǅ�%�KI�x���K�>��8�]��n\���5��`�=�R�k)���&1��+��^�
F^ȉ�)�E�\Pa`T�pL*9c����ޒ@���F$1 ���Ό�󮲠��F�˗/���sF�^R��}R�ܙt훔��8/~�+P#s|߽?��~����#���o(�@g ^dǽb��z�����<�l��:����{O�w�`�뎧��|
}���;�����%EJ��(��)�:�\�
'|��ŋ�>�IǨ]�IH��Աj��� 1jTKg��ᢰp!u���a�@́�'��9���
KQ���Q㲷�s�/8x��/���0^��柖)��z�'��x��_������՞qz[���+���'6������G�|}tx�=pY�?<�zxt����� <}v����Q{.����%[ߕP��S�T�#�y�H �����Q���MEFw�1j���-;K�#9;/�AN���U���x!t�!*^�-q���I������P�tv�W��F̌J+.�ȭ��$�;N�x��J`��gU��@F�,\X\X����#w���bd�3�4��4�hD�j.������MmN��Cl�SV�Bh�C���Y��X����Q�Xj��� 
��/(0�qv�X]cI<�0v�h�=&t��RH>n�X���
�(w\�ӎ�����ʑ��r���Tz���ؔ`?�ę�*�7o�8X����G�m'9 �Ez^[_�~�1�6/�����
�֣P�%�9�dX���ኦ`�z*�?�я@�%�/()RT\�z��1,O�K�E���}H޾}���ɒD��c��O*�Y$���?��?S�����*Rs�T����?����=�q��wKV������@�Eβ���7��%�M�Z���mtSBa$M-%���@**Xx���J�Ti� ���h��$�R*����|q�4"�� ��X��/
�=T�� � �)-{BgGbj��^��Ei�{9dO/m����6;JH�J�q���F�C�,�xL�yf�e��X,
c�IeƦ���U�GR+(xH�H`Xt�1
_K�X�l5��%�� �Ѫi��ğ�H���0Œ�U�5^�r7r1���BL�P�Q�)V!�ƥS����,�`� b�ܳ��5-b�H��p��,��0t:�U��FSW����t8� `�hy`9C:L�R��t�����]�#�|��jq�-��NY9�b��Np
�K�e�,���9��4S"�4����(4c�1E+h��ۖ�Z����(GHv� �Q���Uz<���)��k�%�r��U��p���E,�Yz9�L	`p��OO�gӌ�齪g��'��n�z�.����Џ�@���9�O�I깒����k?�;p�WD�ːK��%�(vJ��v&s���T-V���v�)��B�alψ�Ѫ% ���,a� E����^;pv��T�e�BP����|�6Kcq�-�L�L����dq�!W�)�6��������h	�V!�,����%_�0���F:��d��￹[�^,�,
	6�w�j{���3��_�v��x���c�"����<������x����乯ۻ*�l}�����;���C_�W��)�g	#m�v=:��������/����?�z������շ�����<��;���o�]���h�K�f����?����8�]O潡�1�t�}�:���QQ�����|Us!�`����2/�0FF# /��>��R܎H <V�)w�xI�杛;�z�B5t_<t�v|�����?�������{7������k��i�෰w���gwg�����l�wv}�����oN�����_QuM{��x�����;��-�Ý�G�n�޽?��C�۹9��9=��y�]���C��Af����+j]��@��ZQ�L��	Y` �,|K96B��E�VgG= θz +KF�����3�ڷn��x���x�{Ͽ��z'q|�qkU?=������O�����<�;������AC�����nؕR�����w�m�O��O?��<���������S?���;���g�:���}������W�}{��%�/�uC�n��TQz�P�M�rV+�Uz�RBRx�z�V5�r�Q�V-��9�X�"��sDI���*E���	s|�7�����m����?����{��T�Ǿf�2r�����ON�<~�������f�����nǕ��ru�=r%ǽ�k�Z��z�N�p8�µl������?�C�����l�43�&{��}{~y�d=`'###"#"��9��߈3�N�\�M��8�4_������]g=�.������~�V�XY^�«�鍔3��Z�����ye<��VT�}z_xH�Y'0F�$2�qTxũ�m=���yg�R���<!:�:2Vh�Y�K0��\��ltm7��~�9�6w;�tz�0?���ǲ����z�ݽ�����Iм}6&/k��녃�f�Y}tg��J���sS��P��ӝμ�3Z�φ�]��,Nu�g�+SO
�2�����J� VĢ��U�������=#��P_q]���:d�XГ Y��+=>� �+ "V,K�W�&���Bݒ �E_\�K{��,k���B]��*k���+�'��i��T�}�R�I_�Z��(��kl�nrc3���)��j�ܿrf�j9����ts3m����e�'��hi�����_�����V�Q�"E�+b5�i�h`�B	/b/��I�'�9�)N.	��x���5�I��RD��8���x�Hu��ZK��Uk�o�A�!�i7���rշS75r�݆��]���R�f�XW�e�f��,��Ŭl���E�^>\f{��Ѳ6�����v5��F��x����5&N7�q�q.�Sc�̉��P��]�%.�V_�4G&)N�d$ �K�0�������+�����B,M~�� 	�����ۘ�HƂ��*H�ʅ!�MAG���/ZUkn���^d�5X}��v����f��ŏk�z}=3s�	��5Eo��?N��Ʌ�'��|Q�.W��^��{�dtk��s|oh �},��8��Lq���R�X2fX�W����!�W��,�
\�>}'�e�� &*�I���9��H6a�#P�qWXHF& �а�C��3��l2M��/߿~�������|��h��c�I��=�j�&$4����6��lJ%&�W���||C�F�ȗ��r���3zf{����Z��p>�wr�����:�ї`X�AVT}f�
�N��+G����L������iΓ�u^#Y���G�P9����c0��o+.�R��%�9��5�lx�'2��Q[Q[ �"�χ�ht��]?~4�ze^�(�-�P��Bg���&�r���֫�K�m�-q6m�}|D��Ӄ�A쭦B˃��]���)���i��P)�uMGQ��FNL�`�Ac�c��ѨFzUu,�pJJ*E�.���	L�A���t2�D>�$C V�&�\Cͩ 2%��O��x���a�xu����k�U-G�!�ҿ�wY����UPe��hryy����Ls�ܚ����i�L�7b��v���5�M�k�G-�ni�����č��A���v��o�I�wx|082��%�}g�Z�<�ꊅդ[���iE�jv�O��sÍ���������qv�x$^d[��թ���b���}�W!.��=I��j�<yb�����OiEn%9�.V��G27뢝���L��_�3�\-r�O�f��s�%���(���uVC���E2VUݸe���u���ܦ�/S=���˲���[c���ݞ�u��փ�'{���(?�ʓ^�t� �-���l��М40M��7�c^v�uq8/!��[EK�	��-�H�*!^HY0���h�0��2rMG����b� ���'�}��7T閫/Oυ,�'W� Oh".�
GO����x��!F�K� r�X$��GL8}<9��B�#!&�9�����*��B�bB��eі����$�E/�^!�)B����x��8�Äx[#D�`$m�LT�[�Fg z�3�v�FC�rl1���q���oMaRF2^�y��uq����_����Or<�������KmO�S&�3@��g?��������jC��(A'#II2	�2կ�S�T�YD2<�,"Dl.�(�b��������)P�;&�����Fjt�o�� ���?��l��^��!��������E|Z�^e{9�?*�K���o�[�æ<e)Z���� ���b$yY �Z13�E�Qxے�#I^#D�qs��\ ����Р�$D�����xǊ�4��X�Hx�����+=�>Q&7\����
exY-��Tk���P\�� �.q��䐹�BV� )n[b�(�Q@$v@��V�d�۲ B�8�aWb��$+dQ)4��? �i(!�"�
0i�"\���J� ����#��f%Ş��A&�@5` Ĥ��E!�w4)4x1z�E\<���z	�����\H�$�qx%�F�&�d5 ��tfi( NA��b�UP��%��EI��L�Èa"Jn�C&&�L�,u
I�d �W�X��c;� �b�F��\0��"?d0`\�0 �.�o��r�D�V2���$���B1�?�'���P"V(9�ٲ(�� )YJ���L@�B�HYd�A�iɊ ��������-TA`x��Y���^E��d Yޠ���ǘ KR�rI�RZ��-��JTHY�j�ڲ�*��8�lЩ�57>*�&4�YN�ZF.��>ݨw'��{�E�Ѿ���ˁo�>	d%���r��YT��IFs�aG	)(Y��"0�aASi^b*1@��B�L�VJI�,:p�P�}xŴ�*�(	�`+��#A.�,p�VxC�MT�ą,�)����
\0������!+:�Ȓ�ɩhK@�r��n�b�d	Ar��%�����X��B�rQ��?kfw�u�	�/��4mG�;έ���>{��W��M#Q����c�R]*6����ڶj6�m�Y��� q}�o������׽��'��������W�~E�P�k    IDATތ��?�����������dvg���3�M��QJgiv�,H�R�U�FN+�W�ދO�T3%,�b��m�^ �I��dI&	)�,bC�8M  6��)�&�}�
 4@˿YOAms4�������ɽӣ�;e��cRy׉C534�-�1};�l���jNڑ1�M�`���c�9?�[w�釗W��޾��s2���n´e�6�����l�iX�ͬ��[����Y4�k�LqV�0i�1���m��0B��=I���9���U0,�m��dq�䦲 [���m�%���;���K�70gi��^9R��k��!�;n�;@�ɳ��㮏m�|����.��![�}:��4[ٴ�6:���w�cv���S�1�֖w����߼���b9�-O�7kӕ���Kc�Ʀ�N]*ۼ�ܕ#;�����\�x���]�V4�?OB�(F��[���.؛�3��$H�"F�[��\v�0��(o7�4`p����d�C)�G�}��3�^�ڶ_!�r�:6��eb�����9�i@ո����ߠ�(N�iy�)�Mv����m)�Ug5����lZ�r��|4���8��p3l�.+[7W��X���1����:���˥��?����^�O~�O�R��ܥ��O�plLM# ��,�����r��_"<�cQ&w�Or�^��4 ��DQU�zX�-غ\
X�d
�`�9�m��1��5>_5g6��'{p����������a��Y[wR�	/�2oW�-�?5hm��*�MS���������嵕������椽3�o��7���l�iu[VM��P���-#ťCH�Ǆ�瀷>���r��y�#	F��x@#c<�,,[A$ ���B|�B�C���&���d�yi�	D���m��C�5s��|k�Xڽ�/Pc������A������A����������IԚ.\�Z�\Z a��|��������x<wl�P;n�N�����z����7��{�ٲ*H�s�6����2�J��y�(m�:X���yۓ�u�ho�&�-&W����딯��{S�		/!�\�@�
L��â�DP9�����k���&l�7gl�{�^��:<�z�W�S�G�j)���u�v5���s��'�����ϗ#�����h�^��h<=�Gs�L�Ѽ�~�iڹ��(�������+-Ly�X� N�ULC��ifL-@��	�`#"�� W�8� P�<,$H�K�D	��Ó@#PI��Cb1�`x���ώ���M���?m?0�ܪ[�k�͚YGߊ���ǋ�i��v4Q*�sf���׍���dc(�#51_�+��!�/��m�}7v�|m��ʞ--G3󜖖i�l�3���ʷqX`[� ri �,�%M%��j �������0���-.�`<D�f�М)������vH�hI�Ϭ�(sge��٧kSw�3g�N������l4�������r0>�ܱ{�<8�I6���^9�zmo��!���8f�vf���)�.�z�o�z�������%J/0k�^�^����N��X�������vP�lN���'��3�?y��㙍9l���c4��!��jP<��|���`1��%>��C�ʊ�R(ɞ���VR;7/��W_��4"l$7��Õ��F�Rq0��ECo���ڢiV�8j�>_Ϝ��>��X&�K_c�i3���lq	)�V�t ӊ�r�g4t0�h|_��Ʃݐ�:M���{c��h��x���$X���Am;��'�
� �k�伞�Xb`�/�� '�΀�xqQ8uNѡL&C����6�Ys�p���rJ�piu��X <�:5k4o'�^]oon��:�~1/g7]k��k�}	����zd�f��ѴA�t��Վ�l&��İ��ϖwc�w�ƍ��������e�V׹ˍ���*��?u��n�<�XI��������! HI�r��$ƦY��[��Op��n��HIBJaU#)h��?�J���y�V���}��q�����wk�t�YM��`�����j3_L Ya9�_}��9�����Z\/�W��m���c}ݬ֔Tc���Ɠ_��u�՜})��OPs�I5�o]�l�ڎŨy;�|h���ɤ�������?��k?k�(
�i�FB��G��ys��|�dB��%M�?���x1����Q������ے� ��� $����A�P4Q�X�&-FC+�A�i+�1 chR(�)��z���]@�tr(J�
��e	A��(�8�(�$�NyHE)(%��Ӂo��!*�c�"��d� �3P��	 ���ܴv�A�OE�PV`!A�`4 Aq����h��ۜ>�a+�K;=56��E��~�	�SF.Q�k��|�Ch��'� �,^�'�!��cПn�T������kϯ����R��;���(��RL_�O��n�{Z"�W$�q�:�4�W�^�F������А��/���w��
�����8��
"�� �I�8]��c��A!�5�Hu ���7љq�,2=��|g*��<~��z0EjR�?��?T!)���_�����)H�lv�9�2�J`�cAO1��i�ɳ`,��I��(���b0z�8� Y')&��	� ��o�$�DIA��T4�_}~\��`��U� ��U�|��=�QuKO�&*���
�)�e�.�'Vn�R`���e�$�i�L,I�H�̈MAh$�KZ���O��1bG��� +\�0�#P� )F���dA�1h�m�]�P�Ax�E� )fdh�˅��Vy�� $��)#<&xr ��J*���F���%�`�-Q��ū�	1�X�o%G�,��b��(:�8�O��(��[U���&k 䒓� vULO�8�	%8�H+��.��&�F�\I��ĸ�!GI�D��,�&eIƓr�X1<�� j�	D���0�Ȅ�(1zY��mc삑�E!��(+1Lt�c�ƣ��P��%3Rh�/BW+���9 ���Pʫ��D�R��D	�(��H2�����%j+�� 4)���
�vda�`U�'��r�H-�u���7��Xk���f��i��NL���L@�@i�lRI� ��;�v�Ȫ1-�0��v�^�(X�gj�h)����4�i�)�b�Zf��h�u 1�$�x[���dr�@
����-&��q	 ��*E>u�� 5�ٖ2�$!��1��$� 0J�$�I-K��^j�O��C��� F���!7�Đ0�� �W���"	�2r8�8V�
�x[ r�F�mY�z�W���W��e|����i��SF�>8}���_������.�r��ع���h8/w���vV�O.fS����޷S�T]�1��ힴc������������������������ߝ��=����Yߵ�[׼2���G3󋎪��0�w@u�K�ܴ@ ����C��b8}�%�J�B	[���G	/�ش��Obd��P���iB.%� B� ^]���V���S�Ҩ�{�+��'NOˮ��-�
�r���_u�c�ٮ(��K�r�e�.G)�˘{���m#D�^;�u��:띃����ï>l��u���������*��j8YLv�7��e}��o�t�Ȋ�T�H�:�?P�â�o}/H��V�ϼ�F$�P�+�$��%�H�+L�m)����]%2a��q%���z�|ʒ�F�����ɇ������h��<����g���=�r�cwSF ge�����V|n���r֣		��w���V��D��w�Q5�n�Jc��u�ɇ��}U.�_��������ne��A�a�h�"�Ƽ^n�2ƦvO<��-1�9I�3/�u0��Ր<��*kb�[? `8�\YX Sb��Jl�D��&aG�-%40��N�٢K1���n)�����4������Q��~�kס����͞q�Y��#�r�����]����>�)|3�;�����������V������VH\}���/�����l�j^5ۣ�fx�\Nfns���a�m��˫\`Z�
EP$/���ϑ��z��'�!��F���?��^�[H������m�W�ܰ�#<�����/k��6�Ӷ�f�n�][��7\<ղ�ʂ�'G�����w�l�,�M<ϊ(s�e��z1�?޶��}]�Di`�U�\�m/�.�����b�{�d<��������ٴv0m�f˛��p�<�m^�jͪ���:e�r>�Y���	���  �2FR�%qqZ�h�Bh��=��m�܋�c	��.�� 2	O�k��+��@�.XI��W���`�dз=a�o1���������Ç�'�g�o��j.�v]��	�Ci`ex��>�4���W�	ڤmynt�=^�^���x�����ͫ��lx=�m;bϞ�Ű���v�f��U�ba/�CA����	�>�\}G��?�FKY�U�����-B�\
��� I�4�rT���$�L.��$1��FI�T2�C:,���i�&d�5WS7zp��lV�'�X��d3h�����ݓ�ݓ���a��m�ͷ�5s�Zf'���;eV����n��t:�?�|�L�w׷�������|8j������1[\������՝��ld�����O���%nd��K�%0C����@���������ȟ�PuM���,���SH��o��Iq�0$�S�8I߁�鰟~׊�^���q��Q;��@ۺzttzt|r�����v�����+�<4k��XX�m��]��f�դ6���������b��f�a8�S��h�V����Ͳ���8/�p�9�� P{�<�7q<�4�,d�8�?(ɉ�!�I��$v��H��Ad|
2�i\Ҭ�=�vb�B�q�S��(�8��oO;����V�����?q�DݲәN���ڇ���R�{�j�n]��5{��9�c357�Yܙ���np6�b�^]�N[� ��KUkL����Z�v�JL}\].n�������{;�j��A8���E� �y��M-�b�g��T�#5|
2��%2�O`#Rn��0q�\!A�,����|E@n�B`���+��ԴsMJ)>�ZB)�*BK� ��;5�x�3ò�kT	�Oj-+�|�ml���
����2�o�4��/���-jk��9��z��m�/�c��������R�Ӥ%+�� �i����Jۊ��*�Cz��3?�4���$S�9�d}�P�<��� #�AYt�BZ/��\Y!��*׌��r5o{�y;#�(#P\4�\>��-d��M���+�(�/�w~�]^Ln����Y�Ө�z��:	�pjYO�c�}N���o�j)��'߲���*3l˱#���3��t�r�QΚ��;���������u��G���کCB���T���(^b2���3��m�>n�s�l�~`@C��S	����ɍO�ѣ���<̶�Ԡ$��PU�J�h!f4Ӽ�H��( (W\~8T\�ήw#���F��hlE��y��I�].�w�鵽���r�O�է�����csh;�K�!H"�c,�2��Tapi����涤��D�nS7�6���_���F[^:>޷[��ς8�9�f;�ɕ�0R�&�t�n�7ҞOƁ�� 3r(NL 9��=\�cOA\��u�H+���r $���{S����F�$Q`�J!�n�J� Vvx���I�\�=�XA�b����@��0Q8,� �JI �dHY��8�`J���э�i���d*T��WD�\��Dq�N&F0@ ����$�I��d�/�v%"+��8l��C7d�	�$zI}��I�K�*��4�'!D1_.sj��,n�4� ��f��-��:ӊ$�����N�>��� #���<%�/^�7'���ߛU�JԐ�\�;~�e"��xP��=,��l	�$'s/�b�%F�?$v�3��ȍ$�������� � 0'3�A���1��~6����8(ľo�����#� ��TZ�OWe��֖YR�����/�0��0�5s+�"���BF�\5M%1i��C�d HV $� �&r`�J�&���(7�H�KmIYJ`�L� � ��,�"H���+W����U	E���e�^.%�"����8J� ��O��N��R������!B ѣp/�4�e²0��|�!��B#���> ���&0�BS�0i�����H@	I2L�&�n�@/Dm\�	�ǙD�SJ�\�JL v�9���*��Ll�fv��21J�*WY&Y��Q"C�L}(s ����W:��A,���X2��\�1�)@2����	G}b,!(aĞ����&-�Y�ɨ��S�V\E�JyH� ��L��:.O�,��VHTJF��@nCȔC��$b ���]� ]?$�d�'?.
W���L� Q>E�\Y��K$��B^�ڀ�贖5��Nĩ2I��B��d�$��@�&fFC.EC�,x� ](�2� �H�_���@q�oV#��
~w��j;��rm���0�;s�����j<)���옫������^���kvng�S}�V��9l�U�S�cDJ�d@�
�B��>�{%Y��ռ$���0�����p�dy�r)d�.@ܫ�s���c�a';Ue	�$����*���K���$�"$��(�s��-	[$zddb�aO��Q��:�9KʅǵM��D�(�)=r�F(�
R�,5���#��\j�ڣr��چ�|��������/�<>�g������t:��������jD�ZZ�yS��\h��]_�t�]�o-��=i���jt����^�뻳���l=�������xx��Oߞ��y�q�s>2�[n��M;#<��N��i��(X�
��.��H�E*7�@L�  �?ȍs�d�R̖@V�+�?�(���N@)0�.x,0�R��b3�6�@���͕+3�\{�������~9����#�f1u��x��Z�L����!������CG��t|Y�T/b��6v���7Z�����n�4[;�/�s��?O..O���W������zؘ ��sЬ��[ά�6�aմ� �D\=F�%v`�`���T��i����`Ĉ���@|�'<F��&��Q�=�Q`[)���V�<qu���n{������~�{������/������Fo��w:���v<���ʐɢ:Q�:����˥}�k<=����5y*r�5�W�4MZd�����i�}��W���?ݾ��폯/��Q�f��w�׆[{�I������t���{�(�6��+>a����v���x���
�I)�a˅�^Hx�D�R�X�D#7j�o*����0�`��t��dG֕�|5���p�;=|�������'��~��69lq1�t��8�E=Ks��eP�}�2�.r���lX���vR�'�ֽ��e��^��������7�G;;�Y�`g5����1+clFite�Q7�mƢ����e�aIp�!�]����N� �Z��>�W./!�"��N�廢P��-ı �� � +L鲼`ݣA�`og�nA[LZg��ww������㽃#cўQb�08�c;r蛁�r�jcA�)L�8˂�����k���a��0o�����q���/�˛�o�0{���w����ƾ�Ý�`25Y=�7&��s���F��9Ny�����Z#d���X6"����8P�+��q#�g��dƟvp$((U�2�� ���(	@Y�|�J�F�eF�mξ\r��m7�-]/�v�߻|����������Z��MX��|2���,�>���F*GȖΔ+l
�W�*SέU�a��x�<���/{���?�/~������47WW��Ƥ7��L}̘������tE� ����4�Q��1��� )���+1 2BdI�W� �	;�|�0�%�B �G��2���i���`�H@&�i�P���5B��\�M)?<�=ztds�;��VoPo{��88c���6��C՛�v�\������g�O��б���>��j�z�jy;9?{y�vd�k�^�F�N��O;ף��>K<��ϔdN�L���\Q�U�,e2R���R�ފ���C.0� &A�d�#9���0�$�E��N    IDAT�$<�HS".�XY��o�e:�0+�9��4V=w���tlx�s|������3��G���a9����wDW����Vmr�������Aڻf�j������_������ߞXOj��f�z�|��^�sW��N���]i*�-�����lQn�K��'���f#LeKq�,!~F��dxm�7��|�I��ŔX���'�䇛����4FO��h�+Z����*0[`�q}}u��O�?�?�8{oe�z:��_�ѵ�;x��e�������L(�w�{n����4�����j�,I��8Ir��k�E$���u��㫳�]�������7��}�[D�P�������=-D������{�����8=[�(�ר�3�d��\��ҋ���p�QJ-���X_�|�6�j�(Yu��Re ��	qb�~ �,I\a�%� �(�.��ϟ\V�6+����(Q \��4z����a���2X��lG�4s�G8֠o��#X&5�`��̀�5��"YOi���=���m61��G�_E6�{�~���L�س:��{6�Q��R�Mk���x���2�I`�uȟ<����?�e��G/c�	m��1P	qQ92n$� �GoS�~F@�����J�d�)z�D	Uѥj`4���{]����j8�3i�q��+��k���ttöm9۠����Ҡ���n��ݷ���o��Yu���I;=���:B/�Y�u�ŝ;!�7��+kQ�V��f�n�c�1�lf������î3������_��[��'�bnjsH��9������ ��銘�@��qT#D�G�����ېdjx�8s�:x�Q ﻈ�K��O�~��W�6u/x!ѓ)N�@�]MB���{�n:��.��_�|����||��߸u�!��I�pqNIu�x��)����+�����Y+������\h�n0u��,�2}W�˱�>dꍹ�7��rݯ)lmz��M��j8߻;����%PY�p:G�� ���1��Y6ac���P2���0&�ڳ,\l�@ J�0�L����x�C�OHY!�v\�aI�$1o��1bz �0B�A�wK�,H
��Ა�%£ @,��+bZ��B$PO)4�B��+��e!���C� Pʨ���^PJ�#��Ŋ�,er䢑��^�0�V�8�L�r��8š���i�h裦�)�P&���#$Ē#P��IE���^�\j����$� �@1\a������=F�33���@j��CL=:�`у>��$��K���(v�3�JmI�Cb�.EǂR�t�`��(ze��=c�I���v�����w­����ۿ�ۯ��������Nm���O��o��o���Y_'8���L�q����$z�#V<KШ��'����7���ՠ�G~�A�D�9dᅄ!
lo)8�� _ S�,���Q:5�q�'М�(F L(a��-���*�!��x#��#-�"$+���.օ��F��z0b�[$ ��Ѡ'?ED��)��XB	���X0���4H-�-�c�0d��B&)�a$�ቕ$Y��� Q
����(�dx�ԀT�}���c�=����`A�F2���������
O�8E��8^�"��!�"G��-&�����ƫ �U��OY�*��#�L��Ф� ��mՈ�H/9@X���l��L`4�ϩF���[Fj���\�vY���ph rY����Q���!��T�\1�m��Y�˂�4H�J�V�F`�&!�d�KF������C�\�Z~��x�ɡ�G>��H#�St�����)4V(7� S�X.	z<�C�_G2b�1Lh�Q/� ��!��!��X:�o'�u�$(E,D> ��:��L\bI�RGQ�����$���e�i9��S"XV����d��6���������W���%�G��l:ZN����.�7V����F�ұ���z�{��A�3жuc���dU�,N���Ŧ��hZe���͋�&�Ң�!���\�" !����}X��cl�� = �S�$o�#0H,0��L0FF����L���c��|��U�EҐ�.�$� �胞�� �X0��R.	Ȓ��G�
����9�J�F@/+�(H����B��|� /)@�&����oX��յUM3e~[��O?���珞�;s��c�ӻ�Fqa�ze[��gj_N�	���~P����Z�����F#��Ase������I
uo��[?�~�:�s�o$W�x�����u������;s@��۫��d=�hj�����|6��Ik�2��f��j��jE�~$��8?��B�$��J�$�h�o�Rz0�d!��KU��4Hb�a����+��Y?�<y��o�|��ܮ�����ѝS�ƫ����lW�kP4Em~ǵk� �v�5�r���������!���������{���d��o굻�������w�g�n�����t�~M?��W���� E��,/Ak'(�u�v���9<�u#xVs��?q&|�)K�K�X�R��$S,�S	�+F�D���C�߆��"��Q�j��ޑY5�ٞN����~���7?~rl��z�[��k�6��n�	�E{+�����vQF[�cd��ӏɦqZ��u'�ioV���j��=�ˬ�3�5v�8m=��.j?��������wǗ��F�vҸ���];�PM��z�5$>��d�C�YKy��r�-0�Ǳ`Y�8~��@q0�Lx�)M0$`��q���!�ϟMk��@��~#�o��x������A������狉.��>��ԸU����%ֈ���|zY�]�c��i!�뛮&���pY�������SsFw��P�~���ח?�9�v��kB�j����?�&w^I�)�g�b���8$���!�|��Ľ�������n,��]�`�|Z�!I=1MxIƮ���`�y ���o�t���}�S;��v�œ���<9)Å{��vX_���v�O���	��)+��\����?���Ϊ�HVB٭Sk-n���e��y&>�{6�����Y�÷���s�����,����,���p^s3�]������m�(�-Kc~`�<����&��?|%H�0��D,�B�Q��� S���݇���P,�*+~FP��|i�	�b�k�\1����s�h<8����ɳ��'���:
��]6zg����.B���7���h9�����llE��9_c�ߴ�N/���k+3��۫O6������?ܾ=������{�/������t};�]]�_�L�<���q���Y�F����dA�f�t5��Ů4�O��F�R}��s]X�tP�^^\ɍ&��#Y A2�T�RX�K���c���������~��s�ڞ+\=�ȱ��_���c8[�U,�+M��&,����)�v��XWx��[�f���q�XOV�l�N>����]�>��Y�n���|8��LWף��a��C(�͔d`�'����,x�ifb��8,ra�dY[��%i�b��)ȉ�CL$���`VP�� �����7��%n����L�͕�K�G�޿78==nu���������|KMH)��JQ�֚8k�AU�5��(,;V����,Ϊ��ϗ�߶������z��bq6��65gYߌtэ���vt�HZO���"c>n�(prZ�]��*sJ��P(^��?����+Yԩz \0�^0`.����E����I�]{���Tb*E5H�x� (3���/��������v��||whk���x�Sk�����4����z�����ǖ�����+E�2}�����ráG޾dO����io6ۼ|�LLt�֓��1�\�������K5-p�������fޞ5������}c����]��h�j���5�t��1{J�������*0����;T�O"�(c,-˽��z, �|"��d�LM�p&��4W���D0.j�����(�� /�E��ߍ�cc�[�2%߾}k��S¾(��2�k,?<zx��׆^�jK1�ZM�G����S�s��MSZ�{t�t~���v��.�7�����f8�M'vй�~4������j8�Z�����_}}���U�v�VoF߶�ܥj/�r�4����K�W�^�6l�۸���X��ɏ?�Ѷ�Y �XV��%�x9\�4�S��A�O�ȉ�Ĉ�%��VN�]�AWC�.�x���u�k��I�̆����p����{�vG�f������jʸ|Q�׾[J͖]��-���o�X�o�����/n���������K��,:�-��Ek�����O���]'n����s(ӧ��1�����j0NF|��5��\��ZT|��k{�<F��|��i�0�������  �e��,�I���$OV�%9 �"JY���w��ﯯ>\��{�_�u�k۾�q�9�jMg��<>��v��L)���fYg�ڱ6e��W�r<���E�[.�n�a^õk���|���?��x���˛KG��������o�7;���z'��7��w����@��36�a�M�h3�}��f/_�԰5u�aiLF/ ��b~ ���F�d8 �}�F2�h$���^�(r�*$!�����JYBާ��K�Jq��Cx2��\�Xq�o����&��J!��dI�J.����E��
ɒ�IPVx��JR�,�¨8b#����C" �rT"b ʐI�Lۖ�A�)&�K*[�"PRN�O��(Y(�D�`Đ�gR�e*M߮O�튖K��=j��V���4'MW@vB����e'7y��7��֬|�:�gϞ1�7�����>~��_3�����. ed1���#@[�ƙ�]��D%2%�̠Mԛ�TUY�����A�i�����C1�8R0����ďڬ$�lV{ԍ,��ۑD6���+��芒�L���fN�p�  �����I�O�7�|�,}(!���l�I�{��I�!��
�Lɂ�3�Uɟ���� / �q��")��˒���\��D.5��	2���/�0� ��$$1<z�,K,	 �(��`�n�"��K�>*!PG�Z�D�A�Ƕ&�oY�L�-�X0e���'��Ԏ�G�E��A�0e�Ȥm �AHJ�4�e� D2�����BN�� �1�� aD,�(���_�J����",�h���j�۷�)���C)�����P\��mP �+N�$^�bA&��
 �,��#6Ɉ#��Ɩ$Q�(E�b�Qnc�QR�L�	�$dT����TL���8�2ĩ_���"ޖ��8x���	Q�>�.Rn�%S_��}�t�).b#0aOӘ�%��P���
ڪAN�DY�(b�J�0�.!�(��*TɊk?r�Kx��z[�t���
�,�ڛ��r�'J�X �V�Q�7`d!��D@�,��8ʳ/�:3�r�`��L��O{:Tøei�kǄI�E�[�m�8n� �����g/�?������aZ���x�p��Z�zg�xp�����ㇻ��f�ݲ�t9��n\/�L[��~��I�30���K[Y���[F���sB�=��O 3��x&�� ��2 �IS_[�x��թ���Kt���`Ą`'�B%�ۖ;�XP)�###3��P|����#N�G��T1�Ȥ	$5�-V����CJn���@)l"$E�z1�Ȅ0R��d!�/���(�͍�[O\r��'%k�=��/^X	}��бV������ܻa��,	�C�o������K��]�OE9����W�8e��F,;���U���Xt~P����{�0n� 弾����M?~8�ӛ�oo~z��ۛI��mxW������W�k���,��,
�����8G���%�*����eL[�1ȸA�-BV��� )H�Q
��z��M'f4y���5��_|�"B5���n��Ʈ����3�9���s���];��؊Q���;W�d`�ji�on�in�����:7uǠ馇�G��i����ټ����~���lҼ����En�W��Q�V��%9F+�k�p�+�qi�!��e	��IV�(�@���v �!�^� �p�[0����GBɱ��x[' ��SiV��r�?0�ܹ����_<��Q��g;�!��ԡ.��/)#S���3{x�	�'�w����Ȗ��_nVk��y�{�M�w�鹘����.��uF����&mʺܬ�����?���w�˩7���p����񴼧4��B̧�d�똌&FV��>aB �+Ʈ퉷!\|(S�`�JIe!�aQ)��y1<������������۾w:8�?����Ã��5^`�;�����I��A10�r�&����Uk'����Em
 ���^z�2 �3�g�J5=���<����;����~n�s���~��>[���������լ�~�z��2��������|V+��Bܛ��,��T
���?bI:�%iQ>Ë/�\4$ d��2q|�!��^Gr] x���S�.d�#l�9�=y|b������AϹie��7�t���)jPf�g��ݣ��s�J_�p�p�~`���T��ݝ'�����M���G���mj絋�5߾��?^�O>^��l�[��G�WW���;��Ƈsb�xkf�b�f��xՓ	�oW��a��L5�>OA�� 18�p>�����H��@1J��X$=)�a�Qt��v�����a�?������y��^�3�w��RkP��X��}g+���2m���{:�����S���I�6{��ң~��U��ť@�B�k�a���|�����ץa_�k�����q9S�h�w.���W��+ �	L��89�'F޴R�����xRuD�'�>�!HA�����~�w��+=@�j��3Pw��������~v���OO3��:C����2@U�}t�΁����ֹЛ�E�W�K���A�.���7C�c����Vߥ�{��s/�L}����޿}�_���>�����hټ�7>�,.��&NX���3�@�,�~xa7


>nG��#.�:��PJ��a���"�X�� ���2��P�E�(�c�bY�$@@�]7(W�ڎ�,�[ɰnv;����{�����w	԰���lf�4\{���I��z$�n�zYkbe��e=�%xz���ehiG�B�Ѵ�P�|��x���W/zq�4;14;��_��݌�j��3���B-'B�9.�` )�-g5A
`Y�dX.���$�i`rĩ��4�0��F�"�#_i�%��_�3�C`Zr�
�=������zuy�?���Wg�̹y�Y��o��X��6=������O�뚭�lq�nE���];M����S'>K�v�u�<��)w+7:{��=�\@�l9@�_�ᠯ��n_o�^]�����t����i�=փ�uZݣ��A���I�ɣ}�<�ֻ;:��в}�l�,G<SL�Jq�1
�.���$��1L���+#����j�U
����e�hM՛=!���o��A�c�׬�QS��0(��H�X������،&ek@V�~m�r�����=��o	9J��
�M8Zg�l��_�AcCy/��2�Y���H����{��ݷ^���[,��|���9�woޖW��ݳ�x���O����ٳ/�k��lm���f�L9.�_�^��F1�0�-���g?�	y���C	0\��B��$	���	<K�A�����9W�D#Nš��8�����Û�7oߛ?���M�뛅�m��3[/�������G��T��~�5}6�Z$kȣ�bv��;TVǚ��[w[�f��^{�$E��H��g�6篮~z�8�j������=[�ɠ��\[�=�yy����k����gP�3�`�8�S�֌_����ی��M�r��:n���'��p%W�P
5s����'���+3:���SJ�$A���Ml_�M�o_�?{������a�
N�'�^�9�r����_�;<���5ٵ��鱬,u-�w�>�n���R7������nU��2����+}������������ݫ����nm��h��lZs�%������QM�ܰ[u��E!|����I��Ԏ�i����^�~�3a&
�6Ɂ���v2� �{�	��y�'A�X@ � B	@��Y鸐���    IDAT/Iϊ��w>�4�TڪQI-Q�؊M��zo���
^I�&�Kb��"3e� (���"R�(Y)]�F@��F#Lq�`���*����D/7�#H$M��]/�reQ{삑��>4�t��d��)P��� 6@ɿ�%3^)��+,@�,r2��S�,��(��+��d�Y?�*4 v���K�4T�D����7�K�+��P.��������L���ۊ]�6U}K K�5u�K��A��҇4x7h:�/�
*�E��tȖ�x�9 =iϟ?��	W:��5�����������4����i��;�L[I6#���6\���@�x�Yy��"Qx=����$��%�$��G�L�*Ȼ�����C>��,N;L7��*Zq<�2�j�݈LÛܴH�D��{5'_^��[�^�(1��,�]	^���j��!��^��J�F�ZeR����
��,㩖��+?K����j�p�E9����_&`��LG���|�Y��;�z�U-�[W XGvi��G�F +��m�$��UY�&F �]��C�	 2�4��!�A�F J$�EC&!b��W.@L�X�����¥,� E����)N�'��%�)�L,!ފM.&M����Fd��+��d�d�(�b����@�B��r�r���p$�+2� 7:��p�Fl
�zb��d��9:DU���#M�Md	�;�6�hY���MLOE�QL^ $>��#�(�>�rqm�����rY�
��B F�G�\�Ů�[B/7����@�2ak�`�"<!���ˍ��$2�bdl����%�@=�X�bQMd
� ���\H��WJ��-�L!��.�X����qd��F0�` ��JLU@���0 �BlE��Y(�%&9��e��b`ޚ�j;JY��vK�j|1����|w��l�Çsߔ��k�I�7~)�j��7.Y�^^z{��Ç�����8��˖;�x�貸�AYV|�%�I0*��3�� ��`�	r㓴F�Y�\##E�#G�X.d�I���H2H���m��$yG-r	�HT���V[���E#�W$0����g\y���xqW�+�ґN9���ڲ���?�j��9+(,1J)��Ēx#?��H70=IF�� ���{Q��$�{�k`V���ϯ��������/�?��/���>V�Fsx�YM�S�Р�L[I�0�#���GnD4�UF��h6N��[�i��Ì$.�y8+K����&�"����W����6m���A�l��Mی�_v����<}:����~z5�m���&b����c?��Kg�����d52��qj!�/�<�-�b�'=<g�T$��DI�X@���\>r ��McV����=�&�Zu?���t��m_~�����_����;u޽��nF7��h�4�r�e V\I�������,ק���bҀ�T�����Rr�K���s&�*#�`1�s�<|�jv~�:Գ~��6G��N��=���~�vs^��N�<?�M/W3?��>یk�<\��۫Q�<+S�������J�O(�ud\
)�ce��E۪^"D�����#*��>h�z.��x�H� �����0j�/jc���ڠ4�f�urt���ӟ��g�k܋�[���nh܊��o�2/C��F;(�Z�W���F�^�l��R���e5�
i��a.W��Pc>{���v��O��{3�ȩB�����=�޻��Q�O�迻�wv�w����~8�Y�S_�C@�Ól���e�b��D�c,��Cr��9���9`�gx�\b��H.���74�`����v(#��B��Ar��ۻ��/x���kD���n����a���~����.�[n&�˥��^�uJ�a�:�4��|(;�J�`�Ǖ���Ga;��H8�o�����Rw�u����t�������������G�ӻ����櫟?ֹ����x��h|m��3��L�os}�( �9�����Ӓ+۫�G� 
{��O�AQ90�� �A`:|�)"��W&���2�l�T�|�Q�K�O��O��O�n���c3��/�{���W��j�o��L�#��*[H�TS��u�Ux��-���=�ξs���G*����eF�U��˰y��lG�-V�f��;�[�;�V?�~S�{����ɫ�/o�>ܜ'�n�>u�^�;UѾ�l�p�o���{5��8���.��Ē��pN\)���0�ax�Z���$�U�!���84�W	`,f,=_���}��;p�s��쇵ửŮ�������_����{�D-���mzw���ŎO0/PN�>,��Oo<˃ �ė�I5��(�����
�����n��]N>N�h�����e۴=~�ݯ�??��������^]���z�$�����������;�C;��<�\�p_�l/Z��*\��< �� ����vqH��+Ir�Ʒ!�����r՗R�ޏ!��St�Z�*?���$�T�/8��.p�7����ѽ{�<���g&RC��]ygre��ʪ�Ҷ�r�o�]�v�3x[��C���G�E�T���ڸ�(�egc&~��ݽku���#��4���/�ϟ?:>=���|���7��.o:�h�N�{<)�6]�y7ܧ֥�`����P5�O�;�.�v�<� bB86�w�A|�7�B�\=����z;<"�EC�؃i�Үb/aݝ�&�s��t\~g��;h7����_�?���0���rv;s�)X������Q*S�6�y2���,��2c���u�$�{d����~��]�y��MWDڍ�{Xo���6'��Go��w���y���Wg����f�tqF�Yw̲w���}�.�x�%m5]�Lk&�\�8Joߊa��'Kc��jq�HB𒐈a8?�`\�F86|��_�F�:�4.������'���p;���zssus�����|��;o/˟���k��?<~�����ӝ��v��G82���f�g��Ă�b����x	�%�mo^�z��1�6Z�[�f��kʚ
�qo���T�F3�Em��������k3�o�z7�v.'���j��Y�������m��i��~�ص�&K�$-cltˇV�ܰ�r���i���'c�E�q0D˟Bܸ����xL.^R�� /_�ֶ�u��p��'O ��ʓ�}[k����P�1_�U�������;cc�����h���/��!v���\��ޙ�,���c�s�|	�t2��$~�Ȳ���h��S?�>#&���NW����TOC��Yn:���������Շ�e��a5ޭw�H�M�~�vk��mU��/�-jj��OUZ�RT�b+��,�tN�lș�*��f��:?��<����W�4f�l�ƽ�Ǔ�T��� aLd/2��&W�<r�C<I�A��>����V��^�ݼ={�������||�X�=�G��f��<<���/~v����%)�V�Գ�ۏ�����d[�v��G%��X�/��*��-'[I��&�����9�g���S�Ӯ�ԿԺ_ԟ>?y�֥yO��_�;��������坛�������v{�V��^&���|�����]T���3Ŵ�!��/O��R\A7N���v�?(�� ��M�$�9�M�D�vnҁ��_��M��uUfefeU��)�bѵ�/�B��|\�:�se�#i4�dw���lf��~d�π$�@  $��v�JUWL���p��ooϋZ�x�Ԃ�ӟ���$N �H٥�~,3���CZ�_���r��huMr��c7��]�<~�'���u��}�Q�|���n^v!�V����s�C��m̮{���h������?���Ϟ�_��;t����<y>>�{�B�\���5��6W���~T���Cʦ�䎯���SH����7�j�5Z��z�2�����������h =�PBr	MܩHB�><�>9�#X�A)z|A0�0�'!�(0����h����5*)B��#2$�.|R��ߡL�(,J1".8�U,|`�0G$�I. ��$">���}�È�
<M ��$�P��0� ��G��	��wM��J�I��$�ߓ�(&$�0(U*����雒Jc.������ �:��V� C u�r-���P��� ���~ǒ��Hq�Ť��HG`���[�t��wGl��\�
�u[4%n|I�k|G#K�Zʓ'O2y(!&Z����"	���*��P�˿���*��U��%J�
�z���d�Ux)I����0���1U�=������{���idR����/qV�IxR�UY�C�.��Y-j+T�m*��'�;%
eZ�T���%Q���j	�pB9[��@)չ�	�91�'���El�,����׶��yS7r8\j3�ӗ�o��ד9���������N�z�kea~4����b{�p�#<+=OJ����P�<����Q߯׻�{���������Lc�4�Vsj�(��y��A9JN�J|��ur�ȗ���D�^� �(Q2 ���I�����9Q�̗b(����SVR�#�6.��L�	�� �����|kXp���x>�p0"�L ��	��UrL8G6ᐈ`.2$n`���7�O��D	 ��DIPh���%'���GQ,:d�f�`W('4J��'?l��[#�!�)���3M:R%
�E���$���H����$I�%-�#��ANܩ>}��(	�	b|��� 0/(��d�,��l���O>1*��'i��'�� ��L�M� 0	�и�=Y��&A�DH��Dx�8��3�<3�O&���$����/40�pC	��U��Dü@"Ó�`B �(F���mB�DiaCF�stD�
u�������яO~��O��y���W{��'fz17��e�K��������qj��vF��S?����BO,�:�֯(���)��,Sӌ�<B&��d0�� �(�=2ĸ���a��8�B������	�F�S΂8H��Le�'�Bq@@ۢ�=!�n�����I440*�N�^����F��\����r�AapH����0(9C&8�0�&;0�9�RIK������n*�������ͺ�X����k��O|�׿���O�z�\�>p���OgG���}�E���&\5��K2�[{8U7��f�I;�#�=�&Vۓd�f�TD�jb��R��dk֏�P�cw��\��Q���J(��;.�.�[^^[�o;'���v/h-q�$��6Y��Ҁ4�N��/���V�}����Ҩ2��)|�T����>1�X���В�a��p�<Z\2�YXtV֪����O>z��'۷n\�N��^L�_�4Sb���yu��&�
�#b�ߘ>�����U�i�Z<�+);v=)�M��F�':3#�d��m_SR^�3�V��H�ph�l��?{q�^�w�mk��|��FZ�*�>Q��ᦆ2��)>5P.��LEc|�\�=X�AX� ��v=�mC'� ��e-�f$��d�)�A��k���i(�Ν�}v��{w�V]�t��s:���@%\5��*�*[&�J���<j��W,u֋�.�F��h��k����8�V?�	��[�tl���N���ٝ����lo}v�j�ڕ���G;���vwB��V����ɩ+��a���D�:�`�5��SRG-0Q&�9&&��<v�݆Ae��T�D����6L��e6L����-j���S��|Vf�2[��\]�����޿��fRzv|�U���hR_��!�T��;u������gQA-KNh�lRQ����V	���_5���rօ�s��B��Y�K��Z��ǹ:�փ97����2��/��� k��<
�MɃ�!��	��P���Pr���pe���.L��c._�!'�T��:�bu�1'ZMM_Y�w����!�n�dֺ�l����ܼnO�3v/��e�^d�� �j��x�/���m�L ��]{�1J�IW5�)��1��v@��{�^+�yݷߙ�έ\8��ݽyec�z�������xp1X��kAE˷'cފ)E܊am\�]�9�a��$y�y ��k4�^D��gd"�QJA(�)2<S��g��R����*���t^hлX��ٛ�sm�w�}o��])1�p�uM��-N��Jʿ�\JwDT�j�ԙ�*�7c�I��ۺ�_���a(g�V�8��p�[����u��]T���ro�6g�^����9�w.�D}qfD�ycB}����ʽ�Yj�M�D�e� s�Q@]�F�^':��4`��� �f����'���D��wJgc�U��/-�̆�-~�n^�t��͏?�sg��gK��{��kJ�W��_�qj���H�������Xل�.@-�f-6��s�:w�����{f�溓�w5�t1\��Y��/����68�Er8���Ў0�עt�4)St"���C�#dj& �J\i���������q����gh�0����Y�N��6*����
G�#�<�_[[����j;��g;�b�o.����G��V7��poo���MRu=$���3�'�Q����� q��s�ֺ��1+������GFn�����?ff�/�W;��
�Ҭ3�3���ž�D<�֩��b��svY�+E��ڻ�Gzu+�M�Anj�z�h
+�����CH�\�(|Ah��iD��4%ᇤ�:�ԧ�)�b���tZI1��bn���|��7_~�����÷_/�o��9��:�ww�ޣ�;�n�ߺ�pZ�b���"��u�cOf�#�c!�ju��� S�%v����נ��ha��O�cw~0ӧu�ȊƤֆlq#i�o��Y�<���K�[O�S�­@�N{�/��:=�����6�Zp�����U�^)�8���4�9���2}l�Ҽ��HT~KZ�#��%�[#��20b!�+���J�V;(r���L#q�#����d�������"C�G��\��:�|���G��n�ci�>.&���'r�6�9�yA��r��T݀R�:� ZUq/��c��"o��s?���_�~qr8��à̌�p�p��ڊC���5���gɻ����~�g�݃�?tN�&v�\���{��OhY-n���s�����NC��-P�>�N?�4�F4Cu�dte$�
��1>��8b���loo߻w����A 5�8HWC.��x;<�����g�~��o>�y����U��Y�{8�l޼���g}����m��t���?��t��϶**R�lUu{$�J�/���;�x-!���>6��0�*�E��}�r�8��=�^Zҽ����b�=�zuqs��噋�ݗ~�׻�~f*"�Ϟ;����NaZ[�����wk��rY���n;�d�U*3��?��s�I�����qE�j� r�I��3Q���ܸq��͛��
O!�At����K������7�}�_nJ��|�j�?�ܝY�}n�Z}����ln��
�p�Ğ�<����?����+�C��_x���s'�N��E?�{���!j�����`�U�{�^����;��;>׫�j@ox�(����+7n��M٦��iof��Ob{:���X�F&_�ߔ�]h�V��C��8�� Q�샕�O�gb�Q�7�3ŋ|X%�(�)Ĵ�Mق��ɀ�V)�)e"�o�C�#�4-!%_�����s*�f�C0!�$�Z.�Є�耈n8�U0�\e�e$U��!eA��SBQ��T��%�� OC�'�� ��zH՞x"
"��	'#��!g\R�-��i#�1I.���>XE��KD)ꛬ�Y��2G#����Y/0&>Y?�5F���&2e��B����*�Ǐ���S������DM�ʝ��!i#�E��h��S��P�,�
ƈ��"��S�t��_>y��YR��g�������mCZ��^DL���?��?;����_���/����w�T�)ʿEMݤ�ɔ냗u׬YJ��(o�	3>�*At�Ul��z���ﾣ�^c+�Co��AL2=��N6Lh��Q��J�O�EA ��2,
���q>!�7����̄�D�D'?��Klݥ]�{�����m��R�ё�{�o��~�w����m���:��(�V�{+î���E��z����_b���97h��?7��d��~F:?cw��կ�sh��:���h?    IDAT��=�m8,Y�3Չ�L��T��њ1_���$�bA�Ni d��.B�C���3$ e��hէ��L��2��k�%'(|����0��������$=7R7MGN�0a ���>c&�͊��m��?�\��
e8$dB	���$�H�Ѕ��$�q�䇲	R�ئܙ[#�ͦ�9��/dK�������$��!M>a�|7/0q1��ą2��*`�br�ã��&
ʄ&	0$ߧ��	��|���$bJ��c��Vr��)}>Eć�f*	8>	C�� y|��x�bE�%:�+J"�L,@����DOhhR�	g�r�����1�|QPr�p��?48Z�sJ���K�	?��@����	m<ʓzX�q�����$~wѦA�y���Y*.xs��/����������3���E0)_���]�7���N�Ҧ��t����p��C.Z3�s�$��&���ÔA���S�o�P ��-Y �*�@������%����\(a�������D�W���9�@��OA��s��[>��
nA�&�u"m&�ͥg̵��+|DD������ <���."X��B����	%?���$�D ���BtH�g��pN�8 ��`��īB�3���\^Zp�� ����'|v�޽������d����K�l�W�Z���u�f�T���]�LUQftQʜr�D.��Es�G6L��������tי��ڄn�}2�3�Xs�g��k݋������������̄#������:��,�6J!r�,h#*�������E��T~���UE~J@Y|.dM{U�9��	��!h�D�*��)queU��~U����W~��>��Õ�]��?w�꧓Ɂ��b�O[�3�R_�w�69����Z��Z�Y>�~�KMx�ѳ��tm�@=�c;2iFL1�Ku�z ?bk~��ײ�9�;�3S�̮u��׮����ԑ�S�ƴ@����۷H�h�E�eJ�]��G��E��Lh�1�i� ��������� �������iD�J�~�Aw�8w�����h�������?�x{ssÚ���o��Ϗ9��,��_��S*|�5H�Q�mom���)�Q5��kET}�����ː�먦nŒ�$�5�hk������䰻�v^�K��K�k33?��VN�?�C��i�?Gk�>���Ruڵ�E��G��T?}r>�����J� H�T~>�DO�k�ӕ���R��(���Zv�5ـ=oK�;/�;�B�¸u��/~����a��zJ�M�f��M�֬]A�FG!d�^eH,�����ҟj�ꡤ��^
�4�&k��E�E�յ&�)��1}y|�U3����������G�g����`�<z-?�س�@�H�t
�=/!�8��	�i�],}�&�U	�����) -{��|���<#�p���D+Ǥ�o|�,��=���������h^��}��֧�{��pk��*�+Ѷ�t��~$T�����u��&�����vAF���� �J��MunSRemJg5�{�̳���v��?�hUY��ݘY���b�b̨��fН�������౬�U�_��]��&�TT6��
�r��߲�DC&��$k�o	�jx�듞E�:�>�}��P""㌹��nv�u.�̿��Ƨ�ؾw��N�`6������ⱳ'eU�Q�j1Fq��+�2��\��Z.�HXύ���ɳ�	_�r:v�R���s��*4X�X��[�,�v�NL�<`�wh�CN��̳����
`RX�ָW?�Q��RE���´�3��RS4�EX�7�	��(�15&� G2A0������F_C��Uc^�G8YooD��ebq���>�~��yy��~����*��鑩jm����V��Uy�NϭIT�A*����S� z4����5e��|:%0�i�����E���X�7�؆��K�޻|ic�sy4{�s`k��eѺc�����EQ����M�Ƞ��$?J�������|��D��K(?��LPi�U�U95KE��"e˵��Z��
����l�K�3�k+}�ՑÅ��ƍK��߼�����+23�'e��xo�������l���k��.��`k���!t]`�J̰g3����Z���G���9��k|Rw�/���V�7�W{������^��[tIv�P������$��B����fv$4�B�dzW��0Mgo�!`�C�����a"�j�����	��ׯ��j��G���L�ӑɤ݃�?���o�����z��z�w�<Z��vn^_������o]ݼa�?��v�G��lN�ղ|��"�c��T�K��:���P�t��ji�hH��%�aVjl��zTV��)*t@���f�,ԯͮ�Z�ܽ���)�Epi�Qᤧ�v���d��דC�Rzpն-mFgYV�Pq��e�y����R�ۍ6hO+ �5
N�D�Q� ��^x4t�H6��9���x4�J�wJ�iB�&X�pV������4V��/z���?xx�5��f#O'��==&Hm2��9O�-�p#_魪��i��}"��F�|�$j�m�Maci0r:S��~�0ڬ��LKh���#���������ZL��[�.�W�d0����O���F�2):��3�g8�o��@��*`K�zst���*($z�ah)xZ��V����I���Ci���������V���DD�Ch�w_�zx����埾�������d�Ǝ��{~p����l���{W��Ym��������g{�_�d�gP�m����P򂮕���g0N��X��M����E2� ��/%?Ol�q,��w���=`dg���v���Fw��tete�?k��w&���=?��v'?��r�;��B�cף���J5��DI�_Ů�Z�jɾ�xK�ǩ ��4SJl4�萊�+����z��P���ӶK�l� ��ǰ�Sk~z�o�y����_����z�֧~\zGcc�����~����k6��n=~��ϯ~����?������d��Fior�]�n����G��y��ٞ׾g�������oa̓~ӱp������Eo/�ml,�Fv�u�~*2?s�g��ÉY/��jr�4*��M�T�hus>����3"2�t��@�B�ƹ��  �OA	M&�l�N(q0��p0��H|Ab�A�!*S��O$�&N\��|���5��a��`� �1i�K����M�L���0�!X�
i�<�B�) �&<}"�O�"a`"(yà�N\9Ȧ��8��$.Qa|�y���T �" Gv�'_�`��1n�r��eE�n:lEA_܌B}Z������/���/���?Yd���c���F��쐹���(�_X�j���������?���d-j���Ҵh�T-޽{w{{�:#Q�~��W�e�qf1�$�{�$m�[��7o�A��%���PQ��	g٥�uT�c���_�
/�.&�@����8�ɒB"�XV4�����O�p��L�+Y����C�!4���E8�Zg�k9I("�Rx�/b��GC��!�$%���������� +�Sb?*U��w����bV�F��x��;Lr�|��?[�2���^w8�*����1��+��7�l7޺v�����������ե��.-^Y��z�W�W�����+v��.��ƶX7\�f�^q4M�k�\3qi�-#�e3
�s��NƅF� .Z�WQR������"j�,��� �!	�#�� 2p�zHp-�2���'QnJ#V>��T��']~���4
d88B��'& �CO� N��:��Ez�%i����A,����GiB�dAbΡ�|�>�r��u��Ѹ��^�� "�X��4o<�h�P����D!>���C"��F;����#ʔ��5<dB%�.��!EILu$bA2I�Ȓ.�I�O�p��°6�<�%��Ї���@� <��ɟF	@	Q`xJ7I�knڲ �	����"&;�&�6[����N�'J��N<|��|���
M�a.z�#�����t�>�p�|`BW�����P�'��ȸp $
�$���O��jv�0��w��^X�8�ΐ�+��������_O�/��sO~k`�A�]��ˣ*�_�ʽf!M�xua����H�������t0W3ݵ����������V�$��}r))�T`	&�X�N�kN���ħ�BpF�I1%�-']d�`䕮�9�||D�D�2@e������D�?������h�~���c ��tRɯI�r�˩�|d�/���$����p�$�|A ���$��X��}��yW3�"$wB�O��Xɭk�V�nZ���ݑ�������gW/�LQ�~y��z�xl0cT	�
�'�vUJ�S�\!̀������JB��$�r���'S��X�57�������Q����C� ��Wlm\2�b4'�/,���7(�^c~ut6㞨�m���bj	�N.���.{Q.ѰWj�h��*�n�������}�I >&|Q80_Z	LK!@(��068�����Օe#(o4>|x����[w7�f'3�;�?==�ݳ:Y��4�Ge���em�N�T���0�m�1P�PU�h�UL5�UF��aD �A��t��~he�]/����G�_����ޥم;��q�����^[s�'ޖ4䮅mV��Z�H=}@��lu�i	�V�O��ZQT��J�@Fۂ }�ĂI�$$�KZ��a��X�S���n���6r�����׮��W��p}cu��Ӄ����n<j���"�u�4�E*�3���^[�l�+]�($�$��h���R;/K����$����j/���LE�ـ���}?���;��ז��/��/�;�s�sHq�*�c�e��2�IOB!i���ceG�'< =?�k�CY� �^�)H�!�&y�	��Ð����u*%�?2&�ClK�UO�gG�����=|���ͫk�������+�$4Ạ�x.�/�W��2T�t�uW�Q&!4-s�&VT�ߜ��3>P6ʫ2��7Kde��j�)����܂�Җ>�]i��e�z��3Q��p���E�I�t!i�Ҹ|J�SD
&����*��CB�����c
|h�	l&SQ�BNoj�9�d��������>�Ž�7.y�����½zw�XvM2��u���Vd)�����F}��U��[@qP�t?Y4B����1��g���̄՚��İ^PuFv������Z�RT�\���c���z6�=������Z����_j�e�UG�Q<dB��N} z�D�%.$�sT�V#:��O>>��R�bN�v�h���VGC�-���֍�_�����|4Z2UfGN]�v����i.����ʱ5	�Z3�:���Ѡ�,�(�2��/�v��<V,�bU�� �uP��6R�ڒ��[@��������������Q��\��r0W�N��[%�<J��Q|���1�F�mGi��6؆��3
T�VɩN���w����8A��(i���M�ke�q*�1���s���^X\XYZ��}�7�l]����AK2��wt0�V4�$��r�&])Q�&k�eA���q�*'̀��C��`�ŏ�Dϭ<0R��A�tI,~]�|�`��p2W�г����Zg�7��>�|q|��cWs����ѺS���(��3]P���'8��G! �Oxq�\`���p)D z�,|�gbUkҎۣ�F JOg����5�6�+�^%��6�63[�����u�+�
��=�;�(<;�V�I����ƴ���L�.�0�K�O�Xtk�57噀������C	՘�W��J�؆��\��v��aϕ������������W�~�u`�ҙ��Ťp[$jHR��z���OUHy�P�D���U��GQQSg��PA0S=��G���è���ES&+M�������6D�C�|��<�������w���'V}�O��C>�]ܻw�����ܺ9��l({�wp��zL����У��F��/fV	��*
�`�_����Zc��ѵ��ʨ%&���(ICg=(�.[�є�kjǅ�z�����K��������gs��ts˞��.Ҟ��}0\�4�6�P ���{S�9iF��&M������"z��ab ���U_!2)l�)V3�΁ܿߤ�EMx��� 1�JV��U�����S�V{��<�����\Z�����M�y�K�6iݻ���b5�j}��cV���y��ȷ�Yg<�jc�F̬��c�`ٷ����j��cZ&�ꩭ�μ'<�F���Z��Y�;���ﳓ����g�]Vsp:3�aX���*9�
�`ˋ|�:~�jۇ���M���W>ڠ�8y��a��H�h�eS��Ģpά��m��t��1q���]�&�8��Ó���v^�|qrืEH�
��������}kK1N�'��q���^0���i�L7Oo�Zh��Rv[l�ݴT����<jr��i���X]T��Y�¥�z�W/_�e:�3PUA/f�f����YY3!��f��q���Ŝ���ヽ�4�p��i�&K�5���V�F�N��qJ`�MA hX�zغ��O�9b��£�DG {�d�ζ��C�\�����q���f����1��~���8,��������R�΍��>|psk�7_g��������&�ݓ�WM�"��st�l��o��,�&@��H�aSDn�Ս:/�%5�����N =u�|�;��\���&[���V������R�˶��AyM�\ .;{�uk*O���M6U���U���@~)��m4ɧ
H~>����������z����O�&9��%�(��č�D�\�S@x&�I�]�%��rI�83P�$$�i��>#'�D�%<��sI"��q�g�;�#6҂�Z�j�	�!d�	��H�7����$ �>9�F* ��H�Q��'�x8���������L'�XqR�� &�I(JJ��'�)�Fe�A��˳{��,R~��_�����*��_t+�O�>%F��,a~��WO�<�ēϐF�>I�>�^L�F�XҒ ��7tsLg�A`�4��u�C!F��OD�fYʎ��Yg�>n`����Zbt��~h�b�q�g�bDV9`�O��O:N�����xi������!+$��C\4�l��ˁ�=*{���O�ZԔGJQD�~�,E��3b��9AR�8ZF��P�0E b�@�  ��>�B�(͐�ɖ(ί����߅E�	�<V�]�:پ��\vE�Ρ��-��H��'^���Xq�֭W����޾��U��#�sk����\پ��[�o\�}�����s����w�߸u�ʵ���6���o޼ric~e�Ϲ�Ł��L�l�a�?ڄ�p��G�?�ˈ<��1�/�PΧ,s �橅����e£0u�84��&��s"�O��8�)�(��)/���� Q���Cą���pKP�0 уL��S24�ˇ�J*"r&V�����&��Cna� ���Q8�P�&	�4��`�A,0�:�̈�׈�pU=�c� �ϩ�I�O08�$�?B
�=�D#!8H�����䑏<���%.�p�2I͌f �0z� d�!-�A����I���,>�	��|J(> ^��r ɉ��L��q ��OBQ�b�	��)D<Y���Yt̕ �������!�P�t�����^_��+�P&-A�4ΧX��+Jѹ������L�䚏>�� =�7ILbj��%�6*%�Ezs�Ź���|ux�
�W߿����$���k����Dg��Ln�3�t~V���L���t�lf0Z]��&�4oB9o��1έ�ޚ#��	�kP`��bs�����mlI�1�|�f� |Ч,0�]�%�!Q���!� q�#�� sAq"p���Y(aDDOT>>¸G�v�O,���qh3���+Q�.U��d�
$\D�'u ���g�A� 0D�24�+k\�'"i���$����bA&�`��H@3�:y�Z�$dN�����<zt�ʥ�����Ov_��Gߥ{��k���߱ħ����9�����	����O�m��7F�c�G~�4��G�;k~q�yrۚ�����9q.յ%����������݋��pdNn8�ߜ]�͏��v�p:Y��5Sr���    IDAT�����f����ҧ �}�a8@\(q�Xx�X�B�b����P4��I��TL*��^\�'�s��zc�_~��o���K}O��|��ӓ�}[���̈́3`V˫��8u��ɪ+�,l�O��YWT�qq�՚G;,X�F�B+��s Ň�������Z�����L��2P�5E6[� -@ҿ�փ=N�|b_����я�c/j)^��m�E�VQ�k��ZԔqڠ%'����/���/*-EQ�T� �£�(���>���N�%��6����Dl~_�6F���������~xg��r���b�07s�YI��I��JX4��l��,Vӂ����m �B��4����[ƺ��m�����TS�/�/-�͠5V4�8g�1X���M�̓7�c'��+�˞$;x�'Q�C꽘�����;���ST�1�H�'ub��铣7Q8E�p�O]�,D�a0�p��$� 1���L1�.�z��0�z�fi>����rnIq����Kv_37ݦ-dJN"�і�k��D��i���� [p�E�MͶ�V�j8�o�LZ�G�%+�گ���9e���%�=?27�f`����������������x���avn`�YCR���p���J��R]�@PT
/9�>I�K<���$՘�D�+A>C��	=1$N71;�{pyua�rg�)�?���׏�֖z��>�;��Љ�x�!��YN/�I�N�k�����`ke2�B.�3��u�ZWgj�Z���ji�Y;�jb��m˖:S��U�Zo��и?�!U�I=��R���ՙW���9_U[5�=��+��%'噜&�D�i�4��h5p�����r�0I�� Hd���R���a8I�9�k��D���%�Ov������������[��KԪ���ɑ��S���إ�⠶5���ue@��R��M2B�k��҅bQ7�L�m����A���>����z���iw����L�2�n>Ыv�WO{k��������=Y3��Vm���[Zʽ�yk7 tB	�Mu�S�)$d�Wf=Q\wa�C�y����Z�L\:T�SdQ��0<���$>VFa�{y�8�����{�m~����WW�T]J8��9=:P}(��'f��F�u=��͘�~9�mx�J��堀�-'�K������I�2(�k����������m)
�����Wnd���3?ۿ��ѻ�ڛ���3���+&o���P´���N��/~tB-�ɯ�[��&JK(��ZUf�����%<��i�'F��aM�Yh������l}e~c}~qpV[�;�k����p�����ե2Ň�hy69�&MҢ�j R�C��j�J�l,k[+CU���P�k��(�����Q7�Q!u�U���Fe�mx�W���'Lř�H����Xe]�';g�#3S3sG��-�~��5k����4E8J�I	���sf�%kZ/[q4��11q�8S�������1g�ՠ[�o����{�����?����8<m�ऽ��y���G޲�_#�����ⱝ�o
]��Z3lc�v��V�D.ɨ.���� t�h�����T`Q�b���F&zF��o��%�bc�^�,��=��^�]��ۜ[���.zg�>��у�^��3��2���b.�u�u����8���)Mk��"�$�<M��RV+e��N) �s����y�ݻg>֜r��"��R+�ֆ�>5�̘�)U�R��lu�ƕ[7/-�{����`ߎ�Z1���ua$"#�MGU���RU�����mU�Z f�k!Y���ٿY���ྺh`��:KC��ڮɲ���Rg8�]�[�4�8z�p��'�^�g�V�]=��)���R��I�jI�-)��bxn*��=��E�Nȕ1$93K�ѼOb�0 j/~���P�m4��S���msXu��(D.�}�E>y��ŷ����O/N�\�R�`o����>���G��._�[f���;?=u�1�Џ-��.�������e��9W&��Y%�eG)k���VӾ�j}����N{"��\��7��_��ٟ9�xcV�;�ݥ[�W�W6�z���}�7����D��N�&��U��X���Sf���+����+SU*��� I�@�� ��9U���=H����&[/��L��$*M��⦬����޳�������Yo��$_X>��zm����}�`�Ҧ��������Ǔ��J%ZUP��qk�xOtt�g{A�]烬*pU���nh�T��҃6)-#M���ބ���������dg�~����E��~iy}��0s��uY �����<C{Po�:$�[��O6S��4y���6�pQ/$�M{����h�zC
�	� ��(`SK@7�L,Q8x><��D�&2A"b��J��b����%�0Q���lI%���Hx��I��%b�e�*��	%4>�ÿ
��h�x��8yz�$��F�ƛ�@l�m?jp��*T��ydB�V6ÕXBQ�Y����N�@@0�����_ � Q�h����^tAI� �h��=!�>����ji�̓'O4 ��O}��\*���丙�F�?�z�h�"<x 1J.	�6����?�љQ|,������4HV�,����_|a����3��Oq-�t�Y�B������5H��ǹ	����\Y�$�)�������D��s���̓$��keL�Ų�*IfK��A��#�t#-��$�.LL�S:&�p���NA|^�qh���JNAT�Ras0h�!�pn�Dq���Nn��+�?Gf�֖G�{?ܼ��m�3ޖ�����������~x����M�������߹�}gs�������ˋ��,�_�.,u�^��^��m�w���K������psv��`�Rg�roes����խ���˛�6o\�v��3��6���oI�^�Mkhk�:F����H�C]��V�!e|�%yO~�UG]S�QU�� @�bq�p�'8jG	��P�� $��`�F�2邓\��Jt�����Hb������OL�dX�|&h�!��`�U1I@&
�0$��@:ĝ*!�D�D4O~�>�/" &H��'ʰ��Є�U	e'������(�i�a�P��O�||q"�C H1a�Ex���#�%i���* e/�s��� ��GN0��y*�����}��1	��
&�D��gD�
� j�K .�ͧ�$�S\Q���r�OA�ON(G�`ѱ��>����D*���XH~D
^\4����*bvҧ ���-��V���Q�4���^YN֒��l�1��|@��K����� <�@�������������D��O�Ź�d^�K!*��Jo8w�p~��o�~�⇝����V�9I�1jEʼ��)�MM�MW}u�P�pus}���ʼ���8�?��hp�6��P�E���O9���s`�ӧ�5���E�$(����
@�p��傃PIN( ���p0S��(h|r��_�|k��аeMLj�E�-u���T�5� ������3Z�ڛ��@Z#��(��y�q�LcEu�!KDp�(#�%���D#4H��Ih��:�(��@U����*�sW6������<��?��6��祗3z}}e��Y�S��Hڇ��X#��ߜJ�j��&���rFA��U�p-[i�&\J95cY2;�W��L�n��s��,�a����.�\*���h�kŁ�Ε������h��EYSn��{��vfUGNS4�B��(���`I�2u>ED�s�I� ����g���_�[-5�V�F��Q��G���󥝙��Ý�W�O��o:7�aM�$5�Gg�*��[lಕX�%�*��V3h&���EW?��S�f.�d�G��ֈ���eQ��(�������R�=�53��Y1K��$ݙ��i�����}�\��3���-���j��~\WB��f)?C$���6���U�Á�Ҩ+Z����S|Q5���V+�FY��WU��t���:^mo�����7>��მ��L��OwO'�\��MB����RSKa�	D?�3�j�OW��n��Vc�y&/e�R� �e6�V�&V��y٪�M	V�6��ִ��Ɏi�C�lV�d�a�������K��5]ļ� �w��3���LMK�y��z�B��T<��.2����_��A(C�hHуT`�߸ZS�
�L�����ܼ;T{�67>�凷o_�7K�����(��2��Ўv]^e�i:��~3�rX�.ojN��Ш�J7��.�FvTX�J
�(��V�c�-7X2��)s�r1a���jN��{C�5/fm��u�O��t<6�V�i]E��1�W	�^��7m9*%8�F9��������D��?��`Z%i��RAS��Y��1��pv�n//���4����͍O�ރ��V�����Y6Ʀ-:������h���T�j�m�jZ��Jeڵ�ç����1_^SZ�ު������e�frk9��~{)?��崗���n�k����u�7ϯ,����O������Y	]������:�?P��&�cxE3Qx�j�a�p�<��`���}�^0�UO�n���OAS�� �:�!tqq��4Z��(yi���{nC}t��:���w��I3^'���Z�l��%<C`��~�h�,L �%�U+`y�9�u�3'���u.���QQ�)���.�:��Y�i򲮪t[��e��#{�,9{nvƒ�`v}�|f����=0z�@�g;�O"PQu'mh�,E�>I+T��cm�{�/���E̞@���d&%H����g8�������$̰.�pW���?���G7/�-Q�wy�J{k�y����0!f5�:�["�o��R�兲��S�2F�tm����0co%���G�K�G6]5��j�ˌ��Z1���k��n�p�����nMi��R��-���v�&;GF's~	؎$Q��5�Q� T�y'O�!����4�X\B��G/"��,4��H"A	e�.`y�Ӌg}V��뽵ќ�pϖ�޺��o޿�u�~���nq�	�(���#���$���&�5�����f��6��`�#r�y����N�6��ޣ����p�m�5�]�c-7W�[L,�_8c\6�t���	7�b����K�ێv]��x�uZp�z���6ZZ�\�qٗj4F-�(,��h�S��a��a�o�lQl���y�X�E޺uˬ����: ٭��NĠaw������__�x�m���Z�]��_}����ݫ���h��a��,}Wa�[}b-�X�<6��z]:dޛ�(}�e���*��"�Y�R�Lc�$���JP�L$�Կ�&h����d�8pm��ܨ��-�t�;F,/���-6~\Lz�A�A/��z�VI�^�]R��@���j���(��ِ�0�k��Ū��-T�(���{�,[H6��6=(�7�������qa+����Jg`�u����p�ܢ���.U�m��J^�-�i��`�*L#F��WEvGp-�]�Y��B�� �����hk�n��*khV���v�f�Q�FTw�x��zy0�;X��J��%.�w���V��E�N�-����l���Ƚ9�L�V7�z6X�M'Ĥ�"l]�	^M���d5_N�+)H�V�_�n*�A��Q"S)�J���Π��b�嫯�㿞}���h�� ڷ���=���/�oo�r�e�����'��.p7�O�S�-��RCܪ���eS?85��߸V��ȡ�rQ��v��������m�D��I*�s�	K�{���<�f������K���=۫��Y�9ǔ�O'����mbPS���;T]�0��+@�V�2���C�M���eYh�Y*$_��V,�bO������D��?�����O����܌'Zg�V�)��_|t��{������?>�y��`�_w �Uu�R1v�9;�=�T�?ֱփ�~o���'r�Ĵ�����w�0�&���`~�kl�H��.���8�Y��'G&˲��-.'g��c{�<�^�H+���;Td��X�K����Ic�K�µ�n���2�
��
+���Qb2-/� 4��"C���c��xr蹄�2�*bD*x4`N�O�(;�F�óX���ĉIР
������� �X�� �O��	�ɧd�#%�$$T����#mxb�X�E�J����)�qC���!�D	>qq�`T[����G&9lEkD�Cr�"B&	�t-o��U3s��	i���i���Ȼ��WeQSw����,�a�3��!Xv'����t���������gN#�(z�o���	ɬMJ�j��Ez�S�EB����/!-�f":4�㓵U�`R1ײ�U;-����c����+�,���`+�,>"��J#]���0��I2mM/r����D>�@,
ݑ�j%b��b�̌[�ty��5m=;K��~�����-Qb�)EH,��I(E��8���m��CIl�� �`.��!ݮ'и`�ղ&9�f��L�٘Zݵc�=���5�N-��giu}uqy^w�����	OC2bbh{˪�y���1���c:RZrК��!5��b�ƒ
�t=��U#9��.��?{�T/Ԉ�{u�p��X�������w�·zIo����i�e�/� �Ih��(JԂ�
EI]jb��o�R��iq�	�E��	<'��R@�iE�%����0��Ѡ�9D!��p�K�ز	�J�IŇL�0����	��ą�08�P�޲�	ϗ�i6C n0a��S�EQ.|�H
s�}��Չ�a�B�Rt� �� D����#�D��G���Tl� ��������@�F��!`EHp"���Q�+;��*(�UŁ�*Y��|���gp>�CN�&'������A�	��B��->b)�$Iz����2�IH�X|��aL�������,0��%b>��ӂN.�Gqш�a$DC ����P( ��� 4�B�&0�� nRA,�7)5�+CH�1�b�Ty4�1I���'����}�I�Z���~?ֺ��j��
�����U��tNz������&�ұkW_��6"��U�oAÈ��tg����{��/T�ι�ŭ �#W�#�#��DoQ9�M�If.y�L�V�Oq�˧T8H�=u1��
�QrI+l�� Q>N�H����[�+bL�#U�&���淖���h �(�L��ORvbBZA2`�.�q�����&�}�> &���'$2b���>A�>Q��H8�#㋎ F���4�4���ta���'��ݿ��ؙ��G�kT�s���s ����gfDi�.&C�W�(E;���3(͸�{h�k���.��W�}�B9o�̺g�&�u�~K���lL˰��w��cw������'ߘf^]�\����s��\����`�D��+?��o��bN]Q?"���S~��S�o�0�%4A� ���� �'���g���tRU�mwO�pmeDYJ�����7�,o�h�������COk���\��S����	˺]?�U��{�z��Lk��񕝳&���ә���%x����bU�xrw�VC���;YQ��@�%���	vW/�~ֲh�eG;�����|�r�zo�wv�������L�.q���/f���gk�����j@~�ĩ��ӂ���b����)80�.:�>T"ڋ�����r��!K��G����������"�P��hSJY�VdV��ǳss*d�S�K�X˜�oم7���NO�5�Zo�2�j�	��B�p`zf��Z׍,m�G�ھ�^�%���v���^x
�x���`����Y�Q��w�{��+�'�4-�yu6p>hn�EM�AF
�Π�z�E����d�!(1�ZW���L��p!T%y�!Ê/J-�7WSNqͻ��D/)҇7�^����ݭ+�����ώ�T/��Ҷ:2�D1Rs+�'�AZ�)2���U�U���W.�g�W�M�D�e�l����jkT�M�-��B}aͻ�]4�\�MZ�������8�3e�tz��_,,o|~��_��B-:�7�~�;�u�F9�\jW��:"�u��M�QQ�7�'���˵�ZEQo J=4Ӷ#-AM9U���U����Kk�K�چ�˫||��������k.�s� ~���g��P1�\�٣/V����9u���j��Z�sQ��ۿ��e�}���Q��QR�T98|�.T�������LO��4-P�    IDAT�N.�.�ǃӵ���n��tq��ҽ�w`����;K;�"�;�q\�/��� ��U&	H<�s%�ր8�8���Dgm�'�Xh22�jީ�`���~�y.��2��VF�}���/�,�z���+���׺�Z
6��ǎNԪ�k�u`��Z��&��9��P�-YZ��*��9���%1��J[��b�8\�e�]���+�֪=2BJď�2A���gG���p�R׊���kk�f�w��=_��kX���ݥW��ã�FņH�2���9�Qu�ď�rT�c
�Nђ��]�o.p��O��I!�Q�|���	 �O��f�� �G��w9�++��wn^�v��;� վ��C�W�_R+�[�=ŭ*6k�����#	-kG�c��~Ŷ*����<0��y�2g΃Z'��G�yUw@V�LFT�����\�[$�5�Y����dx�w��O�˃�|�_����cS����f+L�%�%��@t�F]���[h�B�"惩(b#�h>��<C&�U�*���i:�
ON;���6�#�?�uw�^z��{~���w���ܵ��uY�3h�*�2�0�#��3:hZ�>����V0&��v��j� Uo^�������n~��`+L���Wͮk�1S�N+3D��������A���p�`�ް����G�[g�3�	���{NѮ9�;vij]�o�T'�s|����rr**��$
�I&��V@���@�����Y`�y�_s��WdB��zwi�d���g�}��/~z����XR�,���x�k�/_%���#/O� 5��5%K��fE�C���Sd7$�2�_*em��!�TL�@#n�6��(�t�Lt(�	�v���>�s�S�����:���<3r鏺��������[���M�t釽�g��������;���]��������_)�D�iJ�v�����%I�ݻwMl�{~�D�ҏ>e<5*�&m4I�fG�a�B3�L�F�	:C�|*M����/���/�~����;�_�/y�ҦK*u4�NR֑n6��y��O>T��Ďw����-5S�Z9kA풒vp�.���֍K�%�]���;�UG6�v$]tO&��g�G����g�W?�ף3�rw�׵�}<��Ov�t�8}n��s '���j�c��V�oXD�Z]�v���8d}��!��%�S��%0� J���Ԡ�dv�2��XJjX�%j�V��.9?��}��/z��d�Sg;3Å��?���G[�k�㽗�t|�S+�͌X�:jO��3����6��˶K�k��n��^7_)+��ڍS�1�GQ� O�' w�����p�n_�;�?���GǗu�++3��y����m��o�����o^������,�/g�o�����9P]+%
����v����� �n��e&�P� ��w
P,�!q ���h���"3&\��[�4��k�J��|D�����������U>[Y=�p�����͚���*C��T5� �v�'^���'��ޮ�����Soe�؞-�be�Fϕz�&�|R5���l�G7���]\�s�c>qcA~����վ'{�#
tnq��'�[��������W{�Nz�[���~������fFKn��~EͳI�Z��X���A�-��ݢÜa��)�XQ R�5�Kۥ���z�9�LK�a���`5�,�Z{�o���$��P>���F�b.T,HS��|���>U2m�$h*UX�r�%@�0��X��e�
�H8�p2�3	%
�i�	���)�O0�8H��+AI1��"&��}G ��2Ó�RMgj�_�?jH�#������*B�Ĝ����R�,dX�LB�������_�R�폟��C����
 Kx��� h�z(�NBZIW�_}���%J�,Oʂ���-JH�ht^l������Kf�����	b7�$�ƘD�?��&��	f�S۩cC�ֲ'����ֽ{��V��$͏odc�v{{۩M���ۿ��o~��[��7'>�tj )�$s!���N��cE�YT�[%��� {��)�(:�#�0�k�ՏTR	�INf���L(J�`�'���i��\��Ѣ�rFu��|�ͅ������������G�=x��ܿ���r�
�T��W�ͧ��������?N^>3az������n]{�������/������m/����|���Ý�/�5�����W/�'/]n,b�i��ӑ�%S�j{�s���:Z-�.�o��s��($�3zK�(��m���8���C��
��$(�B �Z(4�D��LRW
Ȣp�\ʅυ!Q�e1��h� p x �1d�J(<�)ϐ���s�~&n"����bA��dA�$�dM��CrE��"6$�OAI%���8��>q��	�L"	�&��"�,�K���Q�x&��&�''�>ᣍ�֔g>�_����D�ǦR��C2�c�P0O�<aa���)cC/z4#b$�&��	Rt4�H��"���a$?%����0@d����"A�qQ&8�E�!|������{x��!�edҊH|��h�Xa��$�x��B�X����'J��Ixl�@b2��'E~b%_��V�� ��?`dD�"��pB	C�B�oR��E�4������`sq:�&'���������������C���͹�E0ze�1�,��zΊ�z���x���tu���kÙO�L�ǌ����yg�+egd��n3�M^�ɏ*ⓖK�	?E8A��W)��J�����_�{�߷�z����>�c�X�$Q�o����J�%9D'I�7�73������=՟�]Z�٬^���Ꮷz"�psE�v�C���P���(q F�$�i.B/Yh S	��	�LD~��Q���3��V�9����$Ό:��
������{��O�]��;~�ϙ��\���gM��ԟ�;��������{�.YRp��w�m�S�Mӊ'�eXr`J]��x���E�(���P���cI5�NS�Mv�x�p�mw�"m�k���b���1[�a�z=��̮��20��0�?<�5���c�>5���ŕ}�
Y�: �4�AT� *��Ps)�)2eħyQ�nB�fC1X��]X\z�у_}�����_��/�=�^���L�g������k�ˊf����?�%�Tc?f<s�g�<;�c
�t���n��a��x����б)�Z�u˓�=�� ��̆1ӏ�k���P?�-�,�:fj-��Iq|27k�����'�>�,͑C1o˛�j;m����]�K��E�^)�I��$�F$�\;��muu��M�'��>w��L��$�� @b2�6[��:[��)oOK����4���O�9ǽ+��f
�D�N.���!Ӳ����09	l�[5���g�o'W�2-�";��]��vY����v��7n�������n�W�!_a��L���eq70����գ��X�W�C��ͣĐ�4^$�Y��<�E�&KBY�qk��pQ�w�Z}�bsTxLې{A��<����t�yq�bTnT�o�������(�ܞ�+�c�Y
��0�8��Mv��	�֛ �(<������K7���7����E/2.� �]����������э���a?f��h��!2B�"QL�qv�P���{�$�`���5���P5cfݦ�#����`b�P�O����F�ޝG7���qQ�Mk�4�>��q�Gg��!5��@���Egќ]�=��2��2ZdX�6���<~h��H崌d�/qȓ��D�X��Q�dr'H�����}�����=4�tč�=����{?����=j�#e�!��Y�����F�1$�lC��Z�jZ9m�\��KvT%�L8�7�2����l�}-���Fa����v�ٶ9�WX�����8���$����\�VwUݩ���_y^K�L��fk'վ��O�=Y!� ���|�[���ʒLK~�>�� �R����?ĬR�J0���d��&����4*�f��?��ǟ=�\��~�cݲi�z5�ᦌ`1�d��0	wh�M6nd2�n��ψCJ\�x퓴�o;AZ�a{;�P����g�ۙ��_ń��Ӎ����a�`JXR]5��|��t$��,����FT���*�r �^\039�	ڪ*˟,R�� ��L@`�@�l?����D)�8 SΈ�x-AU�{t!6�������'��=v�f6�G�iF�n��G���,����ș�'��K�a�W����m�d��B���H��gzg.VLC�zl��5�pL�<����'�]V�X3���qLf0p+�]�u}����LZ����3�lJĒ����b*{r;Y�ٰqF�@<�nS`����ggxb�L��Ƭ��-�i�M䲋9S<� �����=���|�w����~�	�\$'K��
�y���%C,�f��\>�3<A\q��D�L�r�'��1�;S���<S�q�+����N��6��!��x�^r��!� �.���N����Ț�t��OMȭ�*���N���X���z����wH
�zzC�i� A0��(@�4�9��?�XL�'ɬYJ��އ�!d�� ,��ݻg%Nї�(I �I+�Et�r��%~���������I�ZU�vۏ><�����?{p.d���&�u��q�lm#=V_1ZB^cY�#�OJ{gv>���r�R���B�m5LTء0�sb��G5b
�q@��Nt�)�q���l]Xg��L؞��>�bpqI��{W;��U����鸖�q�����9��"$[��XMqab]/k���\�y���g`\����k��Ukђ�gB,��T
Ni���_S��.���'����}��=�>)���Q��FP5XԀi�c�qRSBZL�6 <��v�hljE�*H�Fxe��]W��N���Ѭ2�^�	�RXD ���H(W�k�6Nj���k[�Оzm��8���.k�A&���|A,b��\ A�ʰk�l�?gz�@�d���p�S4u����>|He���d��b9�v�f�r^����o~��_z�͊����������v���]��~�3��S��Cn`��5m�iݱ����ťգ����ޱ�~ӈp�9��v������D���X�\3⠅	����'&-�#���Ri2�5��Jc"jQ�m�v[���(�5��AeYL7ˣ�|g��)2I7�R�+�
��ń�7��x0�?q��K�$��J,�D��j8��ѣ�Ńy6H���x|9�yiޞ�{󜶼�T����ݽ�����>x���������������&nM^YX�Ŝ��\b�b�����X�3�kG��9��M��2�C�K�i�~���1T���ZÚ(��)\���{��u,�&n��ZL(�6h׺a�|}5��'�*�=�I\@K���N�K�b�� ��b0 ���s$�Ov��s�*9�?���dT��ୟ������\���OQ���t!£��+�G��dZy)��������E�\Z_.i�Q&�!H0�A.���@�3iH<bEm�I�@؀%�ϐ,l�y�f.	�_���� ^�|}?�E%$��'��r����'d�TY.���,`���{^TA(V����e��A8����Fdj��Z���M�94�*�]v9���,�>x��=���8���۷e��B�����/ɨ��M��!!H��(�����ÇI`	egĔ���_��uO?�3��0Dy����~fN��/���A�}V��>�93Qi�!�H��AZ~��;��������]� ��A��%`��=OR�l��)�\nݺ%o����0�a��g9l����h_,�0=IR�?x �����4Ӌ�{�`�5Q�k��+Q%b� �͈���fݪ����[�j��=:ڋ�򇻱���֛�f��bہ6m1�!9�b�+u�h��.9��t
|$�B�y-�b���!�п�@tE��hؚX[XI��3Ǡ�W�׊F��j6 ���#�������_ľ���, Ͻ�E��FrZ�ˬ&\��p�W,�Ҙ�٩�}d��"��hҢ�̏� u	��O�'�M�<
E	����b��WF�Ar ��ɯ��K��		U[�5E�����p�d �(i�&�J�Ĝ��dC"Q'*���gR���Z� ��[����6���d����lV@~�����T�p	#D����d*y%?7?%R ?Iئh�(�&G�\��H�U"�Gڄ��+I<��͟	�8}b<�y*�$�D!x��+�%��2m�CrF >�㛐	 � �2��X�$�L�)>R	�3<� ɺ�ޑ��Q�$հ\t.�9��p�Η����G�,��$C^<�}�L0� C�|A���dy3�������3H���
NƓ��"�6c� ZQ~��+�CH�'��ى�S1�J0ut�f�
��z�-'�����̃��z��u�h0�m�z���g{i�ĕ�8�k�`Jn5�(Y8�+ͪꉋ���
]ڼTo��ӯ{���$6���h��/�*��-�b����K�EʋZ_~9�bT�W`:ժ��S~��!�d�-�~�_ �~�	�d��Y_�KU���I6��H���"r?�����#��Ta�&C�g���m��xw�ZbQ�j����ҷpu��@O�(�\�SoAm9�G��ϾP�|+a�g[�;���"��jC���\�a08�,RD�H���256�a슁�Y�j��7[�F*�u��{=8X�����1�*�_��P� Ǌv�FNX�"�Ą^�Ȣ���\�mY.m�=�C���a�8d�v��b�Πښ��\�*�f,��Z��+�+�Z�dR�tqӞPHc\�D��Y����������)5o�~н7��~��Uj&��Z��"-n�js��Z'^K.i$<�Z������|�គ�?�d즂6--1��v(U�=?�$�:�V�����?���[5�������"�D�����l݅�x�1�cf=��8��X?CuZ��x�͝z��s���q;x��7g�<��Fhtv�\c��zl�ۢ�!�4Z���y�9Ԗ��c��=a�OK3o�հ�^nmg�Vj�����?*���zy:a�_nUV{v�g�hi�4��]�N���]�U�\�A݄?�s��?9�.��\���ۢ�GH\R��5`� �]w���ik�5�!䙝��wo��x��e<��QX֭t�J�E�8n��Q�FPi��F�Ӑ�Բr���!w��dR4��z�b����sg1���]��LG`��+l\U�^��Y����۰���ـ�9��X���R����Q{U:��|z�{z���l�]2��d��ɖ6�����1Hr�#��VB�hB��<L�ǟ�a�h�p�S�(�;���~rb}����x��arX;�5���V��E&�N�����{����+Ov�o�@��4�R=:�{�Zԣc�^J��'h��rC�#8�(ƦE�)tѪ����֤����������mz�>B�M"���NU 
E��*]��b3�T�Z����¥����'�ǭ?�~�t�rp�Cr�^/�.�/�v�o�&�5:f�4���C������ϔJǓ� H �jWB�p��JAt�b�ս���b88<������9���h��Xg� ml����C�/.�E-�e�Pf		}�PlGJj��Z����H3�%��>���,&���b��L��*���2�-P8���O�� 3���y�ؼ&i���|��KՖnը|���j5������f��g�⚵�I�Ъ1��:��
$��p�� ��	��f�F� ���gY8�)U�P��6��ܯ���@s��n�z�8>����;۬)i��E%oʆ�p�As�T�k��;"�X%�cc��Ҹ�F�}�	��82dX���ijt�$�ZY/vd͖��{�*q)��"�-�	B*D�����]�к�e
�Z���i������{��×X�$��M�r�:f	8�A�=��VGX��Y2C�����,��&�$����0�HD����!�0 ��Ĳk3��/5��{i���=�˟|��a�N��G�F$9��-�#=�E1/T������rD�e��t���&!������"�EJ��H    IDAT X��jD�v�i���RS�JiB%νNEq���C}%��C���`�|u���x���v���CP�z����Ջ5��]G�MCM�8n*�b�S��+���:�dr�'�RbDI�J�6�C`���ou%h���T���B�"	[�;����F�:>����?}��{�[����(pf��6g���Ƙ�}1! .@ѿɮ�L�	�ы�p��1�b��)]Oh�cAD�K��)�b��0�4���j����U��a�fnǇ�:�}G�ff��Z�3�sǩJ�-�J;����i��^���ի���f�eiL�l�X3����Fbޟ���g�/�1��_A��DEEd���9����3ڧ�t�4��/�9��@�����xB7���_�^ʦQu	~�ީ�}����7ol;�4�\�����)'0�j`dL�b�����ӑ����[��J&_Ѻ�2q�lQR��#(�d~e{RZ��FI�N��G�ƶJC���[1�99mm�8�o��픚{�v�}�����q��x�X�k��S��'�F���w8W�r�2�4�+V��v���������K�\e�o�=?�h�bs�O_JSLM��Ʌ��u�N�q'���ɓ���g���d��N��N$��^�^��{B1!��6�̀<^Yj�'��j��IY�=@���8T��[`�.����*�t�ɇZ����K����/�KU�r�:.6��;!�ݔQ#�������N����ʁ��_�b�z�pk����}��R�{g�<�۩�4��j�����z����n�ܹ=����A�߸�ꓮ�\��7�[��w�w�YZx�O��ѣG�6�՚F�/&s��8�����|�?�z��'�~��ht�����~��~��>�6:��W��WӾ=�\�����7,+΍�#�{,ڿm^C$v�e��p[޼ג��F!lH���0C�Up�4o�G[q�pZb��X�x��
$�(�6�j���������{�e�a�����f��OK������_���S�������A;�%%0b��s^�^�y�U\�m`ʁ�Q��bQ����X�E;,ڪ@U�	�emh���?��U̀����P�8Q������_�=I����Vcq�������['w������7Ͽ��2f��]2�^�����&���r��>o,˭u�ӄ��7�����)D̮�\�����R��޽��E����F��U+�`K���ku����g�O�g���s͓����4v��b�4
k���⛯��9���0�X�'����ܲ�q<��<Đ�����T�M
���U�9�X��:c�� �r~
���oPS�\��'Ob�!���Qfx~&@6_��ˁT_�2��|�+��<��6�B �Q	BRt �T��������7r\�ېlʕTe.h���	'y�Mj�����x�N��?RiE%���gx��61$�����͵;�Ev/`,�R�yKn$6����x���kP{3����'�%ȿ�˿�a��)�|�����}�򥼞>}�R�Y���Kg��=)�&A��?�#�������P�\;����
D|�T����h<�������F��:���տ�����/~�*$�E^q���>�E�r���8����2Ŧ'O���t�Q�r���iL}|��2��p����fE�h:��� U��(C����J��~9��a��l�/��0��� �Q<��^�s��B, M�ZN\�ل�p+�Z�u��.���k��*���ɝnB���v;�ktK71Lx��(&`�Q�`�Zu�?:��Z4V?3�X�Ƣ� v���)�]��8���V�)r�M�c>��U�I����y��)d�N���Z�[a9�m�l��D�f�����ϟ�:����^����Alښ�X�#6��Q����Q�,N&���g���on
�Xl�|TI"<��p�d��L3��%��K�<��V!�9����VH�xh�a~"�&��D?�ÿ	LH_�	Ll����~&�	� !�6�x ,-��$��O~H��<7���< s&L>d�`|�O?<b9��̯@�t��G��� �� �f�~f?L��Mxf�<��7	� n�u��%�J�9	9IH���%�E�p��t/0& �,�s�$K!/E�$~BR��P�	y�q���'%<�H�B��$2�@�I%\*d��9��D����r�����G,�ğ4 Kj'2	0N� �I�X,U?�\�
�E�p�	Lr�r#���I�U�/�6yI(<��嫌��M�CQ�{kD.B�R�J�|��4��=�W�V_�K��?f�y=��1����!��=p���u�2=3�w��ᚕ"�%X�Q.؟���\:�����0!���a�a�Hj�O.Y�~�h�����J�n�4�^�9?��-	�wp;Se�T�E 0��� ��K%�G�p�I��D��`8���Z�A|:*�4_/Mk�e���@�z����E���WG���h4�+T�MzQeU��Ř�İ�7+���NI�� �HM˗I[��4Ð�A��U�$g� @|�H"-� ��JBj�1++�ڨ�v�〵W4*��o�ɟ�Ӛ��W�A?�ڴ���a�&7��	����Z�����M� ������`4���x�vbB����r�O�YB�֕f=8�~*�a�~����r���D�Y��JM1Va<2�Z�l�J�����������/�g�-P���ܼ����/_^Lg��-n�\z;�6�rJ�@|Fm5�PQ�w3o���d�S*B�	��u�i���"O�`2?�Re��DUo�%�����������tP������
�޳IX;Z����őP�Q�zBW7z(e����u98�\�[���u]�����M����A��jfS%�����e�񳆇���\M�����=je{,4kz:�h8��U����]ZM������a1�ǋ��Imkћ8pk�e[ә�#,+�1ht�K\�"���d�(Yh�
.�_�j��LV�����V����@�{]g���V��Iw������>�y��-��+����bX�P�^ �Oƥ�6ج�.K�0qD�1 '�&��x<���@Î#�؛p�	�C�����JA�74	U����jw�ڰ�'r=5�
uN͢�B+���{��FX(�G���W.I�����v��y����;�ߍ0�W�ŀ���j��S:S�8!�^QhR�L[Ѕ�T<I�����Q��p��!,���I��p�M���)R��"L�uHƜ��nő%�'�=���.���	3ͮdc��.�M�x�T����'�)4d��|���c:2!L�Np��gtZB�/Q$�B����%���by���nA׶w�)nS	�x��c��8T(�b���.��1�ƺ��%�����I�w�r6iN����2+O�բ�qR��$n��Fl���df�(�Ï��O|��s�_�Mx���A�	 9����-S�ZX��o�YR���,7�?����w�Cu5�9�A�E�E	�h�qg(.%[\��#-�؆W���T(�� �>FP`��}dW�m��A�!\����5��b�XL����yxHd�0w4�4J�:Z�[���ݱIGj{����|=��wO��˺�����t��~;�Yݣ-��'��������T�n?o����u<�z܆���+�Q��I`�R�@fem8�5L�����B��޲��{�������k	�x�ޠ����:;JB�X�z7,��:2��C$��2��� BhD���X��R
�!B*�T�hRQ�!B��1�N�����K#�W��k�}��̝��6N� D�!N��È4s�!�F����?�̡��/�����d9�jg�x�4� 3��b:�˾�c�����	TM��ɐ��7�M��)UѢB� KV��(6~���=�|�������?���{5��ېFh���t�`�R�
�B� �7��j���S7��⹯����>��3T����w��:z<����5+jv����P[�8;�Fڎ���Ն�r"i��D̕�տ���\�v�׵���O~~u=�n�]�:�z����Hގ�o9�i��\r7rFAtP���e���@Q��ړ�����r=%�G+��"���VX{W��ݦ�1V�w��}p��G�m��8ף܌dSP����CN�h�俭 s*ڞ���R�g����|Hb�݇]��v����F��!�,D�f�-�m1��f2^5VW��,�=P�ǌ��T:1E��3�����Qi���.ڍw��Y̾/�E�Q�um�Ρ;��g蘅:^'�ԛ��j��9,�a!<�=��T�pN���s�,��f�'�!�� 0�x�j4�3�����of�+Ě��v���o}����ݎ$�Y߂N��G�t��ui�����Ǧ��n�C�!l>�����-�b�dN`%o�se�cPkt=)���<iv�Ls�Wcf'J��H]��$���T���q���)��.w֗12ۋ[��v���ҭǷ���z�d�f8-���-L�O�m=m����ov��׭�~���r���]�5�������8C���"�Q��}5-?9���%��՘UD�0 ��C�;P+?}���<�X�%��?���4ک9��f��R���tDG����b~c��E҉$���H�Z����zH�kTQ�F7-n��L�īlYיS��������G*"C���M���`K{1�H��>3!��m�tw}oq�,e:�����~o~?�_�ƽ֛�.�,���Bz���r�QRݎ��{�y���n��S���Ƙ���#
���9�G�bS���f[� ������6ǅS������%� f����?�䓏>�T�]�]�2*vI~Ĺ�E�1a.�R����j�J�M{&���Oq�#.���M��l��JH[��F�8�M�T����#��i~3q�c���ڨZ���ض6~�[���:]�ΰQ��~�#���?~�<��ۼ�W�?o]^�n�=�v&G{�
�uǍ��-��[l�N�ѯ���r�ab�N9���{!��0�Yac�$!O���j�Y�*fM�Gˑ7��|�������i�z��n>x|��|rpp����'/�~m��"	��QŜ!f�����-�	km�����6&��^ZZ��؞7�35�__!����|3�l2+<���C�V�����H�EԡQ����d}y�:�b���ꎅ�KQ_���i-��Z���z�7�Ί�s�Z2�O���^��0jm��6.!8�
���* �p~�-~�p<O	9	�^6�����z'�g�d�D�6aP`�MɅ�#�X�OHx@��'��Y%S?|S�@Q8��-�D���b�i���t���~x�,�Q��A��̑G�	��WȆۢ�ў�%�}����.�DB��d�����d������H�r_.�
�����WxF�6��� ��2�@
�x��!�{���~_�!iO��G�������3�ems�o��c��K���\���
�9���A�_�6���PE��0��?���yY�����EI�3�ɉ���#`$�*`͈���S�����`tU��ڪT$H�+��� �;�H6łhk����_}�����ۿ�`xV�F����Hi�T��F!%�Ef��2.�W����4O�"!HQY��2�%�W�|g/]ǝK
ZJ�V������6�`q���f�wn�v�;�;{,�XF��#�2�&�&���i�F5�� �X��W�mdZ�0��諕ř�P��� 
�8�T�s1AƩ��X�����#�ߝ�Y�M3^�X��W��5�a	�6���`w�֭��~�;�v0�Aed���Ò75�Z=���d����a .a `��$5`��w�B~�ڸ(TL��?���O�h�!	#�'C�BQ������� "_�Æ���l ����6�f^r89`J-�'3��$#P�N��2�L��ɴx�E>1�p�����<j��l�L囨ĊJA��%�p��(�� �gZq�m}���& '6.=��$�dZ��Ox �@_�EI�+\l&��"<���?�`Y��ȓ?e����-H���x�g8��O�1D%��xh��E1��>h��%1D�䙻���#	����D���LLr~�R�S���e�' Q9�#�G��(N��!� ����J!�(���'�̼��@�D*x60< e���
�ϡa���Q+pSX`B|3DT�2��ڰb�����,��4|ub-��%��I�8�	N6���jV]�����r�Ym��J��m;�&�W��*y>�M�\Y�Ԇ�gKr��-i�{a�ҫTt��6���p�4�:,���M�Q˟E��r!Om�Sa��.������SG{�_I���mx�&��"��MTd���<�Y�� �U��p��cc ��6���im�b��rJ�+�-G�%aІ�;61�mJo�R�j2�Ai��|Ҧ��t6���]�Q%����g��9���$Xlr�W��	�A"\1��`ࠧ�w� s���.]��V�N��we�����!]7��jS���O�	6���G�<v[sꝮ�lt5���9.����߷�a�<:��")��P����Vv��4l�Y�6�''�Ӆ�zf[�{K���Y��&
^[	BE�W-c-?]���><9��v�O�.n]�oW�8H=gkz͸�11g��U4�lX�c���«��Q����9�6��V�L�?��8�1/Wnܼ���}z�}���ճ�|iG�\[Z �R�����4͔�fIWU�b�)�j&G��<����j����r0NV��rh��^o�;G燦c,~P�wb}_��m���l5;���۔��0<k�шe��Ԗ��y��ڊ���>�X��n�9�>��[��a�6�o~~��^�o�/V���+m��j�ڦU�>���z����Um��a���9F%��
|�o�i�����x�����#���qD�N�gE��-��t˞�ry�������k6�AJѧ)���G��n����Z:sZ�3�RIZn�~���������,Ϯ������l9���;3�P��}Hu�OM�I�[�ʻW���j{�m�������I���n�O9Z���E�t1�P�;g���u�l����|�?/��O�����=��z��S��}�C���Ѱq2Y�gJ���]�)�C:�E��Dq���6,J�y�����&�Y��6�=8y��f�lˤ��#�F�}b#���CS� �- ��@�����ڱ]<�����e���7�-�ZјkK��C�kZ1t��0m����[�n��x��x�`wg�m����æ�%@\����I�ٽ���7�>�hچ��N�Թ�|�{3�t�R��Z���e��u�b�9�!א�.�n����<B�g�
.��8���¥Jf�p�O��SZ!�V�:6B?��a�6s���Z[|��G�����x� m�ɪe�)c��T���;�4�v��f�JL�֣�5�"�?b �Z�z`��B���;��j��6'P�y��w��=����Mֿ=IR/�g�Q2���m}ɔ9
��]�b��ګ����J��>���/�խ;7��z���jqUk��l9�b��(V�إҵG���X����ㄋ�=��Q��-�3R�d, �}%� G�dr�%ԑ�"��xz�y�W{po��Qc>�a��ssUWsSCq��B���hڱA����#�]�������=�\^��,���d��YQ�\qmȜ��`�30Nsww���ܺ�?�fm�W��K�4�c�]]j�ź;�S4ͮ6�Wf˝�#/V��x�����ף��+Vk���J��9c=lIV��A����͛2$��E���z�c�O.c�PAYG�AD�6c�+^ת׏o�������A
C�.�`�p�2~���8-Ea�
KнZ;�Cz3Xmc�F�'W�7㳫�E|5�������m�8�`릘_�c�#�}M�*�{���ݮ���L��h�Y�e!�m�O�:ӭ�m��Qu+�zdXj5�k�u��䳺ס~u�=QS]uY/�ż��R��	�dćd�B`or#�hri�oo    IDATU,^���	)m2�O��Q��dA����S��]��{��e�Ư�x��Ǐ�č�Z6�$��|ز��&�	4g+�A�yܠB7Y�:}���d0Z�L����cN�_,%�t:�c���c;��j̯y7��{t����Oŷ�f�қ|.���9!�iX���́�99G�R��z�~��Je���{���:lx8'���}U^^���nc�0VĖHX&��'�i g0��L�CQY&!��\��פ����H��`�^$1��J����7�����<ъc��V��ӟ}v�m�B�d��r�!kQ�xV�e������k'�BR�Q�0���{��s7���p0����.�Oc�K���?��cVq]��$�B��I����~����<vh|�vIH!bԋ��'���0�6v�Ẍ́�lٱ��)����zQo���Y��b�tu9z��W"��ۏ����ƭЈ6T\l���\"���=>>n�s�*�ym ���A�݌�ob>V���[lN?�i�O=��_|��w�� ^.��=������]��)���c�u�2��R��1T���֓x4~=�X���tOn�.��!�o���pK\��~竝�Bajm�C�h�h��6����흭�Qߕ{�e1�OuL� u����h���3��I䶶�ުҩ�xt�c����@����y��)_�f�W�����S�5L�)TK�HJ���/�N����5CL*���8��� 1���|�i`�)�i��y�e�k���{�tFs��o�������s��&|��{}��v�;;���l��4�@��`yM5	�4C2��&r\D�m���901���byfeR�>,����0�����˺��_g�մ�1���xs��$�K�W��1�h��ia�ω 3gb�*���˧[7�n��>��[?n}4�Ogg�E�951�>?{J��?�M��cO݈@kP�A������F�=;���`m0YwV��Y$�7��᳝[�ڹ$�V�T��I��%�򛯾�o�
l����w���g��,�|����y�2�^u~Es���c��	FL+��&��cAw�k7���~r��+5B����\��$6�=Jo�iIkO�g�1�5Fo5 Z3��a*�j���>( �g��������ǻ���͝��~�'��o~��9KvP�e/�^[�f:>�O��[a/-���=�V����8�r<���KR"�����ZQ`�^�dZ���%�	��yH�Lm������0��@"$��6�%I2B����' �ml�&?uX~`�DNB_I2D������%�%��8��MF��H+�??`������&G	���D8̙$�'@�Ζ��%_�a��,�p`�3a|�*`\���CO�k�Jm䕋��+S}�0l�$ר�� ��MR�0� #��� F��x����^��ǯ��O�~���&ZJ*/={��ʲ?x��f��o�������v��3b���#8%Lz�
+��_�%�Ԣ�9��������Kd������3��&��D^I����l�@j�G�_P�+�d�,�G�@( �& !j��H�0j�}���*�/Jf�+���`�Wa��~+*�@�0��~.��0~��f��W&�-���N�% d��'�ܯ�s��kd�@a������o� �j�GF�r�c�'�⭛��Y_Gw(�U5�6����.~�j��*v*Q� M�С����:2$+J�k�d��}ǁ���P��ރ�Āe�
*���(�6'�����j^v6����
�7;-����n`��������SL�����<��6֔��cm��Q�B��"!��p��Qq���-�}�%�r"a���*6��wBD��>�ӟ� �j�C��
�8�IΟ���#0r*�a�	��f!�I���l{�9�L��d�.ӊ��oy`������Ē)����K�L��I(�_��$�J 0�����%�@��,���)JN��h�3�'��	�T���O��̯�<� #$]&L���\�pd'~!Y��IJ�-�/MN�0�	��L��|&N�O^ ?���~~Y�_� ��)G���Đ--���!��A�rF�Q�y	��YI�L.�J2��QBnC'Ov4�rI��g���J8�&��-��K".�"
B!��'�%I�J:��93#*a���T$r��mh��T�X�?��^�UԐ����<6	(g����u�ڑ����sK���h��ٸi���آ�����[�q���g�k�:�{uqi���yq%�2c�����^]NC9Sz'H
6��(GX��N��"����._NK(�E���*�F��FEF��%_�r�2��d�T}��d�X�9A�����OO�(a�	�7u�((P�Z�;�R���mUZ�u��ۨ����Ӂ] 	�ayϑ�R9:m����e���]�t��}Z#S�Qi�����P�aQ� \�����Gl(���@R��>��l�*˘	}�ggo�H�1��h�#�FKy���/?���<}3
#��u�r!%e�(�l�",O���+1�φ�I�OQ��e���������	,��}B�C���T�!k��	DNO�y��m���{�����x�ܲ�y�lr���zw��u���e�+hraTC۶.&Ł��qv����X��?�?�w�n�]���U/Dx\f���.��J�EY�-BP���.앯X`��x��s�8�?�7�WlO��SeNķ���\��ѧnj�)��9�&zq~߉x&a�m4H�j=�����F�r��㑙����R!M�_{�ś��i�3�yF�wgנ�eGU5������v��=d�-�u��0{��U��Rk����Y�G��Y[4l�В��bcy�snv�^���w+�n4XJ��)����W��[���Ͱl���]/����Mo�8Э�(.��"Z;�2�;g�7e���I|��p���.��� Հ�����Ĵ�F�V��vo|���{pX��3U�4����kg�խ7����A��Î�G６��������7߾�K�U�����^�iq3� yHS���qa���m��Ӹ��ܱ��v�v�}��V;V��޻�==�y,�}ɢ�
��*U���rѦ�2�^�����Og��~9p��֭���2w��C�Ly�=�c�#H��S�(\��/�2W�q�Iq�U��H`��r�����Ĝ71�ٵd(�r�����{����z9�?5x��A�<#�LVϺ��"��3��L����ׯz�O/O���x��-��Vڬ���±�U�^�'�הְ.����ŵ��������ɡ���^;�+�؍;�v���3�"�Z
�|+:�}*�[�V3g��Eh�:G��ݓ����AǑ����	��eS�N:�e�� �[,��[�B��\���΄�AA�( ��$	υ��~�I���86�pQ��}|�����zi����h`����4��T�'{(����Y�6u�!��85q]/I��ߜ�/�U_W�kGCP��ٳ�^�hwl�l����T䖈ݭ���;�۫m�qc�`4��(uX@��IdJR+�ZCE>{����뗝���q��>l�������=OpV�����>.��.�{ [��=��=��09� �i
���0��	CFe5e���x�;d՘��!�[U�w�8Ի�>V���U�X�-�����v�A/�}�}�Ѡu~�����s��l�,��BX\��Y��R�hp�͓�p��		�K?-V�v4������CW:����i�9ŵ}�PgW�n�C��FC`x�)9�Kg�k�4�g�Z�n��r~��~iZ�i�|��j%VW	�J̐�3��XeB
�+.%�2��$8�Kf��	 ���7XT4l!��'3�iv4��6Ь��:�C-xX(H8��W1Rۅq�_��.����E��p�tĩ���O{�Ϯz�۬���ڬ��1�������Y&�Ĳ����`�����{�ý�cZQ�Z4[A�ѐ�����Ϣ�_��\6f��xU�Q9)?�����EmQ딻m�zGӡwVj�T�
C|�P�gԆ]`����.R>́�DT2!c%�S#�z� �aÙC�I8 ��7+��������[s��(.هb;�2uc�u�Z�[��N�L�&�ͬ!-���Ջg���F/3s����|�\k��*<N�Д�#Thu1�^Z�0l7�������`r2Y�MlΚ[ۍî�z�� �6�p�P�b��D�#��I����❫��?;n5?)���?_��@��QMc��mC�*:zZ*	~g��'��m;و��W��񐓊BS!`��&�ߍ�v�������_}}����5%����>�xk+V֚s�i&t�b8��a߄�TF3/�_��x`��ϕog�Fg����7yq�gΎV8�e�$~���b4�@8��lnu�[v7�{�;�;��ݎ{,�8 ��tl�1�	EY����M�c��Ŝ��i��Kb�o~r��*��_NK�@��钿���j��ޫ�g�Yǋ�k/�!�IFdz�٤����I|��1Y�}59���T?�q��I���_E�
�?�b��������f�S��!��|�������'cA.��.������6l�KB���k����]��&���ӋWO�_]��Q�{�<u|k
�h?�~��:�7��:H����7�%օ�N��co���!՘��.V�:fBa��Ɠ*��'/�����E���'�G��`��S�>0��F��l�_�_���k�s��2��ю����@�j��7=}��!5��a���k�X����5�v߈�;h.��x�ѦC��~�_h�����W��Iz�����e���O���Uxy�j���HVE�&��B�@:�1<��&b�����$�(n՟�O..��n�$�p|�w�R7�Z���6:���ݰ�lwSovgZ˼���n�?���+��$��Z8@�L�r�utz^*{��j7������N��7�f����f��^�^&B�)�{L�e�,$�ֈ]�&�Z8����.���%��Q�bB"�����:����g��M�V���9ب�⋯^?{5�_�j�Fee���w��|c��հ�K(������3;��JfΠ��I̡��FC#g����d>�8y�3�C}����V7����b"`����fA���ŏ��̷\���DY�IbבQ�ט�ezY�Z�����Ofק�٫�''V��a�ygky<ˀ''�����OW��x�98�u���$'|�#/� 90�XN)�����Q�� ���3��,0��`�|����'�x6_Q	��I�,�g�;�q�Ȭ����ÁA��b��S-K.�٢�g��7i3P�Ɖ�|%I�y<b9Q�*�����)�J�@n��&
� ?3�O���N0I�/D���o&D�p x������T4�������e|cj^8eɺ����K���rx"-�Sz�7��r�d�T� }Vu�D�p#���,H��NJ}���/_������ۿ���3ӀJ�\����cۢP���BP1�B�d]�����o�1U�4Hq���)ѣ �G��Ϟ=���D��7�I>ڭ�L&�����K%�@�٠���Wr|Q$A�o߶C���P*YH�,�)��<~��qY��	����)0���Z������TN$��������c5��t��*i�{r����;�[ІL4�_Ѷ8��N#`1zoX��6t�5�D�"����$r'�)���I[�Ō\��ˢ��k���B�d��LY�u�*���z΁S'�KB̈c2
�sֶⒽS@Ú�->�9�}�sr��{��k������9�s�"���JE{u�
�Ayы�վF��/?������)0��WF��O��~���ye�lE	,0��8�S��p�ˈX"�d*<)�(��)w.�
�Jr!�~�T��3$6���n����I�����]�~?53�C�TbM��.�H����" =p�p�dH��(I`�pQE��d`JƤ<�I@���_��+* '6�M�p
�� 	<(��B�B,? _�����o�n����ȊN�,��L�*K$�'�O`�tRA"�X��儐Z�#�I�zf�b\�f*��"����|C����AT�A��d����LҰ�4IVH+DB�ҏY��`��}3�,�/!�,���<;��J'�˅�(ꇵ/$٘� �R)�&�  l�ɢ%1�S.�B@�_8!%�K\��X�0���]g;V�U���r��[�;�п��ٛ8ƿ����~;�V�5������ջ���*��1�!�d�|t�M\u�.ͣg�I�F0�Mo�+����E���N-�Ɂ	������O1Y���$���~���<C$L��.H(@29���NL�0���V�����O�@�MR��I����U/����r�K��0�uoz5�my6�݋3ʨ�Z�B˳�x�ɖ����ݣ���残W�ӑkXfE��p��(��PhB�����\6 4s��)0I"
!��O�P"����
��_BQ�E��btΎ�#�K����[�<�2_8Z�G��8^m�O��PM�qX���cZ�������|�噳XO��=ntA@[4j��0+��q�"*�6���_/W-����"/����,z�������{��G��7�g������f�m�&1BI�`P�+����e���7���.������fߎ�K)s[���{a�I�.��V7�"<L&I��K��$��vМU 2x��� $��d"�l$�{������vc��'9�ۿ4�F�x���׾i��b�c�o�?���s���u���ɑ����]X�3�\(+�(�lF�W6��$zp�$�!8s.�b��\Ɵ��\��rew����m���>�u�⤗��-E�CeX��Hfr8cr���֑GR�Ô���������{�Kr��Y���ة�c�Ip�y=����,,4� ���Abfr;k'[8>��*�^��B0��훵
��ڻ	T�����nQ�W^���y�k������Ȉ޴��Һ�ƣ+���І&�.��o��zqq}:^�V��������M�$U��1ͪص1����ƕ�^����q��K=~t2�?�u�po���S�3�L ��2p#�$��z6e����L�Vw��f�����n�y5�>��n�F.iȬc�Sz����6̢�*���� L5���O6�ȷ�ĔX��	��B�,P��8�B��
}���d�]�O?��u��Bz�j��U =�ԚJ-�V���""�̘��.g/�]~���W㳾�S6q�ѐdm�6H����i��1{Ȧ=D��m�����hR?;�:=?99�}������nl�9��"�����ބf���Y"�F�n{0q2�;������������'��#�C3��>�&DѬ�S�)ь5QHHu�"�>���Zl$)�.j.W�H���x[��w�@b�+$���dN�T�%֕��{���Q��y�׏���F�P"ƅ�?�h������_��|3y}9�O}��9foY��!����\�I)\����,إ%����Ã��p�{��CK�~�~g��Z��@��1<����+Zȸ�hkC}f3n��}�����|[��F?1��=r����0�c� �b�B������+���}��T���wi�FO�$ !`ԑ)����a��d��ɶ^�d1��N0M��0 ��/���/[�x�i��������?{v�z����7���v9�"s���O]U<�[�Yh9V9G��fvx0�yq��<|o�s���7����o�;8C�ر�週uq�W¨I��T���|l��k^��{�L�����&+D������x#7�n���5�����;:"1-g� 8�ɟ!����d/9#V�X�$�9U` �V�w�փ�7�E\��s�.�&���s[(#%�^�g�c\3�i�K��x�睙���//��]d[��'��`�M''����{����.����u��k4vi����������͓����;�0Y�>طT�؋�5�\��
B/��^s�xM3�Yn�~��V������t٘9$�0�Ͳ�(�Ғ�
�    IDAT	��)�	W�df�X��MH��a#'��{�,xS�����Su߷��f�C����m�c��Q԰���UV�^�f��&յi�#������닧/.�6��͸7^zږ|L�)�bs�^;H��͋�t=��i���Z¬t�5ܚ�*�'�r��s���ɑ��T��)M�э����y��D?����X�\�l��o��;|��2v� ?@��LR�;��Ƚqۣ�fq �&Q��8��+ԔB��(_l��
�`��&�j�zS���D!6��I������ok��l�s��?�wp�5ޘ�9M����FL[>)����Ӊ���I���ͫ������f0��O��cv��C��v�\�n��AG���Rih���g�2��n�[;�;;{[G����[tW]�)�nX�쑾�'c�bi�]�5��ʣ)S/��^��g����__�֌a�FuǴ�_�LO�<\���{�F�b	A�<�<aR2�#н޽{W�i��^�g��*Z���O�J�@%�� �����t0��w�������uRM�C��G��ݾ�
@s1���ۻq�Zg	T6��ƦK&��f:����sh����a����7�'O.ݰ��V\��;�v�Ǧ�*��huX�A-菇����φ�a��8����i�@I~z��6'BL���g�B��u��!e��ꋁ��׭*S�[�'>2v�2Z�;L��Y��^���Bs�~�셳c��S�M&������w����&,>�ІcV'���d����m��������>���qΤ���~���W�!�ʈ{�o��������ƽsvG$4 k�F6�bp'�G!���,+���pl�~����R����ћ7� EOpH���q0��~���EU�<���*Y�7��:�M�;ӫ���p�aB{�8�K��x��vbzdoSI�~-&^��=;�Ӿy��u�����'��^_�����Ӕ�b��GË���aS'd*R��梀@��l��ˆ,�P�x����^I��������!�8I��Ǔɗ_~����Y�����r{�ӟ|r����r��j6곤a^�����nY�XĠ�J�X �����5Y�'�vXw;hu~en�zx�0��������mX�Ʋ�c�����.��|{;��-��Z�kF��y1�����U�w���8��+^wץ���n��ɟ���/�����WҎ�:ϯ/���𾺍��]q�6��vά�h�Xg�"7G�00^��Ʒ��"y��@�Q��w�D!n��"K�e��/�$�r�?  ��/$ E�̉���/*݆$?����)S_ ����!~f.r�Q?�I��*i&pC?�̝��Q��$c!�9i�	I���3K
�__Y�GB���̲��	9���@(�T�<RmB$ϟ��^2#�U��?&�D$<B�)_�:�L!D�/J�ohB����������i�刷F���L{,����mF:U��ؒ4����?'��o������_������e�<{�쫯�B�@�s"UT��>����$8Y��֭[�P(��H'�O{��rq��<y������1U��Ek�?ҥG��ǏaDU�<ld*0
l��n-j]/�#ݾ�PB6{�HG.0{�zf��eM�G����w��(�� �N��U����gV����E��� �$�-v�`=[��/h:����ރ;�����A��t=���<��"@ػ�2'ZLcI��8D�,����[���F&ŏC`$H�I���v�+z������)z�֟ŊN�CQ��7֔N�D����.V$B�i��h�i�c��m���j�#!�''z�h�8���jR痎	Yhi��F�c�f�%�B���E���%����wD�ój�d�d}���(���\`"߄�� I�&��N�z��B0~�|9?3G! ?��~�rB6N�,��"��T��&$=`�� ��t��4���I��J !~�瑵���,��f`�_N�� �GZ�8!�� f���]�_��L�#6Q�r��W80�����������J+$c3�D%$�@�4�0Vy3����4��(���O-��!��!C�"�o��-�~t�A���O�c§�RSd�ǆ�K����f�ďLS"2S��H�X� �9��(!Ъq���,a
��*X&��O��c6'�0���1�Ll�Y�1����
L��]��4yq�Dx"���W,��be��Tj�&ᓓB6���O���Gb�O�~'*�C�����$.�@�ꘘSM�m;:^)Y]XpԪ�WN3��Ljy}��	�n6�We�o�`P��Q p��|t��7텙�Z�����.�<�5�'W�t��(T�A\�7�ʃuY��F�!	� �W�qe�72I~�Xd^�j%%0���f�
@�Å�QZ.�R)~�A!@����U/��emW��[��>}����~��io�Z�ñg�z$�Z�+W�{,�f�|��}ԥ�YM᭑��M4<�� +Ad�|e�� ��O�,K�� *Óx?3\$�S#�B���Q�e�㾖�����������O������������ߵ�Xb<��{:�h��-��0ZC�&��t2臒嫯O�u��*�El4�;��ҍ��ks�dUvJ�l��EE���j�w�'��C�e��M-��C6�������^w���b�,����ʜe,go��.m�k�����X�*U�ON�������U��F�9U�u�d��B�f��7<��'�Z6f]`cr�w�[Q�f-��`x����'��8�����G���f�Uћ쐱uD?K���4��������p2�:��zxzꮏ��V��i�I+O��:l��ڕ.������O����"S�qǂ^�6������\MF{�m>:ܧZ88�e��`'&JQ.���4q����q}�e����z=>1o�n�ۥ�m}л}�ہ���r���DuX�wH"ƯW��ZIǥ����q�� AO�(Y��/���l�*E�E�plO�K�r&�-����,T���8Ӳ[[�ݺudh�:����qW�U�B���cU&�8>���؃[M�y�Z�ś����}?ǵ#��'9��0��9�޻ɻ��s*Wm=��i��_�+����zoT��Dr89s���ii�=��08�F�4�F�q�qp|��ؼq��_}���l�N�%u�Ⱥ�1�UP�8����Ԁ%}�v��?h�v�E3{qs�����Ξ�Or�	:��8`4��%2������l�W�Q�µ-�����y>h:W�
<�-/uW	�د/��!n��.���� F�(��",F[���700b���;����QFY�;l��L�t8Z�l�����ճ���U[:%r\$QH*�{h��8dE�bd�#�����^�{z��'�Qs4m�7�Õ
W�t@�觢�!���&��<ڪ�����s�g@YE��֫�<o�L�.n�x~������/�qF���PǪ!��+cO�b�륵�R�<w��������c�io��ey'�n3�4P�P؅���;٘a�g�[a��	Wq[��+&�YA~&ϕ�$Q���b�e�K�Xܠ=xz���[U��c��ݭH�BaS�D:�U�
���]�ͱ3!M^��fcpqֱr=�(���=�M� �a|��}�!�C�E����>�HD��	���nm�Wo�9�}���m����x �p�iu#�1e"���oDAx���82u^��w�s�zX~����_�\��S�Y���`c�nk�Ex"���{p�O�  F �5Ԭ�L"rQReud�L�Sz��:��;��Ϟl?�U�����0jU)EP��u���n���|�߽A�qݼ�>�p�$�3~_k��v�׭E�DP��q���h�Yl��-� �Ov��1����lw�F�����6�{í����6��5<�j>jux,����}���L���}<��q�]�+嵍�֨�1L1�~z�=~��R�OAd!U��|�>���J�wVG0�XL��<(����8���WV���~����-�c�f5�!�h�*�Q6-6۞��כ�(;�N���Q��{|eh��Ɯ�^�v��w33(���F����g�C�P�"ԟ�8W
������;�v�j�Uv�mm"g%C�_��#��q�t�;��I��{����p7t돫��/?�uZ��d0�66��<>xL� oP �ϊ�3!������Zx*���{��-�"�ϫoB��ǖ���dln���w_?zP)�=�,����J@G�p$�c�ܭ��\ӑ��X��l�?�{R?�L����Ewѭ]��-�-��.�	�_
O����e�9�(g��睬�l0�#1\���g�{��}�Ю�����VXJ�@��&�cT��O|������|�p���y�R����fgy��6k���]۶*�<7f"dIro�˃W����1?(��dH0��(�M̓�Yq �t�����u�����l�A;媁���{���2�ٌٖ�Q�Fzʫvb�4"��ȹ��4꭫Z���C����:���s^���H����18ᄻq:�K�a!�ޒ������f��i�5�[��[���W[��ߙ�Y�a�:���nOW]z�9JM��D�M4̛���V
���>�W��Sz������3�msW�[I�0�e�q�!�n�W�8i�M#��M��4�yT)�+��pjR29c��C�}$q�he���Q!������W/^�~���E�v0�{��?J�D���ب8�� ��@7���V��&��L�J��>4�����l�U;kј���ܪ\AM��2ϥ�QY5�7kե��m'ow���z�q����n>��h1����:��{�a�~3߹����3�}��o��t�_���e�)^y�4��gv�WV.w�mB:G�?X�<�����<�ֶ�)�z���z<q�x�m#/�TTq�v�W{���y��@J��|V{
iH�v������釷��w�.�ƓǏ���!?�	��� k&+<D̝u�`��e۱�K�һU�^~��_�.�75ך�t)�o���Ӧ��^)ӎ�nM5c�ߎ�YWV��L�_}S����r��o�,xco{˥k����N �(����T���zԚG�v��~xw;�һ���s���?��åQe���f�n��F�*����Bf����˵R-Y���ſ�Z)P��>��0� D4>���8�$��T	���9=����s}U�͜)���W�zs��n¿k����'74hM�̓�UT&��ܜ��v,���É����5~���M�ӏ����=���wO�����>�
�A0�`�\�7�Fjf������[[�;���=ĵ�����)���_�u�݆E�����n��2rk����ͺq�M��Zpr<�h����I�l���R��D�0����Ik���^�d]�}��l�j$XQH��Z�:���A�$�D����� ��ԧ�0#��H�T��0Vx@f3��� UFJ��5i��D"2i�`AD�d ��i�o��& z�a)�x� z<����E �H+2���U<l��䧄�H0�3�� -`�L띹x'�_�L̒��H2R��,�	3-Hu*#?=�
Ãϒde�U�|�)U"���k������n��
���޼ycC*��O`��}C=����|�O�����?�9<yZho�`cg�P(�T�����ɿ�ۿ}��wh��o�0[�FR��t�0����br9S���`W�Q�0 ��]z|||vv��Y+p���۷o߿/{ê� ����XYry���;�?��Jݦ�H�,��&�Q�_P���k��,�x�p~JI2^Zȕ�[<z|����(Ѻy�i��Φ� ��X���{���o~��~���r�4lZ�=�7�ǦK��%��T��k�1o4q��2���'���7RI�����l�_c8_�a&	S|�6�Tx���]J� ��EC�
5P,��8�J��2Fу1�0�ŐY5f�V���x#E��4�F22��r��������b�5�@�@��yc8j�����#D�V��&���G���x`�'�d �=�K6���DrI�`iQ�	��|-�!���,,� !�ܓۙVB00�r��'a��$@���	f)�G*ɡ�PL>�2�O�f.)y��wt1������ Xro�I��H�-Uf��M�g�����'LR(L&�Ad�T@����KX�~fL�3&��|�0��)a���#���ܳ`��~A `a�$�Az����W��{p@rL�A ����3���*`�zC������W�LB�	������]�Ȕ<&��ʬ��L+;E��#l��dl~����r�P J�Y�`$3�%RB`�I�'��V|`,�����e���)y��#��A"�༯R���@+S��T:�$���`	����� `�0�	�p!ȈV��T�NQ�T��P�
C���7����ۭ�����w��Љ[2�wZq�F���Q:����Zc�f�M�1ז�/_?{�x�:�f��?]��0E�ymh*�zZ;sFQ�F�'˅�~
(��2╘���2�/F�����Ȣ��9�|N H�Mx�3�-�0�L�x{$��46,��,�r�A���[�3:
�m��?k����o�}}����RoNC'�'g��rzh�@ݍ�=T��Zi�����|Ʌed����r�ƨU��ѐ��R$aI:�+�������d �� _=���'$�Y��Q-�Q��r�gu�����ɳ�zy\�۔F����W������JA��*�����n<uhmh���w����.�^�?'﮻�=�RW(�a��Y��Ɔ�M�=�'�������&Oȗv�各j� �k���C�Wd傐0��AH�	r:1#�N�R�J��<��C�ϒy�:w������� ��2�R��.�
��z�"�LK��d�l����
�$�����Ox�a��*��r��%�o~�ۯvg�4��ԙb��=&[s*}̉T<��s���<�o�U��^]�pu��u~�=�w�w��Ѽ[ZmO��~�+�-f�8�����c����	k��]�3����U�X��7Ա�n&�3/s��3Z,��wn��G�hYa�nw�����ry�zq�)�ujj���~��~�u?u�A�0ax`K�
����²/� i S�78V<9jdg�0���KL,U*ܬB�'cC�*z����o޼zugs�_��u�B0E7#d�م�A�+=����a�q���A�_Կ��vt�{5��9~���dv�!C�[.����($����>��-��f��XB�Q*�%ԮZ��H#Q)u�8;{��n;w�^"f��Ģ�4��H*/���ؙ:�8iͻu7�������=Y�Ŧ.1O�o�T0�(]�05Æ'�K�m8&�і��_3|֔Tb�����vw�F�������Փ�����R�H��yE��1|��7vġm�2琄�u\�~��s�,��'�y�-h˫!iG�Jo�^�EE�Y5�j1�}��*�	=��얩�L�+Ey���u��F�.$��c���$�C��+$j`a�ZXrލ�,@�˛�L�6W]L��@�˖��v��	���$�}���!Y]!o��d&�%����I�# ��$X�]��ϼ�ڍ�^[���/~���m���LK�ۤ�ۈ�q�cSϏ�a��]�㖨p`}��u���������_��8m�.��͠e�s3�Q7�,3���*s4��[	zF҅}�+��ׁp^6����ُ��cg���6��dڎՒH�؁RuB,⿐6���X�2
]������A2ť��tsXdN��`n㘄��L�L�J ���g��E�#R���S���,�v6oY|��������^?����z����=�����m�6��0�~z��8�rټ8���_�ޞ��]9IB�L���A�j��M�֐�L8�s�R�ҀIf��R9����D�=�������1.�;s�����LP21Є�<v.�y����ȏ��Ů��|�/��rk�k�[7|>;�EayR�V ��.6*Y6��9TQ��
3��䬂d�$�L���~&��2`��� �@�����W/=yrx���]nk:��Ρ��2�f��    IDAT�M�Ry����t����?��Ij7�W��]���9q�3�D.A=ä"�0uC͊me���`etp� Af��pd�t⚷P�O2Xb`�#m��l�rÇ�-��%���*W�v7��J�A�ղ�=A�2�R$�J�	�@\�ટx���F��frI��b��zG�K��d@��&�;�M�����/�~��p��9��&z�"j�19��a��g�m��ۻ:�~���|s��E�c�5_�s1�^nY�p�Y�6��>%㘧�[p>&�9厽85JUd�ax�U�m$#��\D�ب�P�v�H�h'N�Jc��!��k�Pe:o���y�Ӱ�2*O/	j�\I|�@�o;��
B��@��Xt�N��˄�^�f��k�h9L=h��'��A�Ę�u[��w��v�T˛������Ƿ�e��_���:D$���P�ƹdr��R�I6�j�Z�~qY?�>~_��ǫ�W��n�GS9m��!����Ew�K� Fw2��Fu�G;�f��m:h:7�a��p��o��O'�}0�?�\q;�IwA�#b�æ��*L-�i�=n���&��[[�+�J��l��g�'����6����j�L�l��I�Cq�\4~aoJ]��T��&���`!�F���^<��z�r c���԰=�4EgggN�P��r���;�_=�w�S���C�:%fk�%��F�0�ĝ����X�����_���۫?zr�y��^������Շ��fw4p�:���ÅeN8_�Н|��#F�},E�]V��r�4]���_ֵ��mzM+,H�Y�3�X��6��|/�̈����%ƺ#�F��Zүu�v_Ʊ���RF���˔��#�l0�DJh_1�9u3"�D���´d�c�Ƭ��x���˗�ҩ�)ZtLc�P�U5Aex�o���ѷ�t�5�0�v�������w�m����2o��[���g�/*�XVĢ����Χ��Ggͫ��[ӉY;�$���m#+%+	f�$��W�x�3��(�Q���lh�Ӡ˂��N��s�r��b*����/[�� ���^�V�,'\�������\��7��KT�^r�.U��q�7�e�
�ggW,,J6j�����`��'?�����0�k�.��&G�@Ky��ٶ�u��>r�G�G��N�r�淿x��ߎ���/tK���$�b�d��!�/��\�[��F��o�v]k<���>���gb���B�d��?��DB��ذ��Us�������M�]�n�>h�y�)΂ƴ(�7I�{�!�DN�r47r�lP�#�'��Y�G����4YM,O�;�{k��]~�#��F+�z�WME�"�+��?q0: $cEJ�H�h>+N���,���I����0Qy{D��SX �Fax�=�)<"Af���l1`t�,�xx&ӊɼ9���[���$ޙW���0h=	�x�|�r�~By����S���������)��� �R/ ��-�o&�G |F&�����O��Ll9���$�~
K�YH%�Za�p�dA2m ho��`}��@/�VC�H'ONNt�?���7C������,��$-��W_}@�;��L�U����z;�	�,0��&�٣���($����(azl4 ���H���Jۤ�^�HR�aOgK��?�CJC���/��j҃8��f����=8Ɣ�����r�Ch���o�Uf,��qt'��UL�^��y� �Oo b����?�����	o%�6�l��v�b��(mnl�x�������?ؿ�VC���!�����!�~�������3������ �-|e��)n�!�b:cl��p���8�HҾ����v ��r �IҌu1ݵ9�7���g<�w������T�@DBCu�S��-賓�b�~���σ��H�����
�e��W,���*�J�����*�V#�๪�Z���y <���^��+FBo��Q_ދO�G�0g��Y�"&� �O��Lz���)��YJ(���D�_��xT�3Ȍ�6ao�I�2af )�"��F|&�^$����b���6z���-����HsR�a�2�ؒ_�{�?�[X�$ ����@�Lr	�H��4�$��1�g��@�6��?�&pҟ�&aI0�� �P p���2�I��Lɛ���� 0}�L��@�h��ϑ ��&/������L���"��!	s~���$���$�[���f�d$,S���O���cI6�lc�����0r�bP(p>��d������7���x��F$,n,��sI ����	x��\�B�GZ�)�P�-�`i�S&�P@�$���\R_	����SV��(�>+%+Gé����2�騵29V��H�t��߉��÷�L�[��i5G|��\���N�e��L�򛕻������vy��eFV,V�/��e�B���	ڬ��$�����.8A)�'YF1~�č���.�5�,(�+{6T��J�Qb-�x���+H���;c|�*�,DJ �ޒ�PT�qz0|�[T��҄��u�Z��Go�ߝwN���]Lj�i�"��P�[h��@a��e�h7�n��C3ZP~��+�ʵ�
��F>��=W���D�a��@�4'�H �H(y��S&�Aؓ� �\bhHS|��޽����g�;�2GVq1����{�pj�%n�
�-�P��]c9�}օs��4����ۋ�IwR�\�M3�r8���S'������<��q�
@v�V����:��N���������`��a�p�b;Z,2c�A���@�,���&�7&��ɦwu}����ڹX����iL�tV�ޏ<ul��X�.م����J�f����E��Di��~Q<����΁P�MuzR��w��������Ҹ]���V���3��&��Xs�4ks9ju;��󏍓���E���Ʃӝ�rgV��vseܦ��Ӱ�9t���c�Mɭ�T�H-H
{p_�j�x!�T37g}פ�qf���J�N��E<U���$X[Y��.�	*�(���Shzw�:9G�&���`^j���QT;���W�d&�=4���`ƪIo����d���~��I�����B q��W�:xe� j�t���_�����ʦ!Z�\(�Ь��rb���q�Ҹ��ʭ�����o?�?6��ӓ��[��j�?�[u��
�u,o�ӄ�I�W4���G���n�Y�S�2���%�n2�;M��+M����1�r��ES.�R5S,�!�$�S������������ȍ�v\���u�c=ξq,��1NS���'�����<L�'{UG^$̷�� �����L&��
�ͭ;����oo�v��8V����%��3Z
�{l�+J���_�z�kkW��ּ|^ou҉!��1�5�fc�Td���d��_CNV�~�]w�E���X ,�͏X�7 �K�M�('[Z����;
�*��ЂO�����;!�G����6��,���RY��'�㠱%9S��)�Z��'�c�BC���Z��lQ,m&��W�,���V\ص�����j�[k��$��!B$���4+�%�<Z����X>qi�ѻnh��ߞ���"9��M.�^)^��и��90��&�c��/vs���TtT�:N�;���W��!{;ԓ�a��x�iغ�õ�i1O�B�IYѧ�b�:��L��9�bȜ���
���5�C��|�Xԁ�՜a�ˬ�P�d�ĜL�E.8rѪ�z�������ZTMV$����l������9��˓��׌�^��q;��zڛ�(���\���4��M�Q;���Oo߽k~8�^�Ä���4�2c�S��'�by�� &��2Q�Е/G���b�a2V��u�.�#�Kt���s"��� Ķ"�KYn\�(�ȕj0�� >����~��n�/\���.1�������d��������I΃��Ixo �Ĝ$��H�}�?�/��^]٨�޾��7�=ا��v�l�q�������P��i�;nM�x	���W���[ߝu>6�W���N<X�j[�l�)���.
��IL�<%�	�.��=F����q�n�6��64�C�y};�h ���Q1b+��@|5*2�1�P�c����P�q����ft�%�h�V�5`�(9�EEO���?E"YN.ڰ�"'�5Ԝ'���D�a�$���*?Nv=}��_����u]�~U(t��`�a1G�9`hJ0�>|�Wo;Q��wg�}h~[��F�a�I1��2��L�9�dܼ�V$�'�8ɻ����X�F���D�i�Y{�F [�6f?�G�vƞA�`�&��q�_���>7�r(���h����͝�U�z�V���	C:��u U�߄ݽ��p�@<Ɠ4e��I��3��~��O<��锡����I�x��8��M:�g.O��7�.8tz��׿|���a��� fj1��}(��Ѓ��PHLGҵ/��.�>�pq��v���ۮI4t¡�ؚz8:H�Z��m�䱙˞O![�E�+:{<�����a�e�'LN,��Gw��6-�L����r�`��(�ߥZ�;Z���o5���!j��s����]~WK��⿁��.VС�I	Lj���Z�j�����^<x�����ζ^�0���������o��8��v�?������hiس��q�r�SKF�1e�G��;���V�5�/O�?���;�|�q���+�8��G~i��tR�.�Aq��Abp�=c!�ܴ��xh�6ύ]���B����e��0�O�͔�>%�IvNà a�<�i���������$�9x�=(M�Z��y�_���f<<�����mU�ˎD+\8�0Q�IL2W�p3̾�l�FcY�R��0��yLN]7��!J�G��6I���N��~����H�aCc����޼��Y��`���a�VG|c]al�3���u�p��l�+k.ܧ~���'���xѾ�N�{�?1�/s�jހA6�I�b���ﭝ�
�Jl�Z,j�1��j���c7�=�j��Pdk�(v��~��1I�UA��f����H�𻻕�z�S}�g�WU/�8�[���p�]��P�yR��1�@F@�7E��-`!���!��ӧ�4r�l 4��DQI}�pt���l�^��Y��������J��5/52K4�"7�\k7�U��%�Ӓ��y�v��h]�ꨟ�7>~j�=����؄VS#C-O�h��j����i�aQN9q��ʱr���ֱY��]ν�UӯQ�cg�}C��F�qA��R8a�e6��!N����زK	lp�q�af1d`ï��iլe9(��˄9y�?b��d�j�f�h��Q)��;�Jb�Q)�&�&�Z�,���z�2�
�x�K" �ןf*2[�D&iQ+\���Q�3� ȴ	槌 �$�L8i�"�p�K
�L�,x�����Gv�D�h�0���g&L`	�J�K�˴:2p����J��"U�Z$0�~J�I&��$3�'		�;�$mf�Fv ��0o?��D�O��G�0�� zq"�*(�U_���@���i�A�J�Ղc��'''�v��9�U����>|��͛7f9�F0�5��(�����;	��"ȗ�W�$�
ɿ�˿8�dS���mJ4C�%�a��(~�P�Չ�T�S���qL��#�/�K3��`��������/^�Du���ׯ�Ib�����]�2ъ�}���|'���b|U�I�#�O-Lր53�R=(&�O�8��;[�<mol[2YN�oߺ��/~��_�:�C/[
EW�l�kT���$�5<��õx3�
�?�e<�M:��2/�f�,B�c�Ӣ̗C-�>������nX�������]��#��s�P�(����bU�g��^
F��Yf���@���V�r�!��q�Rh�!�LHP����[2f�L&G�^X�8w�o3���p��	�q�D&�;�g����1d�n�,��m����#��q|Cb<Hʞ�v$Ϻ�0�@Xti�)&�x�U�H��ޢK�A  ��/����H���Kj�>�MN�$�H��&I.~�֓8��WI�<�J��~!����e3��}A���$eBo�"���P}<����S*1"a�3�Ͼ#S8}Z�)�L%^X��3)\�H(�m^6O�
�G�`�x b>��L���[|�/�����ɊH��Q~"}��S��'����D\��O���0���O�
a)���{ȟ�KE�P�71�&6o,�H"w�d�h�L%�5[��SY2!`xr,!�<�Up%L� ��R|��CŬ��& �)jZ��6�Ce��U*�%I$���w���gI����r��Z��d 01�&6?!��z�7-I�¤�J�	�X[���0�L,�)d5oE�������Ae��Vsd�eb�ﷇ|ϵ�7��tzO֝t�f�۷n�x��ׯn����sKI��a����9�a;�E��D9$�Ԣ	g���'ċ��G�$� qCf��ģ	e��I�`�����d`"Qג�I |��/�@����*�'�FaD��e���fenW����N[g�W;�g�TF|��PJ�r��/*��;�E#]��fyNb�&_aYU�i�=ފS�d'g���-V8��w2d��1��	m�G"�U�<�&2A�>�����'Ϸ6��v�NB�����Pbsi�*i���7F8�����p���U�u|�9�M7n���O���Ee����}�9��b�^�Y���Կ�ź�A�EA���t�Ҟ�����*�?��7̹�3�v��>eN12&������nQH0W�YW����P�ZSV�V�`W'��E�;gKj��|�Ƨ`��l��d vᶺH��y,�u$>?������dH����(oXܙ/�˛���~����tܜ�]și����GT0�'ޅ�΍K�~�׹���������i���w�N{�2��4]V�;:������h
�d�<Q���FDf�d��V1�����Xsz�>�����v��w��ex�}sF��b4��u�.��ܘCC��r-]��]F��U�ҐF��5,QoqJT!u�~Q���1��6*����g?<Zx>b^�潡�g±R-��+ӵe&�{��{����J�M����%y�3����tYzW���ye���n�vV��c��ԙ~ޜ����B�hզ	1���mx�E��m�D��`,�c4�2b���1aσ��QEw��5��x�'Of�7�#�f�TEő�k:�	˕P�g������0/������ze��^�cZsUbWQx�&�'��rM/�T0Y ���	U�c��? �S*��|����X;�̜ߞ�z�y���յ�]Gc��WO6n�`�E�ʲ�����N��<*w��ԯ���{<���և��?�ױ�"b��R�=-�X������r���uR���p�4��;E�:�C�/�^�E�&(/,���?7n��߿f\�8}���#���%J��~����@��X>lnUV�3v+|�9˸D���l��5�w�+��'5Q��$'�z�$�Z��%Ix``ċ�'!�ʴ_[#.�s��͒�Ϟ�⫇;N��{��z�bd��#M�&�U��}�x0��O�����U��ݏg߿���mػ��8�mY<tR6����Q�W�B]������ը>%!������	��\�J��w�%AɱV�(�&cJT���8
!,R�`v���h�%�'�ik0��me�~�_��%8\�=��̇���"�#&�ӂr�#��"������+\;:#K�-S���ݭ�Ow����` UL�`BH�[/!M�
�wG�f�Ӻ�T{����Q�ѿ�"ue�;)1�2s���/^�f.�AV|T�d�R����o#��Ӑ�em��E�96ɀr�WA����dkG�J8f�AԠSh�C?���ݠf�������:�;W�˦��-Hc�k�W�1���Pq{}�SXE��yY��?5!��v��߸Y�m�oo8i�t������C~#�>��&�0*��ch�y���!���=�|j~�}z�����_����r�Y�(k��a�Z.qa/���8K>4]P���O�(JHK�9�8��M���<��8g�juF�    IDAT{:��@�n�\[�E1��<�)q�m�(`(9�֊<���q��ڨ��q�v��Tq%���c��4*�����!�0��K`�G�7�xc�@�lWY�6�Dq��en�q����_����p���H���c:E�O��`R�s�#����Wﾭ}s�8b�G�6��\�5�{���.�B��,�]��T8�I�AatgC_��1ԜIWi��qO��_ݬ�V���ڤ��g�Avқ���y����i��4i *@տM;�Q��X�����9�B*2:Q���$����!k��8Y�/�֌y��z��@��H��4�ɤٸ<���~����_���!^�����m�Ĺ��_4��/�X(�nL�]+<��e���;Kێf^��^�[9�ϻ=�9�>���h��C9�"�m%7�v��$�2� �f��5;�ђ�S~�7ĹW1u���͚6�|��E����E5��r=p����b��ꦽ�8[��z��J r���������,#�Z�0b�'�ҶLb��䉡�ހru�|�&��x�p�Z�R�#"�ZMEi
���o��������?���}�����wͧn��qdhic��P�0����fR�Q˅��f������<�wϝ�4�i_�2�JG��[����W�U�9y�:c�ʺz%7_s��l��!ř[���E�y۴g�)�Pt�����.�a�1��Р9�f��,[MWq���k����w��3�@��*�G�w�;�;ش��k��`:xx��t>$�
�
��+���nL5lL3�ӭ?��]��
t-���;_jn�o������qe�{�%�g�����y�=l�(s�5����n��� �������={��޷�>6>44�0"���T��)\�����1�1��T�hI;�X%��m��q���������ɍ�X���om E!: S
��k��XO����3I���ֲ���(��'��y�q����_MZ�pm[Hi-m���̖��s�"2&��Š�ۤ���m����S�ϊ#0du 1ѢQ��y���OG���O�YO�8����߿ٿs��iP��gE����,���Z��1�?KMg��di��Z���O���?�teVzQ�=wL�L�^f�� F���Ч�ImWЅZ5Z{ث�xv}[+
�2w�M�![�V匩X"�p��8�.h	aO{$�t.�)p�����t�L�+���\-ϻrxؒ&�qtd8�Aa2��/'���'��,����Om;�XS��	�N���m曟� �a��)0��$��B"s�Ӵ0 ��z���ل3��# ���j����������I�"!<j�/ %	�$�<��x�'%b Gd��#�� ��w�%p<��� �dFP%�E�@#��HI�u�*?�f1 �� ��) �'�T\�|B�OYS��2  	xo���\����Y�?==e���{یt��ￗ
�O?���MG��
���"}"娠�w8à�ŋ�X:���$���a)#�f��#C�ܚ����p����������ۃt��`_}����w�벍���"��e^���Kɲ$�:g��&k�.#4B͇Ї�
if��ޤ�Az�Q���?��u�R!�ό��- Y��J��V�j+�F���v�*X_�2�=��Z���8�=|����W�0tÔƪ���n�h">�<ƘHnFϱ  mI��E�(�`��D�a�c��W�l�{5CG��h��	�Y&&mSVٙU�^�Q+J�{tNT(WhC)�"�x��3��v�6'���0�ifq�A+�&y3�`);MͽY����)��b���˖��͵*�{K�7�����O��7c�� M����aѦXA��e�f�]��5����DLF*���� �$a�g���L��g��Ⓦ�E�LJ�$r_#e�V|���9�MJ�)!o	��#��>ed�,ғ�$�W�!�v����C�)���z0x��Ua�uL��*R	3�,�O`,��&WЖ��
�Y	�6�ͼ�`d�ڌ�������ĉ�D"�,����,$I����T�� �O0��, �[��h��D�%%0��d��'�G8��F-9�o�J$A��I�$r��y�%IK��.�HE�U�;9��'�<Y(o_�$�`]JT�1's~⡄,<���O]���R�fE0B�z���D�xeL��Ic��)_}Ib+��J�4/� e��F�\�e�y�q C�d#΀�5���B�Z$ycf����CR+�Hie�0 4�# ��xO�(�X*L.�]�A�MV�����>�����w�,U��n�:oO;�+���܈H��+�v���8ڬl�����/n���8t�`DS%̸[�����c��f晴�yʂ�{c�G���b�,� ���?~z���A�����N<v�O0�1���=�7�`D"�BĀ��0Շ��:	μ��5�=�Y�B�']w��������Q�q{0m���T9,�,WC�-�"�:I}��t).�h6�cco�z�I�i��v�t�Q.���[Yezނ!�Y�'3&��H?1J�Aأ8~��	��'�b������@��hJN���xx�����TW{K�np��G�x�x/�Mq�Щ^>�
���ɠsq�:9�]�f���y{vR�7{L���]T����E#㊓X�+Vl�KK�qӝ-&b�Q�h9���jW�����y�t��F���6Y�X^.�)��f|����X�ڰc��6�)K���y�c�=v%J������TZfX6�`˗��P���(I�Ra��M��|���b�J���V�����er��d�*;���Xc[�fS�
��I蛦�"o7�̍�[��O��'�����B���:�<ScA�)��`a!Ct"������W�����#ԕ�yq���WE�������ٮY���L19sR%��1��Q�	Ͳ�f�۳�Pl?*?ysp�q��߬߮�f��!�i����A��Й����A0 ?��� ���X�.��@�1fN�>x���ݽ5;�w��������H�.V�f��sl7����ק�?��.�����M��G��|J?����O�H�U�E�G @��i�˕�L�)��Xavz�F�[�����8�7���kvթ��I�7��`u.&�5����$Ȕ�����ビ�E{�_.]�66n�ݜ������"��&� I�<4�,T� �F�Ph��*�� `(c�X����<X���m8���z����[�y�3A�M�щF�Sr\�)z��r��}cv���x������{y/�ۆY�Ί����2b�� tf3s���+V�H8��U�7:�BJ�b�(k�\R��0�W��;�Χ=XE�[5+��8�-oP���B3E��Ba���Q��ʐ�Ӹ�,�0�������~r5v�릜{,.���±v�1)O�㹟�?m�?����w�U^�'k��r�m}�l����Ê�(]��!PC�y�����%�����{.�tMQ��r8��O�{��Zn̗ۤ�\�0u|�v�`�2��ŀPc�$��	(�z�b��]v�#�UZp��M�����Zo��c�C�`�e��ȷ{�>�8lolכ��Կa˯A\"9���1�����y����/W�2���~���d</�9 	=��A�z/�&�yg|���r_S��� kJ��*�z$]�%%����ۿ��Kg6�ʦJ��I�^�OBD[V����xj!
G�x�!�Z�q�x������ѿ亝��Qy8�(m�@���r�GD�P-�G�x�=���AH�®mqF�;���g�Ѩ�h_՚��L^^��Tq*����'�<'��Sp<\Ì!�޹z����gWG��v��&U�5.&�J�Sq)�'��}R�7y%c� �	��x0���,x[h0���r��t��s3�W���`��\'_��¥���ea,�y���΀}��{��߻�]ޞv<o_8Ne�J� �y	c.�:���E�k��a��gs�.�;��Ŵ�
�1��\��N��:�cc�� k;����a�ԯ�ݠ�D�����5�<!�4�e�UC��K��v�5nW��V�p��HW��@�<�����˦��"i�:��Yi���T"I���'�T�?�]ucߝ��nTt���xF)*f}�MC�pN� �,Y׮_���~j��������ޤfu]�M���z�y&�:���G�?����$1Ȗ���Z{Cv�F�T�6_鍆���cw�V��܋��X&�QNU�k� �6{T�d��1r�ѕ�E�{?���åF��p�Y�����L����?�C��d_�K��M ������${sՀ�zS|�VQ�쓉\�qTo̝�������������{�^=ٌmn�KL�Z`��m�c�ZR=d���5kg���o�5K׃�e�V8�&&q��6D�U�@ף��߄��㠽��V�.���{I�#��D�1R@��'�e�ư7i��7mI,��mTϖ���'5ZP�&:�8J]㡓CF&¥u⑳���3��A{�w�7{��PX1��4��1���EE̚4-3�ES�6�� ��#FI=x���0��P�����[�2�6�u�G~!Wc�6�	f��,x�rK˸Qk�ڧ�=~h���-�mrE�qB��Ć�,�L¬�S�ѝ��ZJ�d�ye�P���)V����ݭm���k��q���&ym�3�g���Ќ�J��ӌ�6���(<����Sw��6Y�J��24�ll ̐R&�;F�3)ԭv5c}e8E&+�z�W�V@Ձվ�w0��`����Dt��\#��4w�4ܯ�<��ޞ�\��5�SFY�
��$s��,�`��l���O͏�O/;����r]1�X��9�c�A�"#I�)��P����%Eg�٠E��Z��ڊ�(N�o��F��;��i�s͕��X����^f��aL�:Y���1���GO߼�^��zvp�{�;�a�9��ݜ��Kv�T�xc2f�`�=HE$
1V �R<�ÓL΄ ��X��Zl,�;�
�KÕ���O_>�=<�kU���bX�!��$�WM���Ôp�U�j'�'�O׭�F�����LǷg�ۥ��'卣�1�}y�/q��hN�P���Cp2Ů��dN�E	��\1������#^���������smf�:_��k)�)ϕnԻah_����ݶ��Z���K�A�vqI���=�OŜ$��ڇn���N�#�lD���`x,��`�O�"�,؞��H*�hs?����#q&X�",���ӓ5�?3w�2�!Ioa|��O/ҳ�Z�Ѯ���%#�GZ�*/�$�-0�|J�x�) �wf��#2�fZx�$��%?}�'�N�.R�M �< �ZRx��GL �$��C����A��GFؒ0!��$�7�����J����O0 C��J�A9���"�x�h�#U��|��Gk-�����R������0�'������I
1��=�x@w��F�#���tB���z\gd!x�5!C�w*i�C.���/:b-�V?;�Tt�OaP)�G�x�B��t� r�������C^9Q,R���#�1��w�ܴ��H�#��f���Ϭ�r�����"L ?anQIf���H�(4Z�Sskk�B-��<��/������ؽY}+0#��/a5"�Э�� �AC��NU?���OF��	��7i���
���Uq$A0�J��%�;��M�+�
�O�S�6��w.���#CD@@��P��mJV)vai�ɣp܅oPP�؊5Z��v!�YZ���DUg`�޴k�B�ۻ\Ol�l�,Uw+�����7�{rZC?�(�X�4�4͘���}Q:%��Gˑ�|pb�J��dPGb���IA���i �`%�T�H ��� #�{�����U@�K<�rO��NH����EXLF�-1�a&�W��$2���Z�xo�2m� �<L��3�C!X�GZ���x$)��Cb�6�z���7e�I �E)2�|��`O"DI&I0ad��Xo������T����'�6I�,��W���\X���zK����ϟ�1�Ґ����E$��I_�Q"�L2O�a�g��гv��\<R�0�(a"1+��t���xr�5�@��Y�B-�,��P�-Xr�J�����I�<�6����$��@�J�T�����"��0 �L�Aa�2���&�A�*	$��-G8�<Lfy� $b|�� ��q�NH3�d@���������b�fjA�Y�!l�L�R�,�g�g��ʰ��������f�6��t|�WMMSm�=�����݃7����ׯ_=���Qv�58�#״����k�9�R��Z�PR'�I���{Db23���$8[�",� '��O�j$�h}�d��xa�O3J�Ra)<�`�P~��d��� �U��\�ܫz{���땭�j��vzt��Rh��\�����1�/4@�?1ұ�2lT�����������f��>WM4���(��u~���w\��N$!槥F�}��p6��D��
��#����[=$7Bc�L7���c³�w�n������8,�bH�������[Z��q���x��m�kt��fc�3��g˟F��}ry��~����q��RE�R`/:��hO�U����66���J�^���� �J�����U�[�p��,�ʒmB�F�,m: K	o'}|V����Ӵ�[]E�Q�}�{�`��CqV���Y_Qji(\�ȱ�����d������ 	��0�k�q'��2�)��ʈ��ȥ�q�-VX/�">���sMG=^�y��.:��N�v����r6?c���I�S�rke��$��$��H��P8/&���j�I��.��tl��D�(+�Ve�|��U.��k�l���bH�d�b���:a�ƃ����p�����;g+]6�sG9�1�c��a���R���>s�� �[�-  ���f�eԋ�~�EF6��z#����~t�����յـ�6-ü@���\�V�MM�@���Io�s_Q��hՎ���Ev2�^�f�<� ��&3Mz�M�&��V��x�B�
�s�Z5;��g*��ͯ]_��wW�i4��'���I��݉K%�Wŷ-�w�!�Д�zר׋���|��}�`������j���~�N{1�`I��lL?Ѐ]ɱl"Qn�P4a 4+����f#^�t�+R���D�D�9Ҝ'��͝��޽m/��f�|`&�B*t�Njƞ��w��}�������Ykt�V�ALQ� ���fԊ!&�W-�G��Yi�I���xאL�SW��Ŕ��7'�S򎎺��)�����u����[S���M�f��)33��|��wqz>�S��mVv��=iޮ�V��Q/�ۮ�a�Nf&o�Y�w�[�
����y
�H����_f�DG�NL�'�/��>��,S��ܩ�8�N�MF6$�������̝fsR�^�0?a��\^�/꓆CzK+-���U���Ic��)J�B3�B�g6_щB�E��n�Q��Ҩ[�ӛ��ha���n�ۦ��F�v�
��f����S5q,R�c1F8�o�e�o�|����sx>��V:T��Rt�PIK�Kx{��aģP$H�͚�w�b �%�e�3zh�h�
ⱇLŪ\���}�`�i1��'��� ��fٕ��
�,��V��e�.=�8~W?���pջ�-�R�k�,�/U���P�mdG��F�����
�,��X7|~��8V�a��p���7�ev.�y|j��!U�lSЈl8�n��/��b�"v��m�CǅĒO�'kK[��n�<|r��|P;l��)���fH�!_m	�3�,�m޸���n\�0>��X*�y$�r���8d����Hͬݽ{���Ƿnm�GQ���,9Դ��jID�v�]���-Z�Ƨ���?�t/�̴I/��L�"�cBbf�7�FCX�a�BQK�*4����C�����@(�����l!:��j�����.9��uww6'���`
��Lx��}�x�pG�-D�v5֗��w����i�qm4�W;7�8��ML
٣�.$��A��=�6�}�-�� �`��hKYwS�Ns�X�h���    IDATn�x�do��ݽv�M�b/$�
q�"�ɬ`О���u�ON߿k~<�u��WE�K=�[yb*��x�g���u���Y"D"ςK�'�Ϥ76HB����&/'���t}��T7*��|I���OK��M�[t���=���+��������՝�����_[7�t�1�r���!��p̑�O(���'
��;JU̯,��={f�i����Dk)�lQ���A���s.���g'�[�[�^>}p{��:�QH�0Գ#d�2��]L�hW�%GZ�ns���b{|ҹn�/:�ΠF�ϫ����zl[�V��lFJ���F�!u�*���XS3�0�8����=s0�u�˻	�k,���U�vY�vL���Z�}^l�(��힆��T�"���V��`p�����Ԇ��Mg6�V׍���&��86o3��Bag�7�� &��[tF�m�bc$%7p!j� XtLU��0Ho������S�onzx��٫���<�N��$|08z�j�p��102�ǓA�M��N��S����ĕ�s�m��3��B��4-�q��@ �Z�G�t6�PY�R�F|��[;7�+����O����f�*�F��D,U���KU�W���U�b�n�ރ���O�Vm�Y�5��bhrX����K<'TU�5]��:͉��L;Qo��s��.[��R�������_���*T
���/?]��[�q�|��?��`�]�o����*l\��	>���D��#`���;�������h���:��[E��UeQßW��0�'G9
��h�Z�ƯlnX�[�L���v��a?��(!16�B���H�'z}�q8�h�m�������Yg1%{t�黫���C�jw��;����ͭ�3^�5S��(I�b��㧶-��b���v0ڌ����ר�\~Z҄I��b&&q�^�9��s����?zqo��ڻ�3��[F|!:�q8H/6_~s��
"W���ը5O���z���6�
/	��l܋�á*g��mo�|	�Z�d���m�Ej�
��&��&��F��1��^^���n��I	ø��\r�K��zx�Y!oC��
��������	!��_���������Yy��f3��X��l��!5Nb�1��j'��$�����s�_��乀��*X��wVkV���5+W8�Q�ޙV ��)IJQ�&~�J�TP���E
/���E��d��$Ur E�����=��h�]�<�gF~Z�J���I���->!��Oh�F��$I �e�!��Ѡ\9�J�3~�h%Ϟ�p����L3�-�7<�U�,��"R|���b$� U�L�=I�����Ħ8_m�'*`��:�7�(�!%�T�˗/�_��o����C�W�ߧ�I.@��"G-KU�MJkvd�iN���6C���7o��ۿ}�V��D" �&T��������\�ﷲɞ,�]��ϟcAF��C�2�����n0.�Ĥ^�ɓ'b�	<��A��Ǐ�������k%�������Y��B({0%�'�p��$��l�(ɀ,D���Y����o�sQ
��������ׯ���ٽ=�EZ�ِ=���m��ӦB�I���Jhǂ6��L�H�/K��B��@���EAVۣ'�?x�,���dx�w��4�����-�2�G9�&��>�;@ʱ#4jZ}v_�P�A��6/M;��9�٬�N��"B���_d[��:���� j��I��z��9z���5�[�:��z��YX������йW5k`R��x��B��j��
-@�ҔBL��(Η9 ?�Y�����e��h�S��3�W�fd��B�z�)
�Y*eZ�2�է -�2Mx`�k�ޚ�Oy
0�;$��&��E��$R`�	�HY��I~*Y�-�Eۋ�r�\�
X��76f��!Ob@"F���P$q��&%`�0�I$���8~�+x�0H�oɲ$$ ��W��f�,Z���	L��gIn�=� ��:�z' ���H���&�������?��#�eL� =�S���d���G3b|J���(N�f�`�j�4ؒ<���x&Fr�%y$!I�i��	t2�"����J~"	��BHj���%��`���Q΁��G��3S|&�B��!������ H�������e|��E���Y��h�O�+{�I�����\���v�T f1��	�*�
�G��P�6h=	!�<>���Y�8p��tb�
6���KD�dƮ��\n�z������ʝ�=�����K�k��y�k�E���7�6~��7O_<���#O���1a�;�v�"�C���2;�{��Ŝ���iL��\�)����h`�O����R��~	}�bzc�o� �uXL�*T�O���@��Ox�����+���K r�� 	��jz��l�L��A��f��T��8�����E�މ|4"���dwS�Td�|��Vw_v�ͤD��gk+��1��$W�A�"s�^~B�O��Q�?��'���)�ue˱�!��h�F/!Iye�<Ӂ�{��?<�����Bg:�T��*�B�6k�!��0c��p\lM5h�O�����ƭæ����[��nB����&��O� ���2��k��h���ِ����ۭ�;f�!�3�Rq&�f�V�Է���*��F���Z����冲���s�\a�dtCXx���\��_]ᑔ��Yu���������h�3��*��T��OL�e�"T��M���s�VjI�r����V�
/��ή���w�����ʄ[��w��S����d��K�=��8�6��d=�j������������j~iC�����1s�ֶ�T)����G*�,���=��:�.F?ׄ鷮G�n4&�g����L�)��棛%�9,�8.6�(:�`��`py�����������[�ۥq!	�Z��G��La W�1�@��$ ��<�A6R�cE��d��ّl�&���l�Σ���to^����LR�Lż ��Sӝ�8�k��]�q���y�����Vϋ1��듅\Bd
�l0��
 ��ު ~�l)@�ź����h����f7W�ו8�}�|?����j㇣��$=�Y�E��Xئ�u��ҝ�w��p�����y������xaLὲ/޸��A�֤��/, �
��'Ho�"b��QWiG<��yPm�3�V־��5Gb̷�C�K�^���8���W����ࢾt=��z�6-I��B��D8j��]dg�G�8jV�N��N�zՍM4[P�_��lǼ�����.J,�u�v2�NG�fg�٩nā��u��P�G�I�J���*Un��Ww�%gn
>����d��f�$�J>�X�����9~��<��ږ��$��*֖����V�/���a}D�@  �mVYB�1=,�f�������)��b�Ga����g2d�T �ϔ�$/�D9TG�"RI�09?��̟�ԉS���Ov�߼�uNV;dl�k�/I��Y��И˱��5&q��..�6��V��u�a�6�s]���Yd�,L��x���F.E���$��S�
b����/Sh���l�)��gHѮ���ʞ����R��:���� bj�Aũ�Uyf��tҘ��;�ͯߍ��t5\���\���,{o(�dW�$%y�E^�`�p?�(� �`��
����tN~3#/H�M�{�=���!N�P�.G��:4��m������������z���e�����m����-�6�b�������+*. I�ɟ��S��Z��X�`
��qG\,��F��m��ˏ��7z�z���RP����9|�l�A�ڐ��h�]LD�?�v�t�_��z��_=!^e�t~+nO�i\�[�uу�@?$3a%^���_	M@�M�&o%B�����aC��)�j�������������q��3��y�f��JQ��ݏd��ʹ��8bu�������������$F∉���n��]���9��ܳ&B�!c?������PUŔ�75OҌ{�r��3�A1�&<ժ>x��?7��W�׿y}�8��s������Vs�VB�l!���Y�-[%w����oN�}zuqu?�<U;����M ��	�!\"�(D��d>�O�3����s"y����H�h�n\�Xj4w^�}�ʭ�歩G�i�T6*�vI&�w�O��_}������`n��x��J�t+�2
YU�֛� w�$��%�1�i�؃6~��yQ����u
����Yq�;����J��~p�pxp`)�fM�έ�̋����B<z!�XVv�
��z���������h<��+f�����khP
-�T���'�W
�Qn��o������q�xo�XZ'p��h��z�������.w���WG'���m1Ρ����v�ڈہɉg\�>E����v������iV��ϟ�j�m%�r�u�4��"��=.�!*���07��2OaonX!9e�]F��t;��
�Q];��Y>�z��^����B����*MSF+�P�qⲴ�)(~�]�����F��eis�������d@꾛ᗫJww�G�W+��71Ɠ0��Ơ"F)؋�*�C'? ���ɩI����$Q�tB��`0�?�L눢Z���7/_��t��a��Eg젅
����-��mcٱN�F+���{�m�+�g�3vm��~B�H��/�I�[ ��B%9�`�|ve<L}i/���X=�Ӌ�#�Z�
�hG2�c�����l�(^��N4�?����vu�����77ӛ���h�(?\�n�ݗ��Fw\��O�a���P��:9=~��#��-�ZE�����ʘ V֪p{:���܌,�Ǔ���Ϳy����z2�<Y�]��N�I��^=�a�ItRC/�~��1����ɭॊͫ�J3�����Lĭl����� ���O�gnK��7)���^�m��Sԫ�T����_o���л|���h8�xg=��!С�t��==�������{����=�^{l՚��i�x�ww6"�b�ahL`���l?MӐ��	C�_1�E�u���:�m~0)�a��k̤�n�n�u��1���cjJL��Eԝ�g��0s���	�8�n�>�/o&W�т(�ҕV1�IPWt�<k�$c��x��oNA���f ��*�ϴ�������fc�q�q�a&��	��~�1�����Z���}�1�eS5c������������#�� ����C��^��7؈+j�����j��"E�"�%�+�$I$`x|�$���'�?���m�d ���
 �x�dF���}�G�-U�U�@�p����J �/���`"61$a�i��ə�W<�%܆��P|�EҜ�d��d*�,�/�[�d� Ui�O2��<��&�rC�$�o�)	��`Ɵ��<~�'�K���DI���n�(}��*�@~��N�� �*�0�L�;��W�^�/xt�$}%ѝ�#0nx��X"�Y��a=�9�B�B�po���u�W9B  "��ba�3}R.2�z�Q��ZKf7��o~�Jfnou� �������TH�]JH���[B��	�hd1�����7*�t������M����Ĥ���K2]F\V0|��
̟©�B$ ��
n;��F�N��������ݷ���Uar��(���v�اoi3�͔��d����.D$b�,����2$	f�E�閭�U,n�/,�Es�p��c,�����9Js��#W �앜�P�0�Ԃ�/B
;���C{I��x���ۄ�4)]��\a�gk[��ѯ� �lv��S�a�;���Zv���^��zy3���xu�00�U�����Mԣƙ�˱?.���-,k5�(_�\�}�A�o�o�0h�N?}3����#�AF�d&�b�!2 0!y� V�$�Q(��r���/�X l��؄'U~�|��"��&�@Zy��p�I�XN`��%چ�G�,E� gZ��O ��.*/�~�<���t�r�dF�$��,2��	#$%�l��ENl�S����72 ْ���@~��˟��'��%%�Sgo`

Yp`��$�H��: ��HV��`����^^^B�'����"#.�~8��
��D*Q4*}-9�0+#�FNYL�
4:N�CNC�������r�%_`�6�#�A� ~���s('G0v����JtH���r}����&&�H��c��������t�,wԪ����Ü����x҉"b�5�35���r8_vv:&�m7�ÆI��l��q��t�v*�p���4;��a>�6���_��,����ݱ'�����,�o�Z���֐�G��ʕ͢J j}9g�p )��j�?���>�EZ���Ն>�L�q@v�e�E<���@������D.�E�|J%$%f!�FV�j�Q8�Ĭw�z,3���h5����})tR�!�`�0�	�i�b�#:׷�>������h���g"AƄ��y��+`V=�@W8DrhC'0 hÏc<�'ORK �~�8�[H�~��|ˆ�����:�{�#�+cmX7��bgE;��&z���q��b애������^\�\��x���X��k/6��E%"�C�Ƌf�jƔ'��:R�x��8�5�{��\��b�5$�XWc��9L�T���˃��}w���3��ÝNcz��)AS_g>B��a���1";ʞ������~�����t���m�Ǐh���|�I�`����7!��N !�L�����!E[��
�w��_�u�=�+l���/6� #$i�)Lv�����n|��n�׷�E�j���������U(����Q�.��֟dcJ�C�QV�I��[tj�E���H5D�η1/�\|j���B̎]�V��I��m}9,��2�"c?&űR�Ck@�F��^���뽸[?ެ�N�#s��d{q/_�,nb,��3~
QD�7e�Y�c�x+�헜�a�լ;`�j�Nw=M��l�+v�{0�HI^��Ra��"GgHC�N���p�����z���r���Kwȕ��t�ݠP.��4��C�=Q�P
D�X~�Hvp
"����d̼X<�`�۶œ�,��]�ˣ�Ň���ݽNsѩ�Q������$,�ȥ*�II0�Q�hN��G�NOzFM�Z�`����B*B9�.ð&#ۏ$��8L(ʅ�.�P���Wx��3o/X�f�j�(��`��woZ{,w1�ol�ެhơǠ^N�`_?[*�]o���O�u�N�YO��-y�ir՗Lb#�!��M�<�0di��j"j�,x���	��V%�C��Vǻ{�y�և��뇽�]�
���J��ul���b�:��M+�D����pN�ѩ��𛋧/Ó1��r��3�]ߒg�l%��ĸ�c��[�cQ�(����g R3	`_0�������mvO_��،V�a�X�����fq�M��vk+��j�v���<n��Ք�Yi����v/Y����Bbq�Њ�O��_��#V5b�`_%�4?BT���0�W�6�[c[��D8z���w2vg���SY���}9*F�A�kМTcM{^{`�*�ה��̦]�����7����3+T��B����?��$��3
��!JJ*�-�C��.c �Tj�����i=���lhML�5>D�1ᑓ�t3sˑcX��<���M�������*���K5��5����{Aj��r㛥�Ԓ�`ȿ/��V�!d@$�^^�w��k��<�;����肊���hI���F!��Fv\��r��������ݸ���C��b�!9��Sh�L�Q~�0�0ٙW6��ߖX�"tglS��l�R��:=9?��Q�7̞�B��: ���f�r������{���������i��]�q9���<.�t��c���t� �()xh�i�h"�Ca��G  �)�m�]J�'iq���:�z�rs����u�7������r��#�Y�,V�<���ya|S�nl�n��x���ݧ��=�5����-b'�\("ܓWN�<!�|�L`��!K�j�F$�I������u qqb�a��w���YW�n��?��c��sO�k+Sf9�O����ܪϝ�c�W�Zs���DLt�[�N֜(�� �?CH2�'I�Y�v    IDATHЉ�����K3	9���5k�����ݝ�n�u�c� �c�&B�D6�Km㠷��{oU���N�����������F��}���M���6�$���`��|~��_����!8�$�Ò��Z����}��46�x^��v��j��^�7�XU�O���G���x���x�4����绫��{�C������u�ax���̕`�$������Oq��	�+&�IZdg6L���������c�!��m;kV�Y�ŗ�;�e�[i8�F 7@ȿDg� ��;ʌw.��x+Jͮ�G3���v������ed泪��w�u�g�����컬�5�����t��U�v}�S3�dj��`�6� ����`]qu��\��ifL��w��:����F������glo2�pԬ ����sX?�?��zv{��2Xp7�^h.k����:dM�mIg��<�b>�QP0�B8E0�7rq�xj�i�E��f���n�kX��nP��k��nY8�e�#XZ��Fs���t.�Ҥ���.�:yw��~Л�� s�{��?���ﺉ�c�JΣM3�>;���&K��ض��ˋ�A�"`f!$??��r���Rl`2��5{K�w�ן����&jO�7߿={q����t��xEKi�]uB�j��M��Tg�������ʓ��xr}n�d�Y���0���#!nc#?R�p_o�����ӱc�HR���0?�'�jL	��Y�G�%��N����f+4���	&t�b�u]R��֫��r\����J��o���{�e�M�w��A{_�T-�x��8��B<T_���E�\8�cZ x�9����ҙn��ܺE֤�-��d�����c�4 ��119��m+�R�M.�v��j9�>�/?_N������t�*�2X���֭�U��8W��#��7�6�0)�y�����M�����Մ�u�+�f��A�����ٕ#㔒�&1�����L��L>�"���^ݻ;ݳ��O�����X}�)f�ۛk"�u����ǔ��r�O���O�"� �<�2Pu�p)c�@g"TA��N���	R��&0���"q&|F���x�,r��p�x�$~�n���=�o�IO����'9<����"ʹb
�
���ƣ� x�tI��R:�ɢm��٨�E� +�����,i6���2BO�%-H�O��H���˂�'�o��a�I]D%*� ���<e7���eA���NQI^&�B�iP� �9��K������}����껾�������Z�s�S��~�;��V;����^��*i=������EI�Z�	 �N|��<�' Z4�QK�0�:s��_��_� zjȄ�����ϟ?�h�-�J��D���̔F��O�뚐��(fqܱ�)!� ��L�b�֘����lk"�+�.���2������8M�Ƀq���{�G����wߞ�8�7a_=��\{���r�8T.-
��Á�q/@���l
���i@�4�m+���ؚ��:8Hmda̓U��f���@c��;�-�h+�x�ܠK{�EJ��Ǝƺ�a��c"���W����ϐ��ka�b�0�)��PQ��ܔ�ITyܮM��e�P���W�7�]2�o�4�;G�Z����j�ؗΤrT܃��<�		�'U�/�!�`lۉ������ >�(��J��&J�@!b����OQ �����X `��$@,�Q�� F'���_S)�Q��W`�ж��ȡA�&�|����� a�� Qb	 �h��f�<r��K�d�O!�����K�4�e�#P�e�Y"-ZQ � ̩P��A�GB���/��n�� g�rI!`t�����	&Btf0�O�����
I$��4ʊ���%E mO*V�@Z��O�g !���{��WF�
	�h?L*�WF�1�V�hH ��E= Q�%k�@���O�#0 �o�*�$����������ģ
iA���O�+�R�\��(��
�q ��H�����'��x�qT�>Fx��(K���B�I����*8�ʤ�r����I��bя ���nA^FI���W:�f���M?$�F5�b����*-���1%`�����n��k��W�,�G;������smע�m�(!�l��a�8a��-�FLΎ������}"o�t���k�-�8�%�~&�I��R��VхT�������P%� �o��O��!�%�q ~.��;�Rq["�B	�BRȅ(����'o���j/J��M�kb�i�M߰6��%��,���|uh��$������KX4�O7�÷�.k��M�
���J]�����{��D���#��`�׎ )�4!DHr �[��r! �Q�RK($1K�t��Y<B<Tq||dsy,�0R�*"c����6?�Z�f���%��n��_=������䚬i쩯��	������M�YݢІW:=8��1��㕱SjSw�H�h����횲��\�����Z��$�'F�����N�xg���W4{�{�ޯ�6���Y��z��y���Ƴ�w���_B�m9�a�p`�`�0��.�W_�cz|�����Bp�WƬ����V`���3*�fa����'�@�f�Q� P�m�wY���t3�=��&��s��3��}�4��%iY���Hp��l����m]���`���k���?*�A,Í�#\qP�V�7��h�2���Նv�9�;�T_��c�����f�������[��Y���᫧�ݼa�_v�
ֆ�M��x�5Z�v�9#m�eY��\AlH�n[R�kQ!��q��4[�_�}�����~���B�&R�,�jbQwk�_�KF�C/�M�����S4[V��Z�B����"��EH�5$�c/�r�N�x8Tɂ@�V�=�D��5�x��e��'Ê����z(6̄�o�����iy�eޕ�d�3��o��^5�3&�F��g�;a�=�ۓ__s�i�Uw]UJ]a��q���_�/�'��DXJQ
�(�/JR �8�
v=S�JǠ��ͩX��D�q���>���q�([��\�����R��bb�t>]ݯ�z5��ޱS�q�} �CUR���W`\`�*�T��J|脩e�W�qQYE�e�9�I<�<P��mg����ɗ������:
f.�k��(6@�(w�@�v�?/�i#oӟ�^s��ש�'sF�a�\6]�rXt��F�RdB8��+W*���"#'U\�6?H���9��z�����Ú*oJq(妏a�	��E�]�X0goW�n'z�؟_�W��j�n��N3V�@|�ʘ������Dd^&[JB�
�iH`b�;�,�f&N�=��^#cNp���������<v��-AN�x���č�ٙ=m{cZ���c6�ܩ���on���ט���y�7p�R���$\���I���'{ќ.+B�MN
�	��ɕH�ZMV�R��y��۵KL��+��� RS�v�}�⏉��{�?/n��ֽ�f����z��"4D���p!��H?Ae��<�&wu�+P:�
������dV���{r�x�0��:�oi��z6��SFMV>��I�e�l߭o��ΏO:�7o�2͘mwGH���'ͻX �������-�X�+:�}�H�T_e�@d�sB\���ޞ�<��v?(E���X^UN��k6��0��%�ov�q��q5��t����:(L{�충X����j(1�
&���W��6�e��q� HT��a6�a�H��u�X$���e�np4<�g7��Y���2Ǝ��۬�Z�l���ʽ����z����`T~�±4R�}e���!�]<��$��j��t��`�쫐� yۤg��R�P5���o�yuv����N\��A�؄�Q����R]�=>}��^?f��4A��E��������rA�*Z%�� 4 ���_�.�Ҥ��� ����u��Ӟ>�%y|^޴������mW(�:�D���ZS�����G���(��WZ�o����������=����r�Y�pag�n��V�yD���#�`G�9���>�b�$�r2�*���n�t^���C���߄������1J5�^.B�כ�G��j����a>%�\�F���7����Z����	�g!6���Cނ<r�rξ��u����~���ʘ-2�
aǆf1�%ȳ������K�}�����y}�a�'.s[�Mo��c�,V7���8�ո��&1cDK��������ϳ�p�U�K��h9�/�g{��l<����ő�P����U#|6B����|�ɵ�FN��&E&9�^���_5�}�҂b�$+gL��?�Ī�}jy��\�W��������o�����dnC�h��G�1
يJVC$�,��E?�+�$��'�
�*��N�5^tR$�r-A�L-6�J*�Y�vDn1A�;��ץ�{
�PgݎZtu����I�p�RN �s"n����u^�y�Mo�Qa'?k�����?�w��ʁS�C�=b�4��#9���R6���r�oPd�� ��_ B�^=��Y;%?��o.��㾢����~��q�a�1)�bR�+{�d�=�p��2ɛM�<W�����KZU�%qU����#��6L��r��b�L<PE���d�z��Ip2QH��]���b�Qij��RѶ���dOo�9��Tv*����FK� э��|{���+���}����;~�����7l>7\�3������.w1�J<v<�hӐ�"���0�Y�p�Cjj?0��D��'
I��h
5��}��d�]�����s�"�-���h�q�/ۄ�w�_[X�9-�ȁ��i�����f�|ԇz����ZF��r'�m�tC"fj�)�zI���}O?3���g���������8f���ӱ�6,�n�=�r�N���I�@�*�:���k\��K�2��f��jV_eu:ޛ��:��l�\��v�����*:e I��#�x+�K&�6��q2Q
����	�r`��0 �� �܅�R��L�@N.����
�ؤ� �������N��4���H��?=[bf�/��frP(0�P����6;���U,g����	�W�f^p&��.�9Q Eqp($�p�l���A �'��ȡ*�x$���*r�&H��K� ��H"����l'y��Byz���_�,����S�&o�������#�������%�T��a'7�U�	���~������߽{�b���{�iB ���D������ �M���x �W����o��oB��2V��I�bgy��A˧
�4'��D��x	�bX�t �����#�^r_y�Q�Č���a�x���i�C'�$J�B'.�(�rON~�ۿ}��p��<GC�5�x��\&l��8WW�D���8|�h,z��Ď'2�h�NLPLŨ8:������z!*�c�s�?#�?�0$�̩��I���-Qbm3ё�|B�5v���H�<��Qݡ������(���)�ć�+� A�4c����Ӕ��Y�U����� }�cT9�������I{o�ܰ3g�vRm�����,���/�v�O\o5[>��٬,,�E�V;�@�E&HB#�$���0Z����U�G1
�|�er ��r�0����� <Ҧ|
�(���"�r
�؄���$[�B���Wa��	�R����?��	[Ƃ�2a��B�*�/�P�h�I"k ~&¤G���a�/����O�~�d�k>	#*���B�b��(CB.�Q~
��"*�~r� 8�C�Y'XfM'�]lz`� 9����oRE�@K]҃��8s�6�����g^�#��6}����+xR�ZѴ#��E.4�� �Q�����i��� 0VZY��T3U��D�D�i?���`�AK/�6��~n��0�Z8�_Z!�D)�I9�	K!��SH�
m�d�3~� _����V.!�~���$����%������a���"˂KB &�BF�/l~
�2�'	.<ِM*CݺĈ����3b7��=�\�`����.��O6��J����J�)3,s�Ɣ���ۮ?��[����<�1���τ���X�d\d2�Ñ���C�6tS��	��J8& ��Y�DE������+9nH��D�gf�KT������ᗅ�� p�(nKI�J��JQMqz��g��.���l^��e-Є����1+���X�,l���*I�{.2k���-�'CϜ�HS_��x�ǝl[q8&�|�<�G��~",�,�G�PQ��r
%*���%$�$6�BHd�uJ�-���ƞ�9zq��s;�q�
�(��g���z\s��`3]>��6O�TVS�nF������~y�*.EH�f�n���؇�?*6�sQ�0H9�W�x����!b�3���(-D�7�k�s�Z]�9>h�[�)��"�z�CbL(��a�Q�(;���FC�~�ؚ�M��z��tc��"�(��L~&{(��Γ`)�ELT��2��T��8�ˤ�\��x�r����X,���"ip>VΌ�-+�[%^<�������������d����W9�uq�J0EE.�����g H�|��T�]$��wV[�3m��T��/�ن�V�n�ݷ��ܼfW�4������e�)�r��hM6�`�yu������߮�w�	󝁚���P��d���O�r�=T�G8�џ��.��l�!E��e��q2��h��˳c�L-��:���DU��žu�!��Č�ñ�!&��������~|�\N�'W�1�pR��s/ϏKhӧ$�CP��$2��"��{��Ƀ�5��|3̈uU{���9�j�������˷/��-;�]Z�U�5��y	ۉ���.�ձ{��6K��~w��Tک����ܱ2_J������do��`Qʆo�\R�
���T���FR��iF����W�܉�۞b�kX��s�|�!<*����8o��o*������Ç��(F�x+G|�L��7�o�2r�zL
�o6��b��SH���K��P̬8#��KN�T�^��Ql��Ǉ���`�Ӛ��[����vW
0J����bk�b9�L���֏lh���C}UnIU�m7�Hj�K�r�a�Bғ�	�%�G3x��z	j�
���R��Xsrr���Y�%�"^��5�� �F5cS�q[j��7w�w�0���x7�</��K{*�jBGyfؚ�$�
"��uAdO�x��dd��!t۶���u�����	�ҥi�������;ϟ�X���uF��+fgL�����Ca�8G9C�7��x��s��U��by�hz�pg��PN��Q*lAOָ��Z�a�I
�d� ^`��S@_�d�����D�Ξ7>��A[@�N�<�oƩB�]�k��]y���ӛO���r��z�|,Wg�5S[��%S�ڔ���$q��o]'b��Ƴ���D?H~;Ϝ�(�������tʶ�����!�f=��Ǝ&�*ǘT��}�z�N�*��	�:#�����z�=��k̅l��ձ�#��R$��Ny�$~�jAT�T�JAjQ��(?�ʣ]b��h ������;񠦵3��-��(a��� ��B﹄�ôI����rrq5�}r�֫�a|��J�\sj��$J���y��L�Η����ʑ܎
(�A�d�]� ��#"�[�WX�%w[����N$��zqb���#l`6N�7��k����TY�����і:�[/_�:����OO�������|�il�4y�R��h��g¾*v?Q^�ND�S�,�&�H�a�ܬ�~p���{�o���F�t������!��+�����Y���n��pp������Ҧ�fq����~ޅ��c�ň4(dI��03)�;nk��Dy��U�OS]�D!>K��6���Tr5{4�m|��Ru�T��������%�Q����)Xg�7];DUi�읟�}�j�wO���b�P(l��*j��qE�pOJ�S"T��?Qx^4ZA����	�2|z��������;Θ�v߼>�i��{{ cU���&���g>�ٸuL�1�������ut51���e� >��%L$�%7�$X_�    IDATV�~6�$����f����3�e��iUA|��KZ��Ec������ҝ�KMǏO�O�k�v}g�i�F�������n4Y�,��ff��v���tO��^}��֥��pW�Ճ��z���1C��q:"8��5yG3���MZ�h2�A�(9�<W`��nAQج)������ӚqT#f7!���⽹~;�o�����?�����^=L�v��'1���v��"��ZrD�%�ވ��9�����a>H�%�{���x��H�8�y��9��:UB<���\ݟ�����=�-#[E����8}�-�����r$}Y�=9�v���;��c�7}��>�U�wڕ8�Y��Xg��o"�6x��N:��RK$�(�7bc'7��b&0����3������u��j�݂g�t���ӽ�c�X�v�7j6X�,��x��l�7B[�j�^�\�7�=+`���<y���/���D�媋�s�����o�gR<0��� /��>ǣ�*���}f�N��C�{��b�7�z��������ʊ~,��v�v�7;�e\�^��Ƣu�=��g)��ӳo��	zw=�g,Vӧ~�������.��]xHZh�h�����Cq̖�'�_Bc��@fdW�^^\����V��g�i�p]�������{�c6A����u��^�.����}1z�|������i�8-%i�AKe3���YΉ&ڣ��̢�1G�f�#-~�ht ��/_�����4��b@��4�۾����o{ak�0������JyzC1�]L�����tCs��%;
��b���ix���	��p�Ph�`�F�K��c�R�MW"�AO.�{e@K� �?�`6�� -Tp���#���m�[<	3�[�&�-dz�./~��$j���_`f��� Ϩ��f�,,$Y5�dB$�%�<��NT�r[���0�ޖ �9�-$���S*�Hl���D�B��<�ܵQ�	<¡��7�@�Uᙣ@��S.Z`�|e�3�7�"|�� �|*���a]��m��"
�'��#!0r���i�MھƎ��o�Z����hR�Re��q�Sڎ���9 ��TX7�3���Y0���A���կ4�P���gh$wIL�(RTs�I�*!`J>F]𦡜ƷRꙺO�>]GDA�[e�/J� ,Ȓ�$YR�@5롑F������`�E2����w���8�/a���p�<�S��H��
�k��/_��~}��nǛ{(�<�ȏE['�9�b�m��Z�-�bm�8OS�U��M2�b���B��ъ�}Ԯ��(5hS��ɜ�R#g�%�"�g�V<�=�l����ȯ��0�Q�qJF�qsa60�ID�9Z��h�߰0y���ԕ�*�� U0�.LjšT���4��z����(M�nFd��9k���*`��kk�<=s~w���33]y^OJ�AF�sFy�����PYh �jJ�E� �@�_�M_��_,J0|��83��D>3ʄ�ʟ[2\ Rq<pfȖ���33�
��p.e/���6����3!�f­Z�S��t�*��I` � 4�l8B�IF�g�B.J��<OX�@:� ���Hv�#f��1!	d*PZ	��M�I�$F���_�'�,;�'��&�f_*`�m������<��3TP����6HJ��f���SrDB���-U��b-�J!_�
�-�}�m���?���
Zk� ,j�J�~4d)�h�K%9��?��
��)@~��;���:0e=Y����v6RDp&	'I�'��'��J*Y��"I�C�'����/�B��Ṽ��s@%! `<`�����)
g2�7����r� ]2J���3����$8��ޮ��,5kcݰ8�Ү�ڶ|��W�
1 ��ڌ�����F�L��h���0�R�f��n����8,Q�����2����_l����]$%=(GdV��R�'?`d'�B�ĺ�\�<x^�M��/%/	���@8��\�J-z$�і<� $�0��	^��0ы�`�b6�X�%�r�.���Bԫ^�`untv�����Գ���!�6y4��[u�3[�]�f�gy��?���C�o��X��-,��	�N◴!8��ɒ��ۂ(`�TlrUVH�Q�Jl��j,IT`��bb��8g�����ٷ�����Pjn��)l�]��af�-m���d9d�X����?�q��m�C� !����<?uԸnP��~&��<b��@g��E������~���]��=-�
���f�*;�o<u�a�R������Ys��6�|����Ml����2,�X4�i�X���S�J}����n�H�X�<BC
2R$p,{�-��c,�}��K�˴ůt�C�c�*�����=?<�)W�$�4�.��6	�*c��?�O����|�{z���o'�����\�E��L�
L�;sJ�f��=S,T��#J8�B&b��sIL�ڙ�2dPYF��l-O����`����ۢ�����ZN�k�2#$���Ba�/&O���|]m�;/��o�~�Y��Pm#�J����U�!QX�B�4lD<Vg�(Dn��m!K*I�_`4���8���`;=?b�Y;��4�Eڐ�zdT�Z4�Qy��vf�Z%^���6}�M���������f�`��q����K��g�W�"w4�m�rIf
G!0QM��Q�c�#��Hig	�ª���4z��ǥ�~oY�e��eB��K��MQ\��48�`��+���wP;�n��ϵ�˶3f�+3{�r��A\�Cy Ih@L�Yt�x���)�)��WT�X)F�0(.sZ��^��쟿>ej�֫	"��׺d��vz' S�G.�������m�
 ��d�!-����K6���!��a�Hr��L�b��]�L���'�rN��[9iQ�D_K���h8m{��@~U�=�|>v�]+�uo[5�=+ihC3Si�o�[�gcZţ�Ɯ��]u���Q}�"�v�!�Z�[� ;�ԅl+u�p8)0K��` 'd���p< |I��!�Ͳ�G�{�v�6��T�Ce�Y"R�\���`WI;>sTm�����=�l��Ͳ��Kd��B��4Zo�)���"pD�
�����@N�Ia���gq..��th	o'!I���&����n�R��}��n7#�2���i�����t��j�I����{�G��z߳�n"�.jJ�&?��)��zWȳ(e�/zx�E1�� T��G�V�[H�J��[�zq~�@X4�gw�Z�Q{�����- C':�����Z���z�Ao��?��{�j���G�C�6:!��jp� /�bp��v�_��2�e%0�L�w�=�3�%IQ��(��<�o�c����¼��K<��Ͱ���GG���ż=�M�l:l��I�#g '��G��-���}y�>�.�6��C���Qp��P���`�&9�
Jb+v�>D�d�w[)? ���-�}�1LY��N����wvQ�p?ki�̶6q0�ӚF���k�/�Ç�q��n0�q��Rd�ʆ��ZU�d��g�!u�� �/�˚�/D�o�1�SL��{R�\ȓ�@�jo��!���
��1F���^8�2�\�}y�����#�b�ذ@� �U#K㤸�s�[Oq�_�}T���G���]�y=d�*�[J�`L�dd@�'���XWxr�G,��A�ׁ
W$��R�!܅�T^��vlH�Jǩ���}"`¢8�;�b�v9��|y۟�6mg�bKKmc��c 1f(�X��PV,�F��mt��xlf��Z.u@&цN	���BT)&7�2��hT��HX���m�F�2S��W�vS%m,�m��"ldo����ҹ�W��/o_��\��c#����J�m�;h��E���-���|&��bv4OT�Tb��(v=����l�__}~�4�5������ᛓ�=�^�S�;:���,���-#޼n�C�Es���7N��k�����4lfsCo?�0db%!f�)��!�*�ryfd%W:/��m�g�m�l�h�%\����� jba�ѷ��ho��K��=iMMwi;��]�B�!�j���x�O�ce[���n_�_�j*D7^]Mg���l�m֙}�I�ǈ=fA���8���ׯ�<6/f1|�%ہA��S�a|����O�O��=�+��`��[$�[�����ciX��p����z7����Ȗ U�*j*��~R
���)C#�"�	Y,�DZ��ڐI�:���l-Ftj�Pτ�Xm�M�a+��q�5���?�J��ԹX͸x6n��ƺ�ۊ�M��(�v�����U��S�vOZ���|h-���?ޗ?\n���Dw媁�YC���f�5���f��^���w��y�v�{bOF�A���������I���gr|���߼�v*����������Sm��EM��@��^���.�<��Nw���;ci���`Us0�9�ޘ�-�Ǵ������A����rL?���T�^b�n�m���C�����;�֒f�;���QvZģ:9njD�i�E��Vf3���iܬt0��9�=?;8��v'WL6�^���{8�霞쭚��cd�b�{�HB9��'<b}ɉpC)Z�RA�r�=0������l<��{��9������nʧ���YE�e�E���u����a�n�]c;{��=�k�+�Σ���]���g��:*�	0�Q��#����f��Ȃ흜��W/�\T������DD�d��d�&Pi���'��{OF��W�=��%D�����	;�UT=��Y���������`-ۍ�����C-�>G�ƥN�3JV�Vb�pN��c/b�b#D��t�	�:Rj_8���<Bxr`�
�X!]x@�'��S��B`��a�\l���/ȓ6�	�?�	�5ȏ��LHz���I�B�$��_&dKU#�,�pJ�D��F~�q�V,������ܖ�=�����Eb�_SI+1[���/\�	����<	��y��8'*!T�%�);����4�'�$�(0��L"\Hf�|QEM�IEʣM���(HB��*#��ϒX��$����.0!�ר�J?~~~��?��*���>[d��1u�$�;�I�\^^��4Ē���������ԹJ=l�����7�N�o�Sr�B",�� P#K��ݻw�~��\��'�DX����4����I��prx
'�A��!�(?�'.�r�±�U\>#���-3���(�ʌ�����~��{q�7Y��=��s2�u��뜾���v��б���R(2.��շ(���i1�2�1��LZ� �b��%-�ƴ8d�PJ�!�Q1�3AWX�
Ǌg�mv���0��'3wq+;�d�Q��v����Cg�39�XB�FX��sb`�K��Р�+�"v�MıxC'2-v3h��9�z���{=�#���ը���:��?+ϓV�{={]�N��֯cb.���V��ܴ%T�$H���\��3(/�cK
�R�	 ��L˓!R� NH~.�J�����|��T3<��eB`�B���O�~�S`��\�����_8QO퍟K���Ey��7K�A%V��V�e�0q&p�-$)��RI��Q�x䒘3S�I����^ '#QB�4 �AT�Q@Q�o�O$�
���S�XR�?p0@�_�(�(��'U��$�2n��(��U5Γ%ŀ/�/#�Rk��h���~)S��}����ÐK��}�
�X�_j��:��C��g��z G��
5H��'�W1!/��Z�r �-9͎ń!�@vTqj|�u�(*;�Zr�~�TdN^~BNe"!l�cʊ�_: X!��'IR�	���' Q`�PaP�B<>�"C lJď~4���I.V�}�� '��b��+#Y�<�]��S�^�m��^y�n�\��5�g�)̃Lju��'/1�YVk�8��jԬm�d�	��͜���\�I�<�G�06��/i��᠁'��&�ۯX~�J�I�!����D���"���RK��I+�Ox8e)6~_�~&g@��	�$r@.��g�/ Y���J��H )~��;���;g7mӈ%�j���[K�aSylgv�QӴ��İ�5��ˀayq��R9:��nz���E���Yg��� Ya_+4C��UI9'J	�@~E@�"dY��p����q^�A�e��ч��Xz0�o�7�|w~������qa (������}7�(��n���ރ�闧���¦�&����P��sj��������j���/����F@���F��Q�iً��i{+`���X�X�aG�$L���rlc�&�葃j���ޭ�7u���[ސ��X�sZ#����tU�Y�q������{���.��h#4@nG�L�B���vK9�n�M���Q�	����O�绻��/�:��[�,Pi}��q�!>�w��m�5��5�GO���}����T�9���òh��b䢞-MF.�`�EK�Rz�a?)�=��Ж�F4s*M�{���0�,�2Z!��ˆC�ǻ�ɉU��P��P�ڎ�h���[O��e�ĵ����ڙ��f0�Wߵc%&�����d̐���{YY'�1|��`��-����י�5Ȓ7��N�.-v��x5��C������<+VrT%]�I,G���+br1��>=~�b��[6���ȥ�K��3;;��$�I@U|�
���@��O�!6�#��2�<$��ѭS��S�U7X,=�s=�0�Y��ݨ�p��9릭?�r�U��9���A:�zV�]��0���I�Ӛ�mƳ�rs�-*6�D��<��R��N?1_�~�<pJ$�7+�7k$�)��!�q�m�/ND�Q���6!�PGq_��U?�3c�8��-
����4������jq�>X�3!;�ayrDCQ�פS8J�4�P�N	��yѵ��q� �+a�����hS����.��pv{�?>9pj`Ӎm�Ȇڈ1��]D<�Z��|v����%�}���Y��z7U����ΦO�(�j�������@�P�U�PA�W�� �� ~EDr���!$�f}�ۈ��폡,�𙈅���֒�9�3u����ps���~�<7Y��tA*�9�G����b��δ&�cr�3�c���Q����J��#ל���e qӏ�hs=��[����u��[�+��t�a���"��B�4��۳O��E���^��Sk�Y+��.dX_#Sm�m�E\��C_�O�)T)B�������$Z������U�����w�GG��|H�ċun�|Vd�	�̇n&��=	9x��=��'�b�s�~��8��$ֈW��o���qZ4����,@��5��q���T�!�~e�H�"��F�U[wh��zK�M���-;��AI�<x��z��[�<���ۺ`�뾾R{�}pz�|O��݆�~��Ov�)�u|E댞�}���Ԃr�M�Z���~��$ �K�K8����,6��޾A�gU�FG�t#��B�W =N�a�!�]T?�O.>�>�f�읔k;ݓ���ܜ�=Ζc�s��F�h�ȗ�����X� �Y&\Ҍ����PH�FiUXq֊����`h���"��9]�[�k�u�B��Zg�C���#M�2��PNvݲ�n���`�b����E;�I]���/�{�.I��C_��V��n��A�L+��0�B��/.���j�xmx��0�?˅�ltp�1>�*�
�޳��:x����7�Ow��My��h�֖g�Q��!/i�I��������6��!���i��d*��x�UI��{�Tע�x�ܮ��0Y�S�E�yj��l���`���"��BBjn�*7�@�P�{.jݗ����.�|x�C����k�fҘ�/
���v���CP�\�g�}c(ɍ7i��������{�����^�����~9Q�uc��9_y�QY����n�s���?}���b4u�ޖKa�f8"����;�hzC'���	-*�w�'Q�-�<t`�t0��HX(���%�{��������_X�+�Cu����K�;z���Q���]�2���><���ળ���V���rv`�m�5���	v��2E@��5�mBP���;!�"�C�"���1�ޟ�
O�No�\٫_FQ6�x��0����I謩�ءU)�&����6B3���qt9@e�Y�3��d�D�	_    IDAT8JZ�<y���}"�I��"2��Eqb6ĉ��$�9
�P�|x�z�}x���u��rࢭj��zѮz������r�*�#�̂n���o�-wv^4ڟ�<1�Zwj��r�ѻ�&��RGk�:Ff�5Ĕ���<Ock�˧��ѧ(�֡��e1C!Ď=5m�i�jtw��|9ό���:�uIH�ۺ=CK�hQAh�]�f�X����y�c)�����}z5���6�=�`
���N2'���G3h�Q"'{5mr����li�s��éa�{�нA�|Kl�i?�l���w�ݱ���_�if %@ڿ4�]nD�(�9��յF�G���ێ�9z�����z�Ju�^t�b�7/d;E%�U�����	 �E]�w�}�&F�S6�RY�6��T//>�\_ϧ�I���g'���k��Yl�29�x�&VQAq�ۓ[|��D��/֍�:
�&5�F�J��E_�c9��i<�-�nI"i4�Ta��=�Tll���"�e ���ve��\�[5י��q��[n?��H�I1��B@����r����ai�ns��ݱ�^v��Mm���'�9,�p�ڗ̠�t����Ρ��A'��<?	�ʹ����$�bE%��~ 0��o��! xd��~J�T����$1��d��E�T����N ���\�ITۢ	�X898�H��Y������8i�D`��4�3S_L�,w�L�`�����UP�s��`�L����[�x$��\�� � ��X ��Z���*
�	�����,c)�I��!Of����NQB8h�UR.C2G��Tv�h��F	50(�k���x{|��N��@���?��?� 6H��r�2TzI�AisYT�z��/x-T�������%��?��O��-=L�"r�R �"��i�S�RjN2�^����	Ƚ��D
���s /..���?[��+<�/�HN�
)$����p�@�8��̒��a��p<Ŧw!�����w�w�Տ=�lS
H��E�^u	Ţ#�y�$�X��&�=�(�wwG�Y-����dn� FG��^�Z �n�Q!j�ؐ�"y`
�AD�Q����wB��&iv�nj,�7�@�ۭf�*�]��$��)@�Z�n�ѯ+b_��b�52`�L3�=�ѐ(5v�0��G־Q�P�XÚ��� 'X�Л�z�#X�
~}6�j}���׿5���W�^�e���o��Z-�t����	uO��P.�C�+/Jг~S"3��f3��%���0Ŧ��%ْ���7%p&�-` B[Ґ��'%|��� $�X����_l��j,$'P��� �Rq���'���Te�ʕ`!6�&��X�6Ĉ���8�fF~&B�E�_G����p�e,�}�g�@��9x����%��6�.2
L���&���G���� N'$��|&���gh �t����KB�Qy��x��9�����Xd#�S�|��J.<��)#8��P4���:�Y���8�"V4�(�Q�p�o)X@�@�ɓ`I x��+��\�iZ�
c#�2&�d!k8yd
��ϟaPd�`�R��YSR�gf��Jn+��$��#��!/�3`aD�C�!l2<C|Q�l�~�B,��%ϊ�~����bKL��#@V�'� ���$���E�gO 8#J����`&?Bb���r������HS`�Mx����SB�$���3���tj��H��ɺ��@���,0��+���B� ����b�`	���Fv8/m�����
TM���i��{3�vѿ���9�7Z��nQ��j�z�ٶ�=��;S9�8�V�<N�n_��h��ӆځ�@�����t7�SG��B�"I0zА�ǟ4g�3���p�j�`|3y���ว��>#?ו���r+�ʻ�{o��mV�鄡ڌ�}�zc&%�"�l���!��������w��/63�Z{<���$Hbd�B�E|2�?f)���6��%ޞ��'�������0���7ak�zޔ�����H&.��OO��Ǉ�^�h�}�����bǙ�p�<���t�=Q�ܳ��j��ø�����d��
V�"�B��|������-K���¥:a?��y�Y�r<A]�����wR���Tt��8�fo�co~?XUw^2�,�1��Y�Y�~"I�(�O�@[�&������%<lg�\t,�Q4
�K�a-�Iwe��0���OG�fS���l��my�5�fjrlP�z�r�Ĉl �W��CA���s�2^VM<����4��4G��8�"<��g:�<
����h����:�ףּ������pi[��e�^l��!���ĕ�L�N�nb����?�?]�~���A����ՃXz��H�U��:;=#�?���᫧�1|�ƣ��[	TpG�,,Uk�ǧqӯ��Dm�����a�xt�pS�*!��8�Y��lY2T�~k����V�Uv�V�іifc�|Q�h���l��))W)�x�p_�`26�Y����62j���q&�VrÂ*�[XZ�346�$����l>�29�y{O��"����B��.SyIE9$�S��/�ԦI�a�/H��[�i�@�t�V��K0�\z��a2��=�욈(1T�U�$W�(s�i�`�O/Ÿ�*P{w�ќ�u�����ypS�X�c繴 ��Z�C-R ��m�$���)���F��,D�z�,������X׌�K<e�-&�������z�|?gu���1�q��a& ������6��B� y�L�y��b�*!��$̈pkCq��zT�i����w�'������d1��״�#� �g��E�i!��OϬXݺ�:,�2�7�kM��)�9)#�_Tz|�2�g����$��r�Пs���`���E�pZ�]�����Q7�X��l:./ޔ�n�|������=�U�iE0�h/xe���O1YF��U�j��A[�<���B�X�p_5� ��P9��>d�]����x�	}�XMw���D��9�`�U|��߱�f�E�
�����m�iY�q���[�bOa�xɑ�ǳ��9~��L��OE��'	�Q���g�4w�{''�{-{���yD�RQjا�v��bdc��h�՞kO�8l��u�;{��kN����V�&�����'�E���ɡVA8�$ k(Q"�Y�Dl9�igm-� �8�?���o^���Ȼ� �z���n�F����ņ�b��K�,λW�ޱ�,�U+⺫� �� ���7&/�IQA*O:,�V���Ϻ�&���ҕʋ���e�N��>�<AgfU�Y� � �"�V��n��ڌY�Zۗ�q��A�mmkI��H�A�,���̬���}<~@J���w�;b����ᝑ��v+U�)��B�; �\f/�2)�����O�of7���;Vδ�M������ЀB,�OZM�:m�\�D�qB$T(�r�΋E9ߓ��5{(%�曪w�ڇ��-�n.��l���qc�_��E׺i�]bUY ��Q�ڿ����9=���]\Z*d��j@���\4S�o8�&#��JY 8�}-��q���E����6�Z����8w�8�4+���eJ(E�mjv�]Z�g�<����/���I=G�@�ؑ;٢S�Ώ�(��J����I��D�@_\`Wj�Ǫ?Q�n��� ��#������ʎ����X��;*��X�k�d�h[�Z}������9�:����{�0�f������\U+O�zg�E'a���ˤG�ׄ�<��	�!!~X;w��n�=`���.6Pi%�|kپn��2�qz�Q'B^�|����}��u��	-� �ν��JD%�� C!��*��)'z��#-R 0��~V�k�i��ښ�~������w���s�^�,��%(��[�Mfo�EՆ�G{ww�/Δ�������L�>�
aH�1L�c{P��nx����Z���͢xCW�:�]]��q��56�3�1����'�-�O��0x!^���#�*�R�y]r����C���������?��XM�,��_�;l�#Y#�~�/\��C����oŢYg�a)�h��ӷ�$,�P�:����ݫ�N���-O
W���|��a�*]3�����B�W(���K��]y[m�ܫN��'��׋�/��^�bZ�8�u����2ڠR�tؤ�`�0BU�gw~v�	��K��s�*�����[�[5��@oQ��5�����L�v����2h7s�\;��<?�]�Μ����̶��2 ��T�U:�#D�������snV=�  X�I�����`�	�$_vE�Ǫ0�����'���C���v����@�Awb���y�I���f0���=8����_"��<�:y;=�S}�H�� Q�}њ5J�b�SaV��	���R���I 	�'��#-$~
��"$�p9n0	�[����sЊ��pSF���`x�J^b��[`�`8~�$�F��nB`+*� x�j	#(mPY$+��z(0��	�iU�`�G`@��~�8���09a�T��<���\�pA�� ��
G�0~I ���@��1<�P��|!I �!�O?�#۵���g�}�Z����:���(�M�5Du����OPR�!����'��|��I&��n����;�b����3��ZjD<���C�������X�����^b'@Yi$V��ƀdf�`�-�(�G�ze�Rޚ�H���F�_�0� ! Y�	�\��$���P?An��/c(`��*{��kK����c0����ɧ�n׋KOW��na��1�Յr{^���]��u)�Tpն�IR��n��XӉv����r��m�Q�y��lu~��:�[j'oI\cb�T��b�)�kk�C�����+m��i���V�z�E����.i����򶣆�1*/ �ìs���K����ڂ��m��ٹ��_��W���M����/����'?؀2��P�}p�c�t|�}��3����vzН.�ѲִQX��_J_��(ty�L
���9�2�{�Ҧ�����	I������c�%��	=#З
���n�)?C$�P�M�x4�MlX�$<5�G� ��B�2����b��R�#,��70�� !�|�Q ��@����d�3+�E���Ȃ�W��.ZL5��@�7H�!�$C�� Z4��Q��LrT��H0��%fG���XS�*�H���1�R�Wm��u���}���~8Mo�׫�'l��,�A°�7뎱�$F��ȑ1D�_|�6o<S���_,HI�&ӡ�E[
"��������T�E$G�`��) ��)!X�\`D�I,��(h�\,<���FU
׮�F��B|��;h�hq%	���o������JrN^�	�<�u�j����p0�_s�� $�(3�8f��P��ѭ�i��o������/ !]:֩����kq�PKJrA���N*�m��� �d��<P姒/!�H�b��#ar����#�(l��,����C$`�s2���d?��S�*e~[�'6?��ݑ�s<��^�8����pg{��=,��^�v�E['_�زJf����^SW��;�������{vs�"_F��c���,M	���
Fǃ�kk���b����`�_X�m�*U���a�QM^�&Ǉ����MU
�*���eg��m��r��e�ڛ��S����;�81^]��Eˍ0��,��� p)e��NȢ (���pNidQfLa�"�q+���i�A����C�d�25���~�zg�����!&����CTQv����0�P]�`���c�{��&FV���+�Z0�;�;��
я�P�;R�"y? �o����O`4N�h�X=���wG�r׏e�v�n=R,�a��Y��/ez�s&gvj��|�u�Y�ެ��~^e�#3"�Q���D���5�n�*1���Ypqxg��n�\�$�ߚh���DIUm3���Z�{�z:�T�7G};�KN�8�]���ʫ���*�<ӂ����[0��$g���K�G׋��=m�x�mc���>94<o������"G_�<��B��,-���.-�,���ѭ�g3Ng �6����^�qt-L��m~�ry����?�ì�z�s]�2�-�A��mV�C�IEQs~" 0�8?�$02T@	�=>r��q��x�v����?�Wo����7_~�_�`�]��+������Ԅ��Y����� ]�ѹ�;�n�Mܣ}����`���X��j�6�����*�樄@�){)Xx�	$�y�v�k�k� �f��>Cp�N�n��8��˯jN��d��5����e�\:y}��՛�j�r=@����bhD@@j���(e���l ��KM��Q%w����Ho�b7n���JTTE��0�ʋa��:1R��fn0��ro�u&v�2�h��/m%�v����9�V���{�����z���t���j��l/�*&@�!�Cʅ�6��a� �KTx P�p��,,m����p�=��b���ł���6�imJ��BY/޼8����®{�YF�o��Z?��[H�,y��w�$4��*J��BN�|C�� ��0��������Y��Ս���f7u��]�u,�ʕ�V+S�(�)�P���Ł}���w�}��_:f����FEU�P�#�n���*!o8�)��˻�;O�I)M4�n�w��������uc�f���0��O�%�]�A*S<Rg��F<��Z�z�9�q��ș{�l��-<`Y�M����ri��ł�M��fI��TN `?���H�rg��M�>1����Z�^��+�.E�!���rQ�6[����w?9��`�����҃We��Z�}��i��/�+_�¨Yjb���?��H�X�\�c'�la���aVz���Mu,H+���)ռ�k���oY[�$�vgq������|e��j���z�W�^�9=׉�Z�DZ�rA�@.
OU��c'��g�b�H���O�F,`=�`h�5=�[�L����|j��;�Zj�qm�>im��r�Wf2$=��������>���7����Y����
K�V¿r�A	�H"��14�JK(m)!!��Q*��Z/%�f�X���"���↟}�����UCU�j�=����77o��׮ҭHu�d��F��dC�o�Clu�=����<0�"Lt����޵2�
��(?{B�¦�{�)������`�A~�����և�i����h_0`Kǔ�?U��j��m^6��W}Gyv�]�;w��o^Au�J����Py�D��P���Eg�p	�fB_���+����[.�/�.\]��a�k2��(�`UuIX*�Rt����4��~���˧���+Gm]��aԈ�nʋC2��Q �B�,P%��T����&y�)_0<B���3���m����D^-o��;��;y~~�������vo����h�AՉ��ՙ�-+�Wq��G:~�uT�ȕM��UȩT��o�.
F� d�"C�͈>�'?C|����a(�V|M�Ҩ',Ww�ާB���-!u�M��J�JQ��+���^Ξ�x���y��8�:U{$]�S̈́,�Ҷ��EA <�dH����g=�F<?�Tx�G�h�*!��S�f|�_�ְ�bv�6��]7��>�R���C�1��&�<���Lj%�v{<�3�=XNk��qV��{EM��o%�Qպ�����~�����u`$O��� �0"V����I?�T��o�_�:ؿs��w��c$��i=�Bj�myW�Lk�<s9�>�>�V���������DP, �pP`�����=e''/�.e���$uO�xH��x��X�ԗ��@�]�A�}����k�������|!����X]f���N����z#�*i=�R��o/�ɉd�`|���y����Q4�V�Wz���oԀ����V8m���>��L��3���Y�T�:q�Vt4��0�yu���lT7Q�S��ꞯJJvx�����BKY���6l(�6��ߟ=~ry��^[y��iѪ��K��	���Iz�1�� �Ñ��%^��D��XoM M��Ɍ7$N4�Vm����i�.�n�I���r���;���i���c�w�,���    IDATp_���ǳӹ�It�l�y�����;�P"G�EzȐ5M���R%1���̏T?7�),!�H��[�
����%V*!�,J��(��p0�f�f!Ɏ�/�ȩO �H�\xrb�K�(��6�� K^<A�$�x������2"6?�
�а	�Pȣ���|6�k���_s$�p_CmhBb[*��r�/H�R��'���y|!�ȏf���pB|�>�)I��	17��gh�]	TLM"� �$��4t��O�<Q��S�֬��!IQ.�e��ȅJ�
�������rVC	�0������ �+?���/������VC��������1Ǻk��?�������?Tm�j�^��tP�QɅ �-�f ��Y����.��Ƣf6�$?�� ] �6���.Db8?��
<���,����h�a��ѝ����/~����N�{���k��<f�BmwD��W�H�eDo�/y��
�)���W�+ujg���V?�4x��^cW}F���k�Q�Mֵ�G���:VIo̖i�k6INm��7�c�Q�M����G]�[�>�V��}[km:�Q\�H��JN�,�5F��Jb*�J!�L�AQM�-� %Q��~X1�c�w�)]Mc�������?Z��+��|������&5�zkj����ȭg՗�X��ʷ��bD��sXBYb*�o��l���ݨ��mO�(`��I}���H?}E�Hy茼���@��[~&�/�9����B^|�Ia_r9��G�e��T �Z?)�p���Q��	rC~&$,l��N.�"����6��Z9r�"@�~��%`�I�D�@�mCS�D&< �a��D�i}!����	`�� �/��
?H ���[�@E!�sb�Fs�)l���*F�L��)���0P�����1��g�el�� @rr*�+b!X@�@���,���#�CFr�ȃ��d!LZQ0�I(alE9���@�%�`�!F``b�䫑%�_*�l�i�%��__k�/<$�H�Ȇk��� %�UL8�0�x4
z�rRv�"hCa
}����a�J��l�#j~���/0Hk`��K�I"9:��I/ 4
�v���@rb�n��WrA%JB2�#�I�p��"�Ǘ�Z�ow¢r�`��0��7 Bx��~\ǏNh�p�xy�9 	9H��Vu�x���u�X��w��Ǉ/�7'hDt�|Zg5Yη�N���,�9�`���Kko�����s�̃���j`j�lZ��p��j7�֥B6f��RY�Fm� #��Bd8M�?S
a*�	S ��i�� ��$�C�b�����Vg޽<s�)z�(���c��No��ͪ;�bSDo���ե����� j1x]��z�,S����y�o�Q��Rm�	ߦ�����+w\��ݱ�Ҍ�s+�1���r�-�����j���d�S����i����4�϶����aT��!���5��$�Z��P�	���0�bP鄋�9 `��>������6�9OP/��`���� �R7�NOL���t�9���ٲ�ͫ��������8cD�+PvP�� O�{{wˌW�6"Y8��4�x�D�����bMʰ?hж *�J���(t��ᵝ�i������s�-��J�m}�T���q�>�y��ᨇ[\7���j}Ѧ-Y-�2��zb�lf?��rory�S�l�oMʣE I�&�̮V���)������
ׂw��(�����:�@Y8�~�q6r]ǰ]ձ�������9%V��Lv���{�;�P+msǬ1��Ŕ�T��lM�\�BR�525{����G{��_�n���@���ʆ���d˲!�utd������;{��|�Ͷf�Gf�Z��t��=���?�-��:'b7�А>��H��Ap�ԙ�6v�㇣~��وm;�Vj��<�NRm.��(go��n?��ߜ<y�Wס�8T����/�"/����o#@��'O�ȣ�����vD8Fx�I�#j����W�L�&t0L���.���
ݺ�Z����wQ#����إ�H1�_�`Y'X��|��t����-���۽��/�z�$V�I/��zo��%[3d���M����c
�p!�g�xM �P$Mi�Ƶ�8������bӐ�}�eBj�A�·���Q���;�yu�}z98�찢�Z�o��mk�N��ju��"�� .�hc��Ri!h��yIb����`�_"��3ϬdUH3ph"ASU�9�QUL�)T&}� �B��JU)CۊZ�t}��m�����98ޝ�6[�����BghC^*�$�$�6��#۰&0�I���8�U����{�wt����b�F:-j���i��R����m�q�y- ]Oٔ����o�Цv���k��i�����$vb�eB95B�� F0�7��W�hD���.08�KW�IVKڳs/_�>�z��#�k̓X� 0�aL4�$�	�Sqm��Ⱥp���;�����"�U7��j���l*
I܆���ӗ#�0 �r�E1��9�φ����3G��K]�jRVu�ᾞ��{y}��Փ?>z�bj1��Q�����by>s~�Nk)k�d�N��|�0쑳�(��DR���9�B!��ߞX`��Ͷ�#9A�'�:�-������v���f�Mx�K�*�5!^�*�D�:
3-��|o��w0��gm�?eԺj2*)4ӁYo�B��
�TĎ���F��Txσ��X�L\e�y6q_�K3v�9�R�)z����±GG==���������'_�׫g�K��*gB�_��.�-�Q`�r!�O-(c������xqGԌ<vĢ_,��?�Y6;���<Xv.���pr燯�������a�~ݥo�AO�9|�<Q-��#�:�tO���VR��n�����M]�y���+�$���DEQ�E9}	��FmЖ�&�* ����_��/�ol�!U'Ej�[z^g.��X����s^��@����Xz����g?\�_�nf{[�P�i��1]u� �l(��5�	u���r����/a:���, Nl��~�F�\��ċe(�a�_��_�v������کƾt��'�eu1�ީN�A�&L���C6K�vv�J��:~t�����V���k��R�$O��.�ȏ��
���d��	��ذ�^[���3vn<v[&��+�
QRg����L��+�I�]Q�v�zx%��%UXmP���S���M�m�<��='P���r_. (���a�.갧�v5���^Mg���\ػ�Jc���!��	b}C�ؽ�4�����~�{1�FL���7uXӔe��V�@v�uc��Y���?>C!��Jd��#fiu���Q�X?4˵Ӌ��1�0����p����q��t6Mǔ��蠪Po��稊�����W�_���:�����k���_X�*B��D���!��yH�]�Wꪫ0�d�jd��Fd�"@�NH��FLp�)�(�=|�~
��+�ʀ��=yszt0��;�챭*�0��Mu�7\y�_&���U�ḆP�;�Xxn��%�,�s=�
Z�� CUTI� �VS���_`YϿ��RnŤ�)@�Up�U޾<��w����A��pֱZ-��S�m�(t"tom���^\\�����z�t�C)Iȃ}���g_#A���/���u�֑��_.JL˨p�:� ��Et�
��PK���k�U���6	�4��FK5z�ݶa��LSS���V�k#l��U���5d*/�Q�*I�K��D�  s~�����	@�hQXH��8��rj��W0?7�����+0���X?E�&�p?#�E��$?An~��d<I�l#��7z�����L}E%wREa~a���	��ѓ�Eh0���F�Yժ1���";�$��=�k��SQ��D H�D,�I"0T� �pHſ�P T\&_?!�Lx��C��<��F�*`���(NB.��֒�j��U"��K�B��X��:K����F�-��QZ~�5�0����={&��m� �z'��&���A�XuNTg� �����z[����7}/먤fȃDt��V�}��_�Uʯ��
P[/e��>x��
�Ç�+3�aĮɕ������HH�Sr"��M
CT`"&�8�@�:�e٭:� >��ࣿ��_}���x�������g��R-o��J��-���T����W]�QtY���B����Nt}_�L-��iк�����N�L�~Pi���9z= ��i����g�8\��(��5+Q��*X�&�)h
���n'#�kſj��Ͱ��AiZtmPQ����
Vyu�T�i4��R/�Il�imPMD�յ��R�]ۛ�O�
��-��ť��y=]���ppu^�v��v���?���|������w;;w~|Q�\��lk�Zo@-�HP[<Z�����%!<��5"�T�CJ??���\�q�(7?��J�O�$�X*'T�-6�8mV^8xHT������#Z���p��Ox<��(H(��!�2�mb��:�p �ٔB`-�aY,�/$��O���|����$h9hQ�@`~J����(@��Å�<I��x�I0�̐����0(6��A�JZ�D�J�@_`<0 R��7�53�p1dl�&ɆB~N,f�)��U߱��&�����5�8� y�F�+,�%�w,�p�aΏ��>��
��L�I`(���dͨ� D,�b�r�%P^L1$B@FVA%w��BF���s�S?�'j`���8�*L���H � 5�Ebx8})�9�K�$�~Ѭ����/�@I0�Ƀe�}��,�60��XQ(���"9Y$�ګL�z�Օ/#�� �'kH���eq�߃V.�L��JZY ����W�~�6O +�VpR!���H^�S�@_�'\ �p�H�<hC�^8'_	[��R�m,9 ������`��qoj�C���q:ݫ7���Z�;��s�8���	m�Wu��4��ӛ�#���<���Bޯ~����ۇ��oֵ�IĢVg�a~Ug���N�!����+� e�	�G��p�DA? V�49�Ն�1at=��������$���ƻ�bM�v�Rr�V�F�t�V-��[��;���Յ'�F��/"7�m*�V��'<[;zxG�p�NGD1���櫞©v{��V���/f���U�,,)v�L3Ud��s�i��p��O_L@��iUrz��wh����p��;���W�Yffq�i6�4�EP�4S<�%�6���)pJ�_�XŁ�@!�O����_��sW��f��22��B�L
Zi�1����������so�v��U�	��.'}�W�A��'8���?|o�49+V�2��o���[g�̨�|8ak�so�s�=���!zK(���&,t��$�dk�Ztk�����U�4�Ȏ�:N��M���Ξ�.g�p�c�{5M���_,���"�kB��B�-���l�f����m3j�$��w�'����z�th��d��F�Z���q��;9�j2`�Et��eWs��<�<��("���j3�E��4����0�aO�(�C*���*�Z0}gg��}lv�(�Յ���,Nm�����O_����gww녵-�i�Y-˴.y[��hh)��V���{�����e	���l����a!��[�5'*�p�'
�ͼ)蒺~pۼh��?����o�@55J����	�v�e-WG���%��9��<�d�-��ɋ=�������aLR�b��=4 !�d:�S �T�K��.��DBF���4�@�wy��?~�ރ>��ٕ�l�=e��`�Y�2�$�<������phbf|�s�t�ԡ b�L+Q�|1���e����
;�,P,^�A`<9<>���o�l�W�-����f���gi*��J��I�==y|6ۙ�v.��j��ʸ;bl�R��l.1F�!�5�S*D�`�W��0�_) U�����{U��Ⱥ;
n�2%�e9e9�y��|���}�E;�_�Җ��}�$!Tֻ�Z�;������w���u�k���#'-R㐁 �#J��پ���	�P ^*�j�撩;�kc�zkwo����a��ʇF#��֛����s�Nظ�nw|������a��g�g��v�gZ6j}����P���:�Xf�a�ER��姽�~r�A���BRx���N(�*�&"��ﾝJr�#Q%q��zDU�}-�G|ѽ�����~�U��ʃ�� �B艟$���r��(~�
JoÒ��fb��x�J����y�L�m����s�����r�ě��ǍUvhY���zk�(�}u�9S�PE������މ�W'L!��Ж���`���p\��tc0e<�r��E?!G6^����c�,�x����u�|͙�R�l�˭j"z�m3m�E:n172��O���=�m�0�muf*��C˥$�"�`�y���Sb�r����8Y
fj��pݚIf�����㻃Ѿ�zOP�^'z�wU0S�*zPUf�މ<�m�(S�Z�PU�E����.h=䬽#I�:�IOPU�@B���#O?!���+``��S��b����Ư����O����O���3�Wj�+ 08�OX�y�W@��]'��Ö��]K)��kK��`�͎�q��}M�zV��"��|��6%ăN�*�o�]�n���$�����-u����������w�k���,�٭�A̴چ;%ǻ��[Wg��p��_}0�:�ë�߽*�L�.�B�![]e�
~�Ӏ��=I�)Q<�XM	`���Ģ�� Vüd{�[��wpgw8�A��;7���*n��e�F��f%�6{g�ӭ=[?������Veu�j�����'�[V;X�Қ5&F�R!���/��y�Q ���P9��@jc��@:�):ᯝw6�գ�e�Y����l�j�Y�Fs9��"g�o$k��w���Vh��B���t[8��)J�$0�@
�~�Pc��:A�(!����	�� 􎣂����\�R�: �,ʋe��A�Tc���~���J{3��������k#���UdO]��u�=老�Nv��[���X�u��	_~���N�!ji��giV�l21tK�(e��Sc�5�j����E���<*-TЫ���eDb�+��5��c'Q_Gщ�1Z���/bx�d�uN�Ħ�T��Y�9��Fݻ{tt|��	�A�.WQ[�{�>|����曋��y�XX-[cl����������������X�;;�w{{�w�A�ng�Z:L�L����n��ԅ��{f,��㵟��k�
��$.�Tk;JV�kG7�dS`�������Dm�FP�L<!c3�֍ݙ5�n��Uw�_�T�H0�&��T�~9��\S�[�G�;;��ׅ�2�#pi���P�k~�i3��B]��e�1�!INb�a#y��HR�m65��t���R6ݿ��Ġr�ܮ��ᝉ��4�1T�����3V;���;܌��5�K��7�s;$k�M9�C�.�}�����li���/�R(���J�rr�L�s��P�Q*HQ�,�����W`�0���+<��oBN���	6�8��� Ʌ���ICL
����*X�G��~rb��H�C<z���ښ#���ǡ9�����4��n�����0���%ᑻ@	yB�\�G� 㮐7O ��W��B��+�)�|AJN��Ud�$!�R ���C�%�Z��sqIb�E0*�/T�7t�$G���I�O���: ��;��������LK�?��<���J9z�,��b?~�)0R�]hq`f������O�URu����Bܱ~B`C�j��g�m���=�E����ʯ����a���=�\�_��z�VMYRH���_=z�$���?f��d��_� �G�C�@��"}!<����gb�JML8������g?x�םߜ>�:{eR������Ye�U�u����vK<������y��E�WX�un%��g��*yqg��xK�[5�kkj��x���	&�1j�S6sǼ��1��w�����֓Q��tݕ�Զ~�z2��qv�-��~��S���7�D�e��+*��h���\=����@Jmk��&�T���b\�պk�Uj5���    IDAT ����c�7W6E.U�i�c��Ѻj��&��7�6���?x��'+OG|ՙ��L��K;���7n����a�.6Q�p��x!ZQ	�<~�7����£b%��B!���[MH�,�MF	�v����H'�HT?���C<R�� 6:b���`��
�p��{ǚp1:5?�Z*�I`r��GC�*H$G�܃sC00Lobᇍ܄��*!<~"�?��Z��%�z�p� ǎ�q� }K&`	�����	��d��%;iy�@�&��	�MFB���	�?0�2
�����Ŷ��+<d��		�$��L?��I� 1@ο �D�s�����*SVI�)e�̾���f�!#dC"���[&t L`$q(!7�P=0���.���:rQ��!�C��V���B`��8�W"	��j?�EIEn�D�f6bq._����K.�B�#d���0� ����@����BI��PA�'?�װ]������S0��y�����n=�8����7?`�K��"J�`�#:����}��T.�e׶�����CL�`!D�p�����/�OQ��E�p���XD�srN����X����!9?����:�'>��7�~�`�oۿ;����z�Έ�b�f��~zq;��c�`�j�\�7����쿧����{�oNf�WM��c���jj�њW�;��ē����Hra�S��)�p-���Q����Y(}sŁY������ܞ�>��i���U֭z���	�2�071֟�?ޚ=��U��W����4Τ^��xW()_8!�@~�HԢ��o���2텺*�B��O+�bww�՘�i5�`�?.MEy��uw�3w�w��;���m�[��I�S�qp��k���oWO�9 ����Nۦ��k�q����ȟ�E�@~�q�lBp�/<���	���Y�Zi�#�zG���U].�=Qh6��,�}_��0�RoZ�(�:����Jrd��eƯ.@l��#p����hf�%��ѳ�s��-��f��d�?f�,'�3+V.P	���o�]�ԩ&uU�Ȝ�>���Hg���?��u����z3��p5�':6����U��LT)�_L\�'_sx���P"U��"9�@R�-�:˥fQn�w��;�{0�yM�*����y3Y*i�4���2j2�Va��˓���q�ۗW�S�Ͼ��fl���j��SfG�ɠ�_:�Ɋ?��}9t��
�Ö�	B!���Le���p�\k�^��bN��l:��tzצ��]��˟��4��X=��M\�������O>������3c���h[�C	�P���@�E��K�4%8B1|SeY]a]�6W��4Ѓ�@ߛ��3	3���V�j<Ͳ(KW�<UGY��X��KQ�e<�e=}��r�Z�:b>1�cF�̯��@6S�(Jm4��&��E= h��m�~vf���9������뛫�?<=yy�񑣗�.׎r����.2s.uɲ\���a_:g0ٚ�E�ݹ��w[��EVi�蔖rxA*� C��G�hk�V�$dǯ~%*_� ��1���Q���+�۸�.�rIv���ʐ�z�T�syq�zֹ4U����/`��/G�Q�K�ƽ "Ub�	�J\m�Hb�A �x sU��g�.�����z� �kbLk�^���U` i
K�U�R;=wmR�3iiAT�t[}m�V�L�Su9r�:�TѼ�Շ<�C
�}��
m�4�*���ߤ�6u�wi�SV�Xux�V��56��CV���r������Ջ��Z�ݣ���b]�����m$j���"�KW�gJd�e.�'�8?1%[U�>#��A3�h'0���cCM��&�����g��S NjH^��K9[��e�[kb�/!��ۺ}b��H������k5��� �A,��G'N	�Bަ��6�05�^��L��C����*A��(G_�Eu"�T�Γ��{�lk/�v�doPo�,$3�7GP����8H,i���Ј��� ���<�Iّ�.�pI�T,y�K+�"c������x_�!Pa�4��2OK�w��:q�q[W^���Z�9�w|�x���V�I��OC��EPHE!:(kP�V�o{ݨ;R�Q4�6��Ɇ�^���ޮ]�{��p����k�]\�Բ8Dg6Č�"6I��m⵪�>��<���61�vG{zQ����Y�M��
/�/�����к�9�6�&R�*�Q#8~�v��ҍzKN�1ȁ�DA��4����&������{w�}�Mon��Vw-����G{�;2�R�i�+�����#�y�m2~j�E?�[�jÝ*�s�a ��`L��/����E�hT	���'�/�v��bY������Tl5�Ye��!䩎�ޕ�	a�*am�]��N�ؿ��~��:<y���˧uyd�cK�d���Bz�}h�\�s�!P��i��W(&QA�^�ɁO�-��M9H���s�7K�lG��#�����{ޟ�^�-��\�LWk�P�J7ОH��i>�ӆo�ۭ�I�������֒�Kk�	��^S�� 4s~
�A<R"m~�K武�vK�'�,��2]W�|���=}X�Cn�W@u��5��xT�>�lp��:�7u�.��5VE �QZȉ+�#�Ēi LcE����(VX<��cA9'�/��I��b�jRҵ��*���=l3��.VVY�hk�e�nͷv��ҥ\�eg|p���G�'ӗ]F�ͦ'��_����_��mC �kƳ��˜r (��G?:�:��xK��'��z������3�D��e�<�>���6��T08BA�Z�]�&7B����o�=}~aE���eo�]ZC T�a!J�A2	6�Ah�QSM�j��_�����z��|��2�6v������M�aq&��4;e��+���vn;�_��ں!�-�e�L]��,^޺�����C�;^3=:���=�?x�5��kQ�os�2B��~_�x$g�?�<�}�%��%v������
��m՝��V�ҭ�+u.m��b��V\��Ϟ_��ڭ"|ʝB,��=����+�f���$��6��[\�>�zя=B��Ǐm�*z=F� ����hbQ>�of �W�5��:�8���w�l�ƌ8���I�\����5O������F���d_��i��ZB�`��[bo��HMd`�� �%�w�?x0��9��6�RSd���a
��)�����Y�!����2~��mI�#��pË��%h�H� 4�2�~
�@�`³��LF`$%0^����0\��S9���m7�)	͗�Dጜuʓ���v	'�����+Ð!k!�����C�h �p!D��<�/����#Cxp���rQ�6H r`~�KF�P%I����U�6'��d��A�p���4��4i#����U?`�����1VO�<�����r���͡Y¤�8⤅J�������A-g�������.��82����������������������N䊃���P��������e	����'5�:x@��$Wi#,ߔ.�RaFq�'����'�p~!��O���fb���[���{��_<�d��9_����ʵ�Lt��vמz�~5���EJ?�FM����(�4�v^k�ڊRv��n�3��9�-���� \��-=t��Z}_��T�Rq��u��^fQ���\ۏpu4ۖ7�%3�J�ۗ�(�\C�6 �ۻ���.��Y8=�j��׵ܺ�!�%�G�����@#T�y�Ƶ�<�e*��.z�.��O��HDAT����"dUU��)�i�ˁIW7�������N��~��ѷ��=]����9�-�z %�f��b�
��$�\���hڢ UF͖�5(�[��O <	LZ���K�<4Je@��D2�~"�O呼J�,T�
r� !	�\�P{<�"�
W'7��!�C.��4$R��9`���R��M^X�G���#	
�!y8.	 ��/mJ	��0ߪ��
L�܁q�40�FP��Sb�Ś/�\��ǐO`򕜠�<��pQ��W.6l�"	a�Kr����9`�@�3.si�I>�hc�Dv)/`���Ml�l��`b�)�<��%_��:����@p�%~���&$:X�X�A�X|���%b	6_��B^��VZd$�IgЊ�(`�����ex�	'/�pr��7� �������OP҂Q.)G�H
�r��
��$:槴B��)N.`�УԀA�W�s���x2k!���5��0�6.e�Z�Im<y��
�0C�1" I�y�/?z F%���s��6�J	"�KF�~�6x�GX����=4�r���P��6N�o�IZ~�$1,1�?�>��Ҧ;bfS��K�w�㛗�ӋK�9XR[�%��^��H����C1���������?��{�Χg�39N�-�N��m��k�*ʝ�!�h;	S`�,ObA�݄'a	�jw��P��ٵŸ�X�\�@<������Τs�p���0k@��s�ξu�3�[��Y�^=���:�����h�[L(���>h=��h���|�>+�vQ ��	ǃ)�#��x3E�p6{&\�h�pw� ǜ�����y���`��?��͛?u�=.�(�~ ��T��߬o5����t�jϭ�4��4ﱵ��W��bY���#2BL?��˅$�8��/	�9iE���pL���5���,�?���z�W�l�o����NS�ۑ[DWj�]���Ã�gU�ɐ��a��}Uj�E��4<� pB�r ��u81�s!$)�/����;���:�YJ<sԊ����:�^Pg��J�z������lj�B�&�
���9z�Qԭ���`\'��ї����������5��ՠ�I���zR�-r ;��<^���З�²;<�Μ��4��<�jN��a��� �Oi�Ч�?�kW3����t�f~�������l�)"����N-H���S�x����J�(Z�z���G� x�5
`N�4z ���x�*I�V6G� K��	ə��6�;��ک��=��QK�@�ԏ��ٖ��M�ŕ��זBq��N�V�����`�� 7�<��]�CG"��5[Y�g���+�9���t�u�}�>��k֍���q��@L�*U30ۭ��*��V�G�'g�lq��8ЦT�N^������ C�Dso�a1"I ��?F�%"U)���*Y�Je}�F�,F�R~�q�b�8s����J&/:B���k�ifo��d]ޥ5���B��Q�z�G�m�Be�k2ƃ.��Cg c���MLs�?z8`h"S_�����5���~�Xӗ���K��
�]����nܦͨ�cַn��|��'?��\\;������\�QE2�R�dj<�ʆ�F���x�D�X���C!�WA�	̗��nP��)q��a�;s�s����N��k�>�f���������+�^u���:�7��\�S�.���2��)wT	L����Ȉ���B`�Y��*�2�*�2�5����:k�L�)_+ie�hٕ��M�=�aw��z���w�z�������]��[����l-�qJ� :_\D�ҠM�pŤD���.#L4{�@�JmO��RՂ�ڛ�:�^�Z��q7�[s�o����W�Ti��z&�FwF�f�)��1����.c�HI���� �/BP�S!�(�IH�����R� ��k�`f-�P�Z�s�Z7�A��iV�
U���-�,\�۹\y��3��|�j�v�I�m�1C�SA��-��J @E���;߱#�4����ٴ=M*ْ<��:�p�F��7�D�׽�͕c����Tc;��7X��pUSx�j��z8&���v�lO��xCX	�V���z*2��$���P�Ӣ�&�ay�{F8���+n"a�n�����j�5�4�n׺5�b{
O����v�x<:�.O,���;<)c��t��ІH4D��A�a��#_yB�=%.$$m�a��"�����0X�����7e��%=���ހ���ی2g����Q���Su~-l֙co�3>�:h�X^�4����>|3ΑI.�D�	��_E�X`~n\��#q�?�����5�����������`D,�������VYt-hoq����>x����ݏof�]IM�+)�9���[S�`H�(�1�ƨF���Ń��+��X3���=0�E'��������h����j$V<���=�O�~1Tۖj�c�o#;�\Ѯ����}�o;<���v���4�g���lF9d�b�7jC>	$p~�)��d�*�aJ ~�N�Sk;l3�U6�*Z�g^j{�=K.J�>1�l�a�ʊ�����jk��+צ\z����Y���|���ʗe����$=_ ��1�j��Z�� .�F��TB�\��lh]�R�C#��c�in�6�[u��)Wy,u,�5>��N���~Zm��;�{pw�yv�=��S��fק�z�NMn�V����C2ZϢ�'J��	��@I��Z�޳e���/ޜ��ǘ�ΰc+m6A�j�X�#
T��F�J[�l��tzf��Nʺ~֜b�"�V���m�e$FPh d��{��Vm�S���r̡ˏ/��l�-ي��mʜ���ZI�Bش� N��\O>�qz��s�܎\kHs4�N��TO��ZZ����U���5���*�v<\i�u�]Cb�j���|�"1G�	a�:��G��W ����b0��u��-�u�RU��(�dí(�B0I��V�IeuŘ�q�]Z�~ua�51}1��)E�P�jK�CGc�T������Q��!Iѐ*0�fmP�`��25�G\0)�6��tn�l=q�`@�^�(����;�Ъϵ��d���e+)���ߞ�����F�"��]%�z�*����h�7D�Xu
;���:�LZ��H�J2?y8�N#U0 ���<d�+
w�E�%��x��_8Hiy�a �a߀�<l0��K��^6`����ρ|����/R�����D���x
��auH��b;��}���Es���o�w1|��i��kѦ��5*;Qx)��[�[g�ċ ����`NB�~��@r�Bx�������9��  3 �ݠ�3��rB���P	��I(� x*�Y��I^8x5BUR;褴`�l<봤$.�U���OQ}��Ç������Nj���<y�K�i=z��%Ny��Z�J�����UU,8i����f�~���>~���@IF�U`m@�V�/ф�8T�����7$tc�����|�~����j�� ��}!O`<��(b��U����ņ(?MuYg��a���?���>���xw� ���|�c]W��a��(ײw5)<M�N,�ެf�Y��e�RS�U$U�:��������́F�4�Y�HT���me�"�k֛e��l�6PE&xYSZ�Q�&_��k��IQ1 ���mS5O`��n�x����*:��X�m֤�aVS	�0ء�[;�Y��V-YV���� j99��U5	#���X�"j}T?��D�@Uc��Z������j�<;o�Q��7���e�p�=��-y��M���׳��D��n���܉��S����;�+$��WAs�L,��w�,~ �	}�'�u�C�n��)V�W��,U�t0G�A��'��b���4C/6_H�$�����Wl�<!N'H��*��  =I���9 �0�� J�3�o��AT &\�@�`��<���"
�@��d�'C�h�Ky��� ����%!CűD\r2� 	��SZ����*Q�!T������˒�	S:y�CR(㧬����+���
��Q֡�Ac�bQȐ�0Ky�0�6�0w��A��3 �J|������eSr�=�M8���ƛT���J�$_��Ă@���6r��)�~rb��T�S�,ȇ2B�@�X���/V�0p! �$D'1J��9��iG��<H9J���1+I�O~Ġ))%��D���C
 ��'�$� ހ��;'S'�]��@��T�AqT�Vy�G��y҂�B�łO` ������&� �)9"�r `.�I�'�RA���� �+F5�s�5�����&[�������ޓ~��������k�4�e    IDAT��Q�d�U-��Ù����}�����W?�����3�(���S[W��\�c���lc��$��/� U ǃ)t
�S��<~� _�`#b��BR�iT��0�P�2W]����5��dZ���K4o>��;uo���}�s����''�]w������8��t�?y��Ï�i3��hCvhSF(��#�z�b9�Bm��j�X���(�W�Zi
BE4͞S������ޜV�����u�jG�S�&v�ڿ�i�}�8߉��5ڋ�V��D�&��@,?� V��9�����dk��bvy�s����7��]+�/��Ң�.L�|J���=8������r��z5?��n�ng�lp��l	/�ʗ�$G_�	�诖�M��?�;�����{%�f4��9���Yۛ)��"H��Ts�s�LT�e������}v�v�����˪�k �X�4\�Nԏ"���^�;�Fj��n~�jn��3���X�zk��z�D!G�0�q(���̣E�0���V�!5�/d:$�L���Sm�I�q]�)�k5-��9�1j˄*����S+�I�=��έ�ź�u��OB���UA�s������$9\�M��_�
�f���� 1}���:��x���2Q��pT�Ҽ�H_�&@�X-Ϊ�ꪮ:�-{Da��oYW�=:����K�������n�V��&��@2̗�c0Qmt ��	_��0cȈ��>����m[!�
�)�!ڪ#m�����ݳ^�騺���؜��wx`�H'I�C�O�ZU"ea���eD�cC�T�OtrX��*� Q4x�\���VݱRF�˫K�\���l�S��]Y�7d!c�|����E�\qmz��z��Z^qDHɸ*J6��ۛ��� e	�/�$*_ $}��J�����d����FuX��a�!����VR��`��h�?��|yb�~�1Y��� ��5�J_�2�nJ\Y5I@z� �Q*$EI���=�ė��F�'/_�_�
��T6�\�.]�X�\O/l�Yؚ���D��e�b���][�A]-�����������D�R,"��bЉ�`�UL�d�w��U�i��5��j���4�L�%V�-u֭�q�fc�<�v�u���v0:9{�����:߬�����LG��S��L鲓)by��#s��6EE0.B�/L��@�x��k���U���>���n�:�3ov��ȥKÍ�M��v�G-��Ij��6T�ܮ;I�w{������i��	 ��R(=D�� ?�J Tɶ O4�� D2K�x�0+������L=[�v���]L�TC�.����ة�8f��O�{Sg��n)��H%�4TS._�K��)�TT��%g����f���E��$���C�V��v5(
�2���sԯOO�k��nC4qxt����X���A^g�pJ�c!7=a�`˖��F��������?�\1¥��j^�CVA �8,P$�p��'�Î����y��`�ji�.��Lv���>���[-�vOG�Um���v��K���X]k�G^��AK�=-�.䦬���O.~bD lhK��S �����Ŧ���S��@܁�b�M�z��Z`�:�<?�����裛�,V�ւ�Ə	�3�<Z]Ù�蝻=���:��������SֲVKj�ƛS�K�^�V[sCK�e��j��^iH}�JN^<��G���:�=٪��V�j�{�����\�����vJ�Uh�ѓ��~�������ǳ�k�8�n��&�eD� ��ёd8�����ɐ�2Ƙ�v�>H�)i3,d�MH�ą���h��m�[&z�n�ɢ���v���7�7�C�2mjѬ9�TT-U��3�7];�,d&&��]Sz�7ܹ��u��;�C�ve\���v�5�v��0L!X$͢�[��H�F@1C�A,T���{���$U*Y�O�!�鬛aZr�+S���nݨks��7��Nփ��I]#�5!�v&[� �膬+�F�Q<��d�"d#XI��?�I��Sd�v��κ曋�7g����G���`��{�=��Rh�W;�rM �}��({��"�7=�5��B �����^ܜ���^�� ���Sɱ4��s?�D:�X��!,�u�U͗7����/���oož�@l�E�Ź]�:�Ř$�*����Ӵ�5_��׍�H.aV��"�p2ꍌD&G���4�,;B� "C��I_���Sϋ�&B.��F���^�_�F・��u�Ի�_%�#;�\����m[/��-��)э&�~���^<{�Zw�^��%�m���Ň��u=�}�[`O��Ek6s_����v���:����J[m"U1�'��<H"j��n��^`\�tz~z�Z�WfҞ:���{��)M��q��R���*W��͸Og����+}��8��QT�!Fֺ�Y�N�jE�� ��>y��E���E��Qc`lcq��5���!	Y5�)a;5j�u�}}��'ӳ��׵���9�a�o�T����d�o��������X��{POh#X^%����|�PF�l�P` ���g�MZ!?�@	!GF��3� 8�I(N0)��J�s � �V����p��~�L����*�	��R�A��'$�B���h�+lv��zT�j"�й�?�>ƞjiN7�����~�YX�\��2�Z΁Tp��#EɡA8�����
�:&*�`Q�8�	WA���%�X�cJ��P�^���ύ�@�p�VZ�}C�T��M^ʈǗ��	��,����
��&%:�l���~�;K�(/G�L�&D*��D���F,��ީn*`�!�����#xTU$��Ւ" CUe��O>�R�cҀ?~l�Vʇ� ������`	̯�k�!� �țE+'B�|#>t	K��A}d$!HQ`����kE
�5�;w��#����������֮��g��5bG�&Hw�Ι�����ٚy8e�]m?��o���,uz�d��P�����޸@�}�dT��hĘL���Ui6fݼ_��z��w��|�����s��x�mPs/&���@�k{�g�͇��%��JՈ�����F�oU����Ik��}�j�2�r���vW����98��LR��kv�Q�pcgY�m��~Au�q$���̪-�����\��~�M��ƸI&fG�A)hڝXMo����\ig�R�G�����{~�߿�ۯN�]����0T�O5"�}P�E��=𥻔��y*�e�'I?���AI	�D`P)M��ѽ"�U3����B�' �ȑ�	�������0+;(P��g0�%Y��l�-��H�P��F_�d������J<p����M^`���`��I�//�����_rQ�dʅ�`�%����
E�	���F3��̅�P(//¥��x~���?4��&:��E�l�eǶ�b��0���S�˒s�e�r!����j0 �#.�$�D6:Y����E����o��V������ 4ڇM�ڇH���e�sp�Ɗ��sc��B�	�>b���91�$��N����$�G��^����I��{O��\{�Z`��%���'H�������B/����
Y�L� �;;�Lw�L�?�J����7�UYYYYYYY�"KR��5%��T?��s?!��_o!y�~"~Q`�c�� s��!�~Յ~�P+J�����a;N*�b/l��.����kH�!!�V�T�p
/!����Ea0�@=*�b�1���N�����*#~*H�Up��Y���$0��8���U��+&x!�TET^b#��8��G`C��	��` �by*w�%B�+Jv�Y010�~��D$��|�t45`@Z�d;��l���݌GL?�ͷ�?��d���p����I��.���˟���G�?�������w*��t�=1j�F��z̀g#w��H���"	g�"��, q���R�R�V8xN�p�\����1�3�5��xl1��r����;�ܸ\ S=Y�̾�T�LmsV�\��&{�ه��>���>�^�ٜ���0�:W�"Oe��R��':�$_r�X"~�(���O��?���8m��b]֩�"���8q)�\K3������G���O�[`�+C8��鼛�ޛI.&��39:���3f��F����x.\l�I��Ĳ����/���J�+D����N>��5�Ɩ3X�A1�L��1+�m���1ڃ����f{綄#���8bC��NeԄ!��
|F	�?�P,E�@_7��s#��OvY&Wǧ��Co�M��Xq���z��]Xi���m�oLp�X0�.��w�x�`޽p�*<Z,�@�L6X�0%�m�K1]v�|���k�'|0Gֻ���a'�n"�A�8)#tȽPҖu�K	z��?�m� Rl��d�z�>��7&1S*�?��hS�Oe
t��f�{� �r��9<K�i�PaJ�}ƙY�°�^=�b�?��-a��K��N�����յ!���0�T�!̴=�W��U�/�P�=R�7�0��V]-eu;��Swpz͝�7��8k6��L��>5ffE1���È�������+��n]�����ŢRڤ�d���!?�pR}˃r��OU��c�b�̴��d~�t��v�^��N���	�6z��F�W:�.��G�����Ճ����}g!�$3Ȑ������1�(p���~Y��xBR�< �QI�;�S�z�;K	�#Um76�e6�p�o���|�o��������K��t��r�=MCU%�pAS��-��Z��9���p˴R&R��M�"!f�}9�.����T��G'H?�˴<B�ۛ��x��&���?q	]Za���^��]�0d��|��hy29�6�9v���˫s���
Y�ȷ	a��(^|�d� �WA�$=��x��b'!��p(�R�,���ڐ�̕�j�vսN�q��z���h���#�-3s�fEigu�>}l���]��b�Y����h0B�)�Pr��n����T�!�W���n5�l ��V;G�p얍�ݓ�����l�(���-~��u`w3tP��ۃ۞�t<�/��yh�,Y���or.E�4�Kx��/QT��Pv�����b���XʁG�� ��Nȕ� ���?�7�x��k�!��$�枇?1x��wMop�<a���ֹHYg��"T�aw6���(C���h=v���`s�ꆀ7��ϣhE'�FjQ�� �]B�{�I���ܸ8�'��;�a��>�"#�O��}m���@���/�?�n�^�����^X�/rр��Yۗ#�'�UDXJ�S);QQ5��Ͼ�R S(rΣJU��,�Ȇ�m@o7˛�o�O��nL�ɝc�E5�,�;�hv�7��t���؏ǩ�L9���,:Y����K��f���%�`Jx8��d����m���x�m��=y/�>�]�-��W�����%ߝzD�Z��j}��Z�P���� Yg�?�s���%�H"	���r5E!W��60FCH��5�g��DB�I)�����S��F��_��Mw�3:����R���b�4�a��lE��I{� f���tc/���żqn��6�[�t뿪�/e���n3��D�T:��H�!�2�B�" ��H]l������ы�;��d4!*�
�D]0�����T��v�kfp8x�Г�={���<��7��?ο��_;|�ʲ�uڳ����BJ1��&�h�4D򗬚"`~��X]�JJު��@�"� P��I~�b�iX$t-�o��N�ξ����C�7[+N��g�����&�T�:�����`g���^�sb�k�gri��QXR�X(E$\є٢�;�R��fZ5R��k��L�����~�r��[��+O���BO���q�.�L������|�r+����/O�	��3�0�9> _�I8z�R���|�=`B�L�+jDT�/���N��趙���K:��O��=}����\�)j������S���j�+/��O�G��m�2��v��zW׹�3F�5�����[��.�h��4^�Szpr��I�Unz�ٔf�wrz������|u�"bs�>Ӽ�1�`��H�QA[�>�S���7qD�
i�ʉ������}*E�,C�J�Q%�QH��Gk{�8x��ɣ���gݫ՝�:��ҕ�����Xz�*��2�OՑ�=*���<;����I)����>x�����xv��'��ϟ}��,�ӝa�9��VE�.b���rsĭ�M�]��=yz�۵G���01`�N��c����͖�hʈ
�<
�\���%y�K{Q}��%Tt�4�٣ÃEVR�l�n�u9�ܬ6�d���m:���ͽE�է�w>��sY���o�*�"�ȝL����fΐum�BDуNE@���ڦ���Fd����S�'� �(&��/M<�&ÀT�þ.�@e<���]��7�D�5��n�5h&�\X�'76�>�=<���;��B��c�ˏ ?)��\ԝ���)�d��R*$q<J$\Z~�+��}{�
$0���o՗o��< ����X�
���g*\�
,��D8��� �Ȇ_a+�?$ x!��(�ZaPe�jMh��wz���ht�l#��\$nv"J~`���ڸ��c�&�cu�kҶu;4[Ѿ;��:ug\J�]����Hɇ�"�xO���L���x�c ���nY�ʼ���W��6T�u���%P�9l��/He����R;�i��VT�R`�p~��GIU��xdC.D�"C��V��0���R"0�@DY;z�ڞ�_Ӊ���?G�o�[H����(;hA�cwp��H�!	��Jwǚ�(�EY1����h���# �_�D�/~��FQ�u��T�@��p�dC��hC�U�+KH(�u�)X�S�8!2�[� _]5O�ޗ_�b��k1�4�,m�Ӥ�����>z����n�����һ���Q�e���k"!&L�����i#5v�M����auk1�#}vW���9g%ڕ&���$�A�g��:�LBb��e������2xu���Z��zt�#����ˆ1���!+����ɘ�G��4!k	SW�:�v+#/oD`:��C��j�J���|�g�(Jss�7Y�{�v�3 W��ۥ�����KJj��#˄��Z�U�v�`��
9Rx")C&�Zh2M�@'?8��������M�V0��,�gG����P�<���[.�<I��ƣ~��$��pL B�[Fi�j0��J`J0��9���%��$W��J��@㯖�^,<ڛ��Z!�+V*�ࡒ�=��,�/��~�<��T��(-T��5a���� �hy8 �#l�FF��+;��`��A��� #�b̲.��K��	�_r�{�@�Ur	Q�/	' �`*�"@ ��AV�?D%I�@~8%)̒c��������{��iF:��/��I�r�R���;�Qp@eG��B%� ��0ˢ���E��c%<J$-�ܑAW�*����D�(�=U���	/f����?,�],bxda�~٩b���Z"��䲮��%Q�)'	v����W>���{c]�-gJ"k����Td�	���?�����y��~�V��,3�
�Tb} ʕ�ˡ�NG� ��O,0���Z(�8�u`2UM����so>��{UB�RQ�-�Y��UM:���_m��`&���$��G�� 9~h�y��
+$��[?K&E�`Q�% ���}\�y�/��DU���p���6)'�C��&�Xx@ʢ���_?9��B��+!<�hRe�~�`�Dz`��V>��^��bF�����?���۟��}�շ/�8���o^��:���ɛ����=~냧{����g/�N�;]����NM�e�-o����7�Rd_#1�,q�AL}��Z�!C�ϡ�)g3�$(	�
_x|T�&~��m`b+�i�ic둉,Sh7׮4��9N{��Q����u�#ǫ�����=�ݼ�4�9�X���8�Z�C���5
y
��K2�J 8M@�q�<�D�*��K� XjN��ڑW�|�ض�����l�����M������Q�	��c�w�s�ȅ�=7Bl���&B�o�����U    IDAT#�܋{<P!�<��6�
����D`%�2�����|�p��O�,�5g��!��>�mUԺs�k�ִ�����tXβض��WɿoI2��<���o��γgo���?;y���=e�<~��;o�EY�%��mo�nm��� -�Ү�����ɣ��Yaf49@����?�����`}Nf�,�I�[OQ��],��ml�EwL��b���d�T+XԊy}J�e[D��`��*H����/�"CT����/W�SQ �@��������\�f�5�Y�fjٹ`Je慮��;��;i�����4��w���O�-�$�i$��L.t��30�#�S-�cy��R =@¿"%�'�H�g�����b�;��vw:����|�a�=`cQ��2	mԟ.Vj���w��J	��#Wh��O��[r(Ō-bP^"T\�T�6�*!2�U��̰���x�$����ڝ�5��NNB��^w�6���t�i�vc�Ͳ�v���7���̶w'�(�z��K1Z��HBa�����a��U�/���lq��&�eo( ~V�NNZE���V��i>&e��h��?�������ugs��N�Z�3ϒ�S��b��޲���u��g��8�n���xKq�)��kmQ!��%�=��EG���`P��G�@J��2����i0L��)S[V�"uA�Q���Ň�����&*����m;X���KU.J-�F`#�
�O�U)��K[W����T���oq�fQв����=�v �H�6\��nEZL�$�t��������G���a~;\8_�6I[p�t2��E�bu��ޏ�*K�c;���Xͣ��
%��Ej|m��N2g��:w�WQqΖ渮�)ss��}��7E�;t�<��cV�U ݁�H��j[O�T���L	�u�fH,�]u�;`S,7d��T��+��ڬ�`*!��R�Jd���Z�^��>�ݬN͍!�v۟�g�����h�Yo3���]u�0��g��Q1t��M9�U4!��ϕGa����`�d�d�{n�&���9ܝ��S���j���5ccff���K��T�v`��� ��[?�zC� xLhZ�T
��!F:A�#��t��<�a|Y�Ujz�ST(�p�V]����"\_F�Ef�3X���=�|a�����h������|Iu����������}�p��d�{��p�1��R�����d?V�f(n4�*n�=��Z�����K|��[dm�1�?��t���oo����5�����r��� �x3_C|�O81?�w�]m�!���BJ%���H�Hȏ����p�c;?�ˣϤL�^�9������w�|��7o�������t����iϛ��ec���d~â��X�b���/�;��O����b{�\����|-�	���o1ɓ�_}���~���(*��=|�7_LmK�t��w������H���yL����g�/��䕉�ћ������ܥ��N�*�P��<(�-.!��iI���
"\ @��7�i�3�mԉ�$\�z)`Z� mᬦ'����ۛ����<?�R�Ȁ��L�$D�(��<3��u��^\9b��F�"��&��˂M�+�r��gX�v~P}�,�X���b����*N�D�������m���޾͙B�����6�����`6�^}��l�Z�|}��j��?�Er�VC.eG���f0G!�C6JJ���W��] �S�y ,��H���O�G���JG����|�⻕|et�rH�N2�0�w6O:�1�w���U�U�b��̪z���;����c#��DĨ&eD��4
�R��v�7_}m����7��ho�5PgR����(��9����X���K�_�ăa0�wG7݁�������W9"�ոW?�p�Pgs�����آ�b�7��:\��-oro����[��D�$/��vjb1���m��۬�	­9wooq���/>ɜ�������Φ�+({�	7���������m.�ƥ��&
'���Ӆ�<F�T �G�JZ��+#_N�Xy:9y�ӷ�B�@?��T��+��d)����f���N�ɗs>��X��X�}�y�ގ�M{����%^U�����
4x�R4���@���Eg�9 �^�T鴍b��
^J�l>��������{�3�y��kQ�=�y{+N,iJ��d��i���N��R�[���y~��Y�.��)2P�'`���Vi�K�S�p%����`|E�6Ri�(��Y�&���PF��O�+;L7ڨ� }RF�����Rp�E�8_�U���z��
@up��+�\��� sMQ^ l���664�Ӛ7����t�;Q�h��L:�m�+�ě��g�ј1��ە]�F)���j��a{
�"&�c��w��m�Zs��e�[�/ ,�Hm�l��堊� n(^j3U|��_e,��)���h��pq��r$���2��+��co%��k�J��<b���j�G��<��Pr�c�F�V���	��Z���;�J��ۜx}7��)V����7����~��8d�YM���裏�	ၐk���?��r�[o�%ɿ���g.[(�t�x��/K�'��A2�����%�@��(fL(��yx�W,�)���=��
@�e��$��D!E	���R�g@�)t��jw����w�������x�4Z��H�J����hȓok�8a5�Ș8c ���l�Z���T]�<ؐc���{�h���W��F���q�Ŋ��٥�k��-Q��|{z}�$#SM�����p��c�����g3�ts���92�'{��F�K�!F)�ڙ�3g�=���ld��63�c���vgֺv&���45��^�?�/fg�Q6�d�Q����D� �3F0ߡ�̼h{ٗ�³i;LVw������o�V�����x{����O�`Z��WK{~�Ν&�9E.լR���y���(�@�� oZ����G  ! *D�
$�<���� L�8?���|+!�+k�N!��V�ʫ2�$�:*V8�r�V�\�.�a�J`e
��W����a�'H�%0�H��Y�K32\	��XmPT�P-K�\Bx�	#6�
�� a���}FRa+��c~�H"
r0�_��*��
�Jr��|a���0?����уdr���V	i'����:
�O>��O�s�@�#Dv~RS��&��h�V�$Wp��r�>��c�UFfd Q0JB�����S��~�R���##�I�f��U:��
L�'l
%V�K��O?U"�8yax���V}I�Q�
^!Xq��=�Ph졘��G��
� �h��S.0� ����T� ��Gr�WL	�*B�A*�Rq�D���׿���'UISՐ$��{�������+d����¢�Gx�W��M�"�`�Zз	�鹠U����A�l��p�	Zd�����4�<�C�,�_�ax(<X���娀� P�<+�B`C?�\�J���	:�rH�I�$H�,�,�*��\*aU��iEU���Ul�M�ȚN�.>YvG&v��~��;��Ë��׎_�����>�{����p{�Z��O�^z��17<��oܓF�]O 3�a�2��(j�_�����8`
@?򣜇l��|����Ue�М����8�)L��0�҄�j��-�(¼C�=�����oΜ�qʳ��6�F[k����>��|Ax�L��	d��%��9,��r��D
g����b/;d�$1D��nF�+���l������o%1�eB2��+w6ZB1�i۹���R������{]��Fjx�4-O�� a%��ɏ�ي�`*��_W_�>v�~�s{��Q[`_�#�<T�v�F;P��.�xE��/ӏ&��u�p��Hp Z�Y�@�������`�k���Ç�]!{������zӟ=\�=0�?�\�YJ1�`}{� =+I0ܗ��@w&�)���<�g�������n���<���Y����fj�+�֚\�������b�e�A�ŗI�:��j��	�[���
U<�K����ƃl�(YT�$(�怃�d�|-9�c.�@2�>˲���b�����xЛ/G��\�ý8�TS�jl���,@#Qb��6K���H5��U56��I5��z[;](�hx=�G[��Z0�W$���Zjf����|����9�9ʶ>
�*�f���o7�Ҍ�,��5E^\�Eη�E�	خr����q���boq���
�b�Wr���$Vq�B�8t;�]S�Օ���l�gg���X͙�����T�]�8=y��h��CZ#�S^����`�>0f�9�� C��b�@�,�*�n��ڦ����v�_Mu��⦐��=�v'oE���BdL2�&�(��l2��qR��;���)�k����#p�L�֖a����	Ȗ�O��-?^	̃B j�>�~@�������:ݱiڈM�A�i�M�*�1��6���LΎ�i����ȓ/W5�z�$�@-)E��8��)-I�U�!�@��Ь�T�$�^�ᛩZ����닎�RN�9W.�`!�f1�E��9T�[TGSׇ;9��*�I�����3z)mB�*H�Q҈IrI�TA�s$� �v�5��1�f�R�{{a�Q�͍;����1������oO�����بr。Kҿ;y8Y0>���[�s䜴W�C0�3&����Nv�/�*,Q�*�jΚ��wWޘ�\�I�mbݳ\ =9�Ǩ�Ja��<.v����RQ��|�.��Xv�4N��ms�Xd���d�����<%���$�M��]7�3������<r�ߩ7=��/|���:#3��D��9�iSL4�Ѹg�{u��ś��0�Z���֥���8�0X� ~r���< |V`��D�@J�=7��=�sw�q���9}�ß�l��{`�����ƈ��B��L�C�on8���|bDT.�2U \1e�,h^�_?��(#Wx ����sZ~�]1�v�C�f�Z��+ș7&��J���;���K����ڹ�۴
I���(�����Hv@(CE��!�^�h+�����J�*�PT�:�$�.�j�e�w��79(�3�M��хs��lҙ��K���reroBhr�9�E�ⶋ1�|v�E�]�e�����P���r;%fB����V*+�{Ub|���*��0���/�O��^`'�h��,<d8��=�j9��ZQ\��-������ڼ��q������d�<X|y�����a٥M�H�W���C�z?�1��u`��ɶ�`�� T��H�K%�/)�S�͊!8���$`�4xT�Pwna8{x���1n��6-�d��=9�~�:k���y�#g�ҙZvNOi�i���Db9�s��ҍtC�$6���T��7�b_q�#a��UZ���=Z�S�V��"#���U����8v�N�Z��.Q�N�q�ҵ�nܓT�Z ���(A��XW*]l��O����:��	y���)A*l
��osM�����ӫ�3/	��D��γ�]ͭ�'�جh���F�^�(Je�_5dl��ljj'j*]m��{�m�i��x�8�Cm�d+d�,�
ݣ~�	1�f�8r9���ƶ��"yآ�"siԗ�b�[y���/������<{�8��nB�? 	�ܵ8*���������o�NvN.�D�f��Ao�����S¯	|��;��� ��"�"�'�jH���X���2u�e�>�?z�@��r��t��'�7� ��\3�6}؎bA	�Q�E�q�}[�	?��{�C��m��T �$9�_��SV��$N=Sk�БzД3�ժ�칗�[��'��h~�|u��إ���[�RX�~�jb��Z�E������:"a��l B��$B��BP!$46�Ei�~r T�S��gꑄ�K1���Ǉ����^���w�]Kh+]���jo�ľ&�i�9������G�O�Υ��-��_d��mh�/JR����L��r_�`@J�H0 �H���)	Wy	"!X O�TTa�pQ��G'I	y�"�h��T
�y*ַ�T8�"F ?����Y~?��G�1��kӳv��[�T2������jn\�4�Y[bZL�����̧�k#ގ���="A��e���_F'xyտ\�Y��7;K��ʦY�ş]`Цzh�i�
ȃ
�
 '�j�JAe�;��^%Rg�)I ���!�[�� ������C�XQ<`�,mqҷpJ"
<�V�+�B�"�9H�9�ȱRf~�}	�#<'��4>�g�_����>�L,��.2}m���K=8��������ɂj6����~�+��q:x)w4Ȉb��/~������?���7�GRQ�m��/��/���/�KE�7������O��dÎP��(�)r���Y��\Ð<��£�ʏS�Y�*Q�9����Zl���Gs�>�w�����>��.NY��ʾ/���1�X��jUd'C�(�U���D���Hu�i��OE1Rʍ�4GQE�dy���8�vn���wW˻�[N�fþ=>s�eq��K×,z}*w�d��c4���n��;b��C)wZ٩N��sNu�;��6aE��<����O�5�<����x��ýݱ�9�O۝Y�t]	�]�gS����,b:n&��v�&s��&5���`n��cL�Z�M���LC&|(�1�M�m�ivh���������������H�7����t]�nǄ��Q�+'�Z]Ƀ�j3�K�.���x�0�V�#�\0�EUH�ܣ��x�T���������M�BD�st2
'!EIE�p���˫���0%�����z)�JxOjC�F�I�+JZ��G�쵂��oa+�
�!���d�'x?��U0�ف\`�+	0Y(>��E �A�X��0?`?��JQE.!��{����o�M�QJ0� ���R�������/�I�١h���\�SY���\,���x1R���/����SX�&d��B�����;��D`hQ"�>�����G bd��.����9VJ�Q�C��$�.�)������<��;LO �e��PA�@�K�x?)g�~�!ऌ �WB`0�h@_�y��jhx%�,�stf���_���O?��F���D�SG��	�ʢ��تߒ�rE��_��ER�7�" �W�8Y�?z�Y!�S�*�B0 h�`&?�~J�!��@�-
��E���/��$~J�<2��C^ ���Br�*>l���@�x$Y��r�T�� �XQ�0T<��*���*T��=B�y�wA�`�⼝���������b����x���w�޸�p��bog��>*j�:z��13�sv�}y�>]�.>�
�.ʬX-/�Tu�J��� 8!����]D(��,j��5	+KG>:SH&�����K2�t<%���2��fnZ��#M�pVwo��
a�3�0s�lm���_��3�4I!
˯��~"�V45�N�- ��4y U�U�q�'L oگ"dﰋ;��N��x��a�;�#9T�}��m9*��!�@�gE3��Ow0�s��d-;f~s��!����1�Wl�G��<�� |%�ҫ"�(���%��f�����"39C�n��p�)ʎmYÉ�6�[Q��z�ɠ����%0��N�9�s¿�֙�/�PES��b:7�?=w�>W�@�\�9�O�N�R�KZ�U�������E�3?���|���^�pus��K(ɖI����:bbQ���?ɪ&��1g�ca�6�"�Ňc�gp�ɜ�`��+<i�C����?}q��k[&�];=s#�Zjm�y̶M�LE���g�.�y{�ibM'
xr�~yrꆫFTT�,�Q��Jj�����ԎS8J���@�4 �T5���J+�T�,�\�5�Ĩq�;���=~�ƛ��[��/ϯ�=�i��֝mVk�U
���+�h��K�� K�`��D��eͣD\��nB�!�O�"C�ɀ��`[{q7�Eq֑��ɜ	�T˝�*Z��e2Z�	l:gw����do��z#E�`4$)��#v)�|}iRJW���{���td_~��    IDAT|�|v�ɂ�3l8Q� �`�����-�Flc]lH`��e�,ґWuuyY�s7�Ln���X��k�=ܙ�YG����d�M���2��2��t�&!���C��q�(R�B�*@Ub0��''�#`o��n�B4�M�����p�(a��lQDf!�ʍ֓���]C#�"q��x:�dFK�)���ᇇǗ��
3݋N��9��&���
RBᤚR)��
D?�yl��cF;��(�����anX���h�5��L��uc9Ŭ7	���*ɭ�;��jV=e�P��.��6bE�r��$�	���-C���G��z��-��̘��z�>S_9d�BpҝRym��C!0�Moo�����{��G���l��M
��Ƌ���P��Ӏ�%��!Jp ��+sd��Ry�3�]B%�z��O�+����$��!�0�.�	�<?y��������b�6�MF��Cc��W���[����uh���r��8�/��=x���&�(BQ¯P�]�@NH0���ߨ�N�۬��X��<6��g�����n�v�1~�|�P����fЦR��J.7���Ν��^�.z��`B���d�Qj�OO�5	'��+
�q��Hi�C���  �� 8��*KEl�������./�O�x�w������kn�5���M�6e}Y���ZY������0��p�F͢Jz0
<����G!��Xu!밴�����"�p_:*e�)��b;�x4�6����ԧ��e������m4p���l�ӵvnj5J[��	���bʝ|���W���Ө2��b�3��>�ѯhR���!��T+����lD1����/S��?x�g�{x0�<yu����E�UK��T�+v�(5���{h����D��5K,L��8 2U�b�oD��8J��t��+VƢY���芲,�y/�mt��Y���=t�:;��t"����d�I��Fav�!u��u�p�r�������k���95�h'�Y�զF�`U���Z\�aU&II�!����'�
A��\_8_G��t�� 88qyvmx6}�n����9������۝ i>\f��d��8�<��	��k�c0���q
�o3�B_5�����A�~e74P)��g�%����rB�`3���+�mCɕ���!Ǝ�B���"M�i-�O�z��<��Jl��*���E@*2H0��a�"��0�y�)�U�B.�����?��J�����}sou}~���������;�n�Or����l���(JV';�Ϯ�!�n {�V�W^k���)�&�H�te����E�o�^t�\�ZL�7�T��â���f�Af��(ƐT�ek�B'�v06�m	r�u5j����>gc"G�/z�5O�T�4�/'[ �;��z��1�H"&�O���bk��r!U mC~$��P�{Zwo��r{���٠
:�݉{}���l��.�L�����%.%ww��!��x��a������5�_ʹ�jF��}�
�B�Qa� +G� �uI�1-��v���� �.����"���"�e٪��c#/�q�cO��]�#s�4Y���NG�T�\TV,���1�A��X�KE�!�w�U<�������T�X� I�80� TX��}O��N����ڊi4��^��#c����3O�sY���F
�z&ias}+{,
?KW�IM�J��J8�����O�U*?��/�p��
BY��B�ge�C%PIPU�� ����P~I�!�;�*�p?ʨ<R	,"+���W��*�����	!���Ȋ��Q�N�bh�����3�����֖�����4�9�ˌy�M	��[��]��f�����Cmt-������2�ڸ�}tqc'q��b�w���Kx̰��:�d:��a0���K�z�J��Ö*���"�[L�a�,⑝(��9�=�}Z���aPH��˷P�(8��=�j��.��p�G�JA��`3	����H��A�(��(�~�+�]��t�+2�X�,(C�Hz�<��A��W_������ba���o��`hڙ�������Â%A��$��C��_�姟~
���ڪ̊&R���b(`R�H�Ze+�Vr~_`���3�I@�-0߰E������6r��<}�G��Ǯ�?;v <#>�]6�edn�1��E[�+u���O���g/V�-1Fp��&r�k&��u�L�uW��������٩m�����ٝs�ߞ._���Z�cw�������<T�3���lA����g�k/�k?�Q�ɠZ�l-Tk���HE>�*FW9��g��"o؞��զ���|��{��s����G��|�9ܟ�$�k��D�E�x�UO��>����9�`��2%��vyd���e[(Ef��n&i15K�y�j*�y��������������w��o�g{����^��juz��Wjx`���x$��GM��%A�%ɧ9Q/�P���g��4W!����ON�oJ�fOH -����呪įR�܂3oZ�r��f! ����"{��J�%�V�+z�l��ɶ+$h��C��h]�~�E$����` ���*�r���T��`��K��$0� ��-b sb9ᰉ�ʗ�P��'WyIRQ0�|R <4F�&���i:�Ja� ;��?�)���T��h��,E�K{b>򔈣����C�	��d�LŁg�ˋ� �>�c�������#��Bʾ�;�$���J�P��/�U^Y�*�C�q�:�E�@!ʋ!)��a��� N�J'D+dT��8�2
	�A���NjZi�R�
TG�Y�`��PF�&�ϪP%so�I"a��Ѧ�B�T,�"��������~[�bPʯ8�^�O�*S��,�+����A���p��[��	9'��(x	�@a�B0�a��<J�'H�K�\,����_�/�0(�����/���D_!rQ�` �@�������ŗ��_�y��[?�ȾBd$��B���7J��O��"����L���WH���	?�M�d�Ry���bi��{m\e�U�ko��P�J����nN�����V�±m~r���@	"طx[�B W�B�D�B(t�]Ҟ^�զ�\9���g�����m����g��chaƜ,��O/��v�Ogz{=�~���Bg=��s�[�UrG!�T� �~�E?	! *N[C�M�I�3Y���*0x�k8��6�+9�x%�Y��YӇ�2��ۙo��ݞ�����70�s��bH*k�L蕝X�$�HQqR������Sj44Y�����p��y��o��[��<L�u]��ZA��q�\��ZL�2nt���-��p��p[GĴB�Le$<,M(�Nƴ�R�l�'�)�C�޺�1�˘����d��:�^��j���a���԰����;?��f�!f�����WlF�iR�'�[;���'�T޸r�9p���ė�^��a@��Ⱥ�h�)R]��%iSJE���go?S���B����H�)�&��K�R��V���U�˼&��3�\����3�0m���Vȫ�"{t)�ЫE%�6�[������>�I��ec=H		��_��2����]g�c&�� �4�Lѫ���"b&1hLf�d�βw8�O�yæ�|T�)�v(Zj���@�H���Q��J*�&UU�,�Z�x���U12�ve�m�!r,��e�q���r��tt0��v�.\T�}���N"�U@�S�إ�W��W��/ �EL�0h�U�����'� ˘)�F^��	��YO�Es(�����K�L�`���^Xȕ��t[�ʌt/++�M�r(���;&D�$�!�K�&E0@[N H$q%��������"�668Q�em+��)d�Y��.�d��p��颿{�=��SiZMʾ��˳u;�9�8ʤ��d�Gg�
�X_ꗞ�QG��b�hx��&�E�B	,��HaM�O�;���Z�^���;�����Jr���h�6�l3��z��Q�s�K��;[sF��,?a�g�����{ɽ	p)O!��< ����qS�)���^�[y�F����dM�ۚs�w�ꐳE"S�F���hdY�sr�:���n��p���W�eAWc2
I�+��Sb�˻ﾋ�dU*U  �Yt���Y���N�_4�>ַZAq�)�]n:�=~��ᓃ���p�U���l��I�Ʈ�f�i������d��r	���+�oɎuz���ͽ�qU��J�~!(�Q�~��Eh��i.��?�J��y@kЛ�Gg�gҚh�HU�'��z�,aReъ��y�^w:��ַ����ıK�����"B+9���9�K|C�*WqX	�@��*%0��'"y0ux̜�F���\��+�loڱ��Un��YD�ƃ�b�K����G�ͬ�@�|��Mv�$�+E����'0�B�X�8y���&rh�U�f�̊��\�ey�9��� R_�y[�[��L������<��bR�;�����sPh��؞ (�.��U1���Ch����S�� �$�Ɖƃ����ݾ��DBE#�)1��p/0�.�3��n%��c�n_�һ�+�(�O�	�3B�yn�W�W�KL�XF̹���r��'勰*B������0<�c�?�=�9�&krc��y�C1=t��sP^vX[��
���у��.>���__\]|s~�����f���%b��	5�Ъq̌l����H�k]�I;��?%)!S���,�U�U~�]���c�;|㤍W��=��g?َz�wvztv�2Ϫ��tGY#JKu&!�i0�j�xt8�� �w(��1\��ʡ��Zt����VE�c2:��KX��&q�������ޓl���Zծ�鎕ե��f�.͈��W��t�Ww�ߝ�:�tի��7��Oɨ`{���;m�*�Bǜ�=Lc���|�U��
 n�=�ÑǁW#0h%��O������H���8��}�����{�����v�)mhc�L���R�v����̛�cU��f}��0^��޳��m��L��"<m"�_h�qp�m��
��`P��KmPdj���h6:|�`������-h�Φ0Ob�T=u�A�֍�����ˬhS�����)�U{�X!wY�>0!�g ����ܘ�k^���?��~JK����&���Q�pF>�S�\2c��s���7�{k�.�L��@�\]��ͪZ���#���/�􆡛��NaW��m��l����ae[�J�5Ǧ��A��T\s`
�(�G���P!��$�
,��P�7}7�8p��.[BҸ3ݺ�}gE��ZO�{yu���Ȓ�v���.�B�+Fɫۗ�[ �� 3�h�Ir�z%��E����
�D�K�(��)���iQ���ђ��3��	�pw�a�Q��(��#2�,W>:�ikD1J�rA	)��\Y ���-˗ �%.���A*~�V��񽯗¦^�%����V��-��v��������XTI�S?��r Q�[}ŗ����X���(�Wj�Ъ��ԡ/lԧ�3H�̭����`����v�,��<�ga6q��,/��풮�Q3n����d��T��@U�_�����ǖ1ݾ����a3X�=7��vY�K��R���t���\�ptvqI��� W�5"�4E3ueH��"MOx���V@�������X$V��
�Nx�
,������g@Vr�9��pE ,w��(J�K���_I`�}h_u �ᔩ��W83I�����"S�ϟ?7R��>������ۿ�[�^C��Hh���_�Ag�U�B�0{ߧL�1�^��������Lv+6t(��Lz&��'�'�����-_�#٦ׅ@� �c:�Q~���(K�6�hG�V�2U/:���f����7�����w�<��B�c&3;\��ξJˉ��T��em���e�i��h!�������c�=@���_�@Ķ��hefW���ǧˣW�߽���y�vZ
˒���A��3�v�G��+��$���L� #�JnH����ف�j.��Qi��+ocl������w۫n�L^B���k$�9w�����������ӇsK�{�;�zx]´�� �?ZL�iQv�B����l	knTg����A�8����HSI�,�ױf�zkK�K����i혙R�X�s�������tgq큖[#����~Wv������q$D)����?%X?}E���/`�yR������VQ<��/��-B���Oq�9�ZA%�)'6�凄��^���.�*����$m��*����� �WB�� ��WB؊�
��p�l\�/!�\�*kȹ"F�L}ˉ.��E��l��$���V8H�� (!�2���#��,"U�(��a�D� 
�6��;J�J�����$�[9Jȩ8�|�E�h �'l��"��Z�e$k�0���(+z��H���W�� �G $�=U.dS���*UI���O?��H��;�	��/S�<(�|et�C~��Ą� �0KH+;�Sv�#�������Ta���#JZ�2�Q��O��>���G�T����B����%�I��9\���(�R#~4�<"l̩�,��4 ]Ƴg�Y�>���{_.��T(�A �/���@��3�!
`4�W,�'� Xq8h�%穌*/���RaY0�����U^���}�%&�ǷX�.�i� �ge��E�|���#1�?��#�Py���a�K(9䲐? �E	^U�-!��;�&��;�]^�NrG��N��-��,��'�͎�|�VZM�@{a�8/2� 2����\d�_��zA0�b�S���	��\�Q�+UUO*��v�a�^}��L�0@���Ձ	�(`�Z�7������cdrw4v�䮷�,utb�����Ԭ��B���6�(��/M���_D��.�,$S� �u�%��P+  m1f��OE"̜�(���I[�@ض� ���5��Y!dy�7s��d*_�j���c]]�h�֩t�q|j���	�K^��%0B�^ ��*���\�� �:eV��G9 �E����ԩ��l��c�\zic��弟5!;�ll̬�G#C���ic��G�!(�+��0<x��hi%Ľ���)���ȁ��6,|�[GUI�I+���u�/O^Z�\�5߷��,��iL��8��l"S����^fK,g��Y>6waR �)�K���`VУ(��x�ʪ:jM[��%��*%�AM��O���@0���e�؍5���-=����7I���y1�;���ڱ�٦�z����L!'�X�'�� �ΧT1_g�p��x¬
JP���n������K.	��Q�@?���f��{�|m�Ӏ�;�?�*�;��F���IO�s�&�D�������6�bTR~�H54�v�a+b! � �)��Qd����˵Z0g%��ٶ��G'G�����87Fe�-=c
e2Q&�Z#g; ����T���v����;��x��b��C�EԚLe�9-���pH�Y*t�c�/�	<I&����*SG 9��W�?���Ű���5�э�*��,� �S����Y��
m� E�f��6eL����	��ϘG���%���hF8�q�5�b�r�`&���9��@���)�X� 1�WU��^Z��2#��1.��37�aj@ǰú�z�ŝ'���{���j�Փ����W�DT7�a%��f=xN����R�I"�ʂ*��@i[�W#����?x`���-�d������]g�,�:�t�>��;�(m(���7�&:6�2q��<��A���L�h�b`�$O.�����������X��9��)��f�Lߎ����c.�;��jp!��w.Vν��q��v��θ�d�����T��E��˨�F	&�s�0�hZ��?Q�����lQu�V$�iD~��G���P�p�Qe�����݊����޽���]M�i;�o9k1G8ԧk�^���9�ƀh��p���P���W���UHI2y�U.4#����H���f���W=�2������Y�l� @�s�D�زA�vF����d�wG�Rױ̑J��v�׫>�F��G�}e�cFU��W~C��ϟ�i�b�D�|m��WJ���0��z    IDAT�2� u�6L6�6[̇�������e��^U��`K��K����/L��m��-�1ѣ^�}��<Ȑ/O�)Q�#�B0�R��p �5 �tD�d2'�
�N�4b�%�Q;�i,�l�p�Ӝ�]�ٞ�..K�HBN!��4���Q*�2�9��*�@[z �0
��|�I(i{y�`dG/� ���9:_]@ N-ˑx���v^�ʊ�?��������ɵ�	6++�,<�2ۺ�
��t�ʝ����DJl7��M�5�f�3уH�/i&78i�XQ�[~!��-[���~U/`�� ��V?<XbPΚ�2���jgY4�h��#[�ο����������`L��T����3���7ߢ��CO��&7�D,K��`BB�`& &@ٿ�P@�j��(r(o�����\-8>ж����v��;Ӄ�V����.��j8s�ٚ�-7��ً[���WV��a�A��JS�w�[��p3�9���.��O$A�t���6�_[���*�(���$�f@�WY��$���=���W���幽+��p:;Nn{�\7��S���Լ=���$C��	�z�I�{e��"�(�ؔ����ar�0�G<
%ז�y?��)�C�|����ڟ��yD��;�;ts��֘�C�a�	�M�Ry���&����vB<�a����Tz��1�Sl�[�J�r!��B`J-�O�~���xpf]���&�ؠ�{��y�v/u��NY�4��w���[��k#�������*9�O����n��3��k��z��b�ķt�ݝ����d��,�^-��6O�q�g>4:۫I�F�~�a�,�;�m����&1<a��� vfO��ON_x�\��`D�h��k�L1�w@1�����y����=���ly�)"��M�*�BRy�� 
X O�
a�n�B8df6[8tu�$����S:�	zy���"F��|̸ۻ�����?����bi[d����U���4#�Ku|�&��(��]@QGBt|4���hZ.�*i1��HY�E����ʗegy�$1H0ˈ�z6Z�w����fS��[�f�U[�Z[֤�,��@��T�	����b�o�~"�CF�42 ���o��T ����0��:� �������U�,�U�E��<E	�b���W�I�������W��H(J¢��TK�W�p�\U
��myhrKFΝ������b���ƃ���HtI�X����5M��é���v��U)�����"F��>>�s%�Ԡ��,}���1-�c�����J�ٿ^�2��'��md��Av�8=�M��xR\���$U\�o~��{���
 ��XԌ�&$���Ī1��\ ���K�=��#�X�	'ڤ��*W,;端�"�@��ax��9?�_,�֬���?���i���~(\o?������{���߇��>�����8�ɂ�B���h���1�r�;C�����PSR��P��ɟ�ٟ���?�bx�XRUT_k{JU= ����R�^��SK�0�i��p�l>{�g�]�m|�}�������q��<�:=��$Mߟe}2cاr4��/�I�DE|V��P��C�1�Ry�	����hSz	of21�b������sO��\�8Z�\n��w}s{b�P���>h�a���#F妚(G-MsE�4:kp:e�w�����,P� ۔�"�uR�.��+�.�eriY�/o/:7���dm�dy��;������jtr��˃�����ho����V鲭���I���,6+�w���5�R��t~Y�D�>����)"�؁���ͦ4�|�x���>��6������{�G�}���������.i:�	�:�hh��C�1a�^b�0D�%$��#�B��Y�"��,���������c�%W��/VYTx}�����,��3��hRT	��,��+���"��]K�"W ��^��(YW�����R�O0U�UvQ�B?V���W��x�6�W���V_?��>�{x���oa��/%XE@m�����0��_����#����~�,��.*�Th#c�4��%�An�M��x�n �(�*�?��sd�m�Z"<�p�B���6]�[�k�IpV1�a����OL@����G���90]���9��D,�#DY�04@+w�G,"5=�� ���$�� ��"9�9T� �/_4���_!/���
%���JB�:}��8�����𳾐% qL��~I�ᕊ�+8�DY  ���a������\!U�`���(��X!�)\rᾒU��%;�T:x��
+����X�>9�
�A,�^��_,'IE�E8Y�V$��l	/�+�r�S�}E�V�0�;�Yx�.w���t0y��;=סAz�G;wO��ڠQG������g����������f� �d��"���&x� tI� *TQ��B��*����J��W�g*��3TLL{s�S��'���Mg�8Yr�'T���<6��*W�X�ʬ��70����n����nƃ�d^.�i�����ո�h8~��r�U�Q�D8�jb����/RJ�h5�f�TP��-#زE\Cp��ej���Z�8W��F�K0����L`�&K5��rk�2�~�[A:��wˢ�e��׮�3��+���g���.�<���,��
-Wz��o���+G�UӷM�#�&)Y	l�qĚ�\_:���,"XFf�ؑ'�~�)����kfW���C���.K�|t��H�`�H�#��F�������4Or�c�d<~Ӧ��a�r�Mִ4�ݱ
�v}��5{�3m�g�d	s� �ug}�/�W%�u�4�тvx��,-W��E�9��9d��˝$��X�Z�4=�6� כfi��%枒�́Z��9H7��΀�R#G����ں��[]b�K` T�r,���%�����?�����/����I��w�`����\N���;G�N0cob)� � 2"X��b�#���F���seN]���\L���r��8&�'<ir%I\*�5g�I8��T)�P����$��w�	5Ӕ�	gK5B������h�M�ʩ�e���W�����#�D�un���A�u�ʃ]�7�䀥���&�(��a��R�-x0�&�К$n�Px�K�9���O`w�LW'7�AϦΉ����N�yN/ޑ� �8D����XkkC�����q�u��+��W��@"~���E����u��DsU�	�S-a.jM��T[>��{#:KZ_�����L1����������:���w�{�ŉ�b}i�������Ќ?���#W���_\�Cg�k_�"�3�T%H�I��x�������5�ξ�O-��qJ�'I��9ͣ��US��l��vNޱ�R#M��'�v*�2�S) �E�@_�)�+!0�T���-�Y?���Ԇ�=��!�~�fb3S�n5� �v����v�f�~���l��
�7l��eG��L���g���W�L���!	Ua��)"b�l�@(��)!`ȯΎ�[��d:Á0s�B$K��P���<�3j6��%��m�pg{f���T�l;&e�YSo,����
��V/b�W `@���}��fm������ ��/s<ũ.e�D8�!I�N��Lf����L��lN.-��K��K<�O�U�<(�4��j��!9~�7�d�� ��:X� �d�I��Y�pG��F?{�&�"�=i�Xn���9�ޅ���}9��9�E�N��e�(r
ﳜ/-
Yjs��RhM�@���ʎN�pQ+k`���G�=�p.����ύW��bf�6�|��n��%T����U��Lw�y�g>�L��S�O�����I#���U)=<7?��㡟��:�j�����@*U�f��*9��t�j�6D�M�-ƃ��N����Y�n��;��!
��g`hʬp���ʢ�v:�+e9����;W+�c
��}
%;?J��u����;���qugOr'ǝ�*�2�2�.�}��)�:�32�d6������z���Ic&���]������@w�hԝWU���%��"#<<<<<<<n9Hb(�j�Rb�?ֆ�Q������\1��6���ړHL���pw���R�e���{Ǫl�mȞw"b�C�h�ˏ _yY�/��1�^���/��R��sI"c�{����8�mE�ˀȩ�Ym��]!����0G]�lڲ�aL[�eUɎ��&�}K毲�Ӧ��{+���߱4
6BJ�-������M��'?
coy��)�8�&�"�b%T"�Ѫ�����؏9<<Ng�1Q��jK��8���6{S�o�!R�%��+�0�p���~B�
�%w?�1f��xK@}��L�Xy@�()�� ȈJ�v�a�	���%n�3��&F��F1R����G����+�xp��-�m��j��W�*�n�K"1�a+�\|C�p~H
L��\f�p�4RF_~�����������=n��o�vV�)��1qp������ �2*�g���jE���HT��m��n'��M�P�m��n��~h�<R��%'�{��E�<�`>�6�fD5Þ:E���|�3��34���?�𣓓��i^mq��4��|k'm�v�/�X6��]�>��t�;��SD�>a �Fp��W�,ƒg?�N!� �ɾIԄgJ�}�~��we���C�l5�A��O������s2�����������ߏ�f�:�$-A��66���A�q�"�>�y�b��I���?�$r��(%c�.P���L8�~�b�W��`�ｽ���\��>~���w��d�<Ȳ3�m:d#����v:3���	�b����M�@	��R��T"�j���֓� n�Z����X!U5<�D�Tpk5�A��q�V��\�(���'"����
<��
O�T־��R�ZMU*�)�0��Q�㤈߆���zO˝;���J���ΐݜ�X���9�4�!3��/L�#p��n��f��M�iS��YĖ1�
�T�����u���d��x�6�++;��֥T�����Ԏ�YѴ�ij�j�+�\=��&����㔗�p��R(R��0���C1�$�gq�7d�o}�/`H �B�<RI·�?�K�'��kJ,DrNr��#
�I����՗p��$�/�=!�`{��J�ڠ5Kˋ�Q��4Y����?�Pٟ={f��w���ma�3�����˪Y�4����fغ�w��eh�&�!��aG
]��9�	4�o]�g�o��o��#�7Q5��7�@"K?y|1eB���kQ�\�/�/6i��=�5�d\28���~��qg� �:���F
�
�!����[B�m��x��΀��L����Q��grng2�c�CLs=�.o��|�̳�u>�Ȇ/V��7g�ӳ˛����W�����zcƬT�z�؈�וR�lRk���o��u���6Ic3�W|��zCf�n�� ��?���F/�^���3Vl��9�Qk`�ܲ��ڳ[,o�|��{�ݽ]m�R��hf�֯������ -Y�p�S n��L
+��錫��Hs��m �Gmez0�Rj��T�Z�5@*[3�k��O��n����یٽ�����������m��3�����]�Qk�K�7�l�b�<  s�ȏ���ZI|EI(���/H_��Gl�f�}��A�6����B�g%/�,D�� T
`�G8O��]v�8���=�~��+2?"a#З~~�<�5O)5�eZHD�D$ ~0��'i"�������������<OcF��X?�(|�4 ��*�?�B�����g*�N�_Hщꌣs���J*EDϰ�}��E	y��Wv"U(PZ�F���i��Q�J���*dW,	l���5}ᑤ~��^B?%)�fr���) �Vy�\9*2#	N�0ڼ*E �Uw0à�(�WpF�r��v� C�W��)�
ʝGq��J�5$2&�*O1G.�p� �rI�r�@��ո�*�p����)�줭�@
He��ϢSg��zI`�ƃB@r�R46��(�U���$� PRQx�K~��PօD��w�K����J�#��T�+j%���QB*�b,"q�	<R�	@��A����@Srᕵ/W4�/����S�j)2k�UZ��r\��ob+�τP߭-��P��A*�7�A����˞ž�{�	�"j�4�#3b��&�L�!����D��D٨�tHF�R�jDL:���}���8Pd���+S�(�Ep�Qx�M`���X$S�02��ܡ!L�I��`ޱ�6eѓ�i��Oͳ�y;�2�|�k�?�CB����AKR�H*ȃ�@cG0���nS�~*D�A+�g?)��9�!�:��eFe����
��96��1��.�$� C�����3�J��ɮ�M{����U&ד3WZ�۵?���Ѡ8�5T0�E��mJ�[� �IF8T�;���j���3tn�A�7l0B�Ŭ���<{�0׬̮���D�`
�8��m�E�Le�BY��\�8Tv��f��e"*����AN��ע���R}��RG�{�'L^�T5�^����������J�Ơwt�QL�,}�}�*��2���͇�_���]D-+�f�/Z~qu~56��lx����}�&;�S,A��X���c��?u��AJ�ˁW(�ۃ�c0��ĕ:�v�mk3Y�� gǋP����υ�Fo.j�XN2�@���x!$�~���E����'�R�bq2}�h�â��	��ZH!��5 �����˪�VSvd���0��ܭ)B��.7RC$�1��.����R��cw�=�jV����X�Y��}�9� Vt"a�b�TZ��b*,Yv�=���`1�U���U�1��o�躲����r��Y�v�f��۳�[��k˥D�-1�OA+�"�����)d�H�U�N,̔V�Tq��+V񕰸�C�':]scs�w��:���zem�ۢ����YH������0{������f���EN�.u�X��:))�.SQ��{'V�媌��y8������u2��5?�<�� ���to2�h�?��N<H����������o^ a;�h�`��>��(
'�ol�0�p�r��� �/���H`�B33�@jH�	PD�gݻ�?�h]Ϲ��_��ڀ��#�6{�,c=5��	{�dn�\��U���h����v6�ܣ��M9K��;m��x��O㡐�O�x��R`��LI�����v-�l�:j;V{��Mw�"(7�V�
u.���2$��L�;^�i˲�6\dMi�v��3���$^aN�2��K$�� ����X�h�j+jA�RH�"JB�W��� �ȍ�v��Y�u�b,���)�6���0��z���F�^z�>vZԄrd�@�f��KS�#a`��N�%�a~�C��r�~�������|�Zz��8�<��F�oSp�̏�u5��8��V��c[C��a����Q"f6f2*PA�NF���)K�Y��>��Q�xuQe���W��'�ɅA���V ���q����&�=mJL��o}���lAqLP÷ΰa� ³��@�,�]���pZ��Z�U%겖2��э�ʫ����x��X��ʔ��I��(�t��J��Z����y;��� 3jK���}���M������Kx� +������\��R�T4�a��[=�~h�Mr�T44���)D[�P�H���-��nӥ&����Ӥj�z9�,S)r
o&���JgB�3�=��M��������͘�.5�%W���@��	����W����e�mdO`��]��8g9���~^W�ֿ�k��fw��L7�]��Ѷ7G{ۖG����l�g��m;��h]��2��!D�U@B��C6ƖeR��J��"B�IB�D�U�@BN����%@�Ԯ;$E���qb������s�,8v�F�Ғpk,"���4�'��p��n����4]�����f9��5���B5=���(~�	�7��{ǐ���*�r�N�3ȭ�8n��3���D�C��t��=��_L�K�K!���GIi`:�
 �D����!�(��"��+W~���|9���څ��-mD�5�Q�$�-� ǆ�ry    IDAT�F]���π��i����^�h'�	<�0q��6GX@T9��H.�����So+DI�i��-V�sh�-�Y�,
���an��-6l�;]z�%:ճ�B$�v��b'}Po�����:�s�7�b�g�RF,�A���o���
bP}bH��c�0чj]���{���|?݈�����4=2TɮM3�<Ъ��_�e�u�{w2;l��cj[������YI��|əE��3#�s�/��2+�!Ґ��6i|�;HGm�������R4=O�����.�����L�|z��&cKs�ڣ�4�+Ԣ|�����K݉�5�����>���o����*�X����R�j/U�%��3�D e�+b��$��؀�Ѱ�I](K��CՋ��y#���b�WB.��
�ǟ|�{��������a6�tr���ɔ�P�6K8&�,����	m �+�M�+��+�G�S��U�
�V�
���	@�<�(ɁI^?}�����B���Sx$��''���:��2�H_���s�S �@Q<�$��K�s�|��������������7�����l���w�R������`�m�&���kg!�2����������0�lK%j<��;)� 칰4b,�&C�M�������O̕��Q���~�ǝh;IF�e}�G���bso�#4�������-y�W�������������\�G)!1A�*��W���� ���*�o�+!�U^��B8�B~�g�c>z*	$���J(05UMC��}�@ʨ���S���)�W���f%�+����/��_��5k�qQ�`��?��^}rvS��7�����mu�����!��a�d�i��o�D:�e�\���A�:M�C�%�*���շb���o���ę�#�4��d�to��Dڽ�����ٟ��6/���(�E��X�ՙc��<m�.'���f6Fbz�Ȳ]��y;þ��lF�a�/��z��fz}CzM0��@�Wϯ.?���9���N'����X���4�b>hu+���GC��vT�2��/+�L�[?˵�L�)u��$E�LlW<��f2W�HTX8���F�5��t%|fwˉ�6s�Fd���b���3�y��������M������:�����\3�e�)�(3c�R��ތ�x�;S,C3�5�Q=ZA��=��iK��f�6����~w���8_���k������_;��_1��bc�A��ռ��o�v���!��9R�������%3)uk0aHs�����Q#�B^��B�]�9��օ���TS�Wl��|� /?���1b}E�H%��H��V��Yyで�嗶b��^Q�@�(	 �\ᇹZ/��Y0bK�Z_6����J3W�\H1$� 9��?�K<���x*w�r����0�(U@ɰ��5ʑ�J+k��AR	��~2�i1��H��a��䥳)
Q+G��QH9�	��2&u;%S�Bp$�(�@,���~�JΡ*`���!Ӳ�)��K,�H`�CEʂN0~BhↃ\a����w�)��Ќ�rA �<r�
m~ʚ�E�K�3�����V�W����9��=`8ɫRp���|Sg�), �J��j!������PM������S��/�D  
VH�A+�Hȃ
��Z�+T([0<B ��o!��pI ���[}+�(��?B~5m�A04��#������K�+�|���U(�r�W)w� /��B�#UQ�'�T�()D�B��g�UEX�Tb��!U!���-��k6�U^g����N 9��l [�� xdm����&c5���M{o�(b���M5(t; "�?g�PJ
���T��HTq_	+UA�A]4$cr'��KgF�W��V��ׯ^�1���6W�l^2�e��ݳݬO��,�:~�����-������*:�t�8�n�j9	��b�؋��d�W��D�&,�@�*E`9�T���)=`2Ęls���ٯj��[G�{ۍ�K'-��B�e�a�j�k��~�	�=���ί����̋Xm���rD0���$I���(&"y|����Oɥ���M�I�CW��	c�v޷�F8K�*݄�%��ێ�d��t�[�L��=h�3_^�j�p�������Nچ �7Q���J͒��U��d�у*�/]��P�Ȧ�_���	��*�R�����w���������~ta���k�<�|��L�f{�"kLo^��v=_7:�c�%��Z����Ʈ��* ����)�����_N)*�H`����yn-��x�c6�x�f�:�vAۣ��f���8��%����k�FJ+�з�Jt��
K�"	�b)$'Ea86�g�: <�[��R�z�Z�0y�XI0$Wd_lg;;�������ֺ�78��m�w���b��zI����5do�#�B�mQ$���0���.&�@wrs�7��$G�h���`u�D�Y�A�@��EᆴU���ZO��n���z7y��g�fq6�H��XX�'٨�^�P�9-�}�d��p��ٹ9M��(A�r�Wc�/���a8�w�a�4�Hc��S&5{b�\�j�J�o��0I|��*��i�7��7�����`dN˶JBDOl�4I�]t+�d��d���vrkM��=��b�kt9KTRZ�V�ʈ�J�<�*?�����J��ip����6'����5�te�R�v��w���`�T�Y^/���3O�>~��kg}���R;��b)Vd�q�N��:v���}EVq�5A}o��,�T"��*:�������j��V��O8����`X��W7��G3?h��_���Hr��n{�dkcB�_�,�f�8(�*�;�֒;ǃT_�����ˏ��жݪ(Oe^���p�V��mG���ka��R3WmY��r6i���><>u�ӈ�x	|:;a/
qN�lr �AEa�X��XLj`�s�(�Xx������,=��W+��$ 	�7��o��%�T�Vwc��Eg����k؍��:2��8�k�:��9'����l��{���!9z�)C# �>��������Q�XT(`ccj$j��
�W��t8�R�חӫ��c.��Un�	6�)��4�kMVP'&"�k��=�v������i~�`�6蝳(>�hi�I��Ø��b)J�9�`�R�"�aV�Fمx�N��o4Ceh��sb��p��S1	ZGO):۰c��Iybgs��I�:�iF��A��DBf3l�67ݳ?��j�2�ei.^�a��!��r�;O����[?���U.��R�JE�*5��9��L�7����|��n9�~7�J
��;,�R�n���I���n��U���ו�9���u��������c)0��[#!]��KY
�H%:�'��s�/-��)�$U(��$d�<;ܳ�8<���{�}��v���3"c��E�����ӂ=��fr�y�|�;���'6���﬌�].����F0#?K�"%!Ȩ�hV.��C�p�j���O3QݦI4���L�b�D�j��.�jf�6�K����j?[V��ۻV%�{�����kr`�������6<�-= ��=���-��I)�ʚV����b��ٽh�h-�"��\�M���M��Lv����p�c-��¢�
���EsP��f!G7��:U�w�R*$K�	{�R�e��WnLY�JQ��>�ACq�9���y�*/"� y���%D�j�r���l��9�0w˥�=(�Z�rj3�# $]��������GtQ�E�ؠ�/bp�xXZE��%/��@*"Q�g�I@��BeT( �*0�!!IC��&Nû���#yg��-p�X���ͽ�4}��<�n�$b��ͺo�;sR��f�`;&0Y���C�Y��ay����~�ժ���
A�Pȕ��(�p���"S�a�I��un�v�1�;�W�.M35�L+�6�-T�L��	�&77���Gn3�Pmp�[.�,�^8v��pI��/b�K{��)^����dO�����k�Q�.�֤�m_�P�WC�_]�#g����&o޾��!^�.��s%�+$�?d�,&pc��\�g�ݡ{qzNd(Gwzf!7��h�S��_�&���J�i����WhV�
I�vїXm���X�F���t�j6�]���p�Z&�t��eւ�����e�����N�۟b/x��������D{S#��J��j�)�P��ϟ?G';�j��PAH��]���	a5�7�Q/��_ٙ������0*�7s�"fW�����qV�-bY�B�g���f轛�
!W^IP�˯�AX�r��<�X��\)Z��ܡ*�beQ0�$�C�SF�	�'&�s-2�{_ �-=�g� �yG9�̐(&�#p� Y�)T6	Di�%K8X��.����5�������㣮++�5b`��������<�Ķd#���W��N/'o^]�����������x������>{J�J)6"cP��bҳy��C.�ڷO�;:�?:�^>������O�lfg�ڕ�]\֤�EK�;��bxm�6����~�O���v�����T��+�L�q�+�4و�S2��ΪͪD�K�!������#��s�%r!����AB�+�֑�i����2-T��,s��G �"�3]`I�RH_4'# jMk���/���Ϥ����V�2'"� ���
�����S��D�VCe���`��Ҫ^���,*�X�+��_��O~���錯��Zf<xeS%T���6�K��8���9�-�tY�~��?:���������7�n���LB��mj��}�n�����Ν"��r�A�I�*S���n7�l�����]^��_^�x�z|���ۋ�w��W��y9��\�&�}F{LD��?��L���#9�B�~2��		HU����캣Ӳ۴C��2�I�g��\�K�����QBE�OfWx��*�����9�h�����_�Gʲ�}�������h�`��7Z���f׉�S�m��Bg!f���QO��a�M��H��^#C|zlS�Tm�f.�U���gǡ�噫�?������/��mNV]w������k
��,i��/P�└��`0�X��᭧�B�N�0���@�b���$�M6-	0�T!$IDq� �ǗFr02�U��1<��
��/���$���
Z��,
��W�(���/k~��놵D��G�/�� 9
�n��Q�JUe�<w�����f�0C%���$�����V���$�<�� ��;ؐ�3Ig�m�B��!�(��
���@��<�+lT�_��_QA (@��%��#_�Bx�;�(;�E���4��L`�9���:��~�K�08�Ər)<���B+��>�RS�0�)	���o~���
�g?�Re� �ô.�(R#a�Q�f���~�G**0 ?���x�<$6����
���,#��A*�ɫ��_��]���(8E)��J�/`!� ���-~���P^\�*��<
����!�
N�-X[�E���
G�$-���W�~���<'�*�$��(ӂ��NQUp��,<�I_�2.����p_I�q�# 'ܷh�P���]v��(`0K^HD�/�* <�C0�R	ޕ������+U	�"H��yԬT`x�^<�p~6 ̕��U��� ��v`U�*�$�+��*  2�A����aB��TEU�/�k!�&���OC�tK��Z�{�����������������=�y�����������1��^L�o�]���z�Hu1�>݄t�5Z��T� ��y��@$2�+�(j�ȶ6.�+j8u�K�i!0*B�XPVUy8� �F����ōkh7vG;�ߎ_{�4S͆�3)��'�y0�](�iU'���k3{s7��2��%/���sdc &��ȷ�rSd���S�~��l���7߼x������Ona�.!�@YwU(5�ƈ~/�?��N�����:��A�ε�ĭw�RaV�6����BJ�b,�q�u0+�`�B�Z ����;�M?�PU�)0� �_�cnh�#�tm���WG�7�ǄO^�g��6�������i��W�Y�\�!ӳ�7z]���O'����Q�Aj1��Ê����Ⳅ�S�q�j�*�����e�wV���Q<τ�Αaց2�h�ի{��{�ltw�����<�LJ�hG����EK������[?Ɓ�@��<l���#�B��7�*t��iT�U^ �#&p&C�~���1I�5���g��q6����++\F���3͒1mV�n
SL��Y�7�ˤ��l��9:��tq�`H"	0p���U.t����	L���b�c�{8�#���x>���߻��z��l�U	l5�6��S�!�<��F�ß<z��x�7���N�g.��p?��]�E�*��!�pI���T!`��O�
aHEȋ�b�����(W�r`�6᱘���#�{�x`�J��f<�{�)ǎ��d���Z�܏�oc��׹kjƫ�i�v9�,$�I���h+6�A���<b�FJ����5�F�y��p���$���g�������vQ���������,�j�ny����^~���v��]L��g���b��Q��#�N&�x@�/�(��E(�TA�EʱZ%j��v���Ue0+,�Lhݚ�N���������Z�Ӯ�R�H�V#9��pm��e�Z��[�,�݁$�,�,hS.N֜�b,y Vl/�ؒ��?Ք�'��A4Y�f5w}s��@$ݬ�樑	:���Zݴj5��^����]_O/E!Ʒ�g��}n��^������TT�%��䡙K��6l1Y8�����Y����Y,���]�}�22�ޓq�Ad�ɬ2�$'&V6�"Z7�����6;�.���H�[���Gd�(��&4��S?Q?^��J�H0&���c��;�'��9S�CǕb�6h�M��*��L�&��Y�%���?x�q���뷛N�7G'�k��o4y�#�|��J�I~����BCW��u���cD2F��d�������`��D�yT��5lv3/�� vN�-Qg ���8Z$��(��Ɗl�^�\N��eG���ʝov���.`,j���5��_�*VC*�W`Y!T�?Z��#<Lvv���j�{Dnm0ʤ]mщ�D�y1�Cw���?xT�����G�� �G���y�5\&q6rj�x=�#~�R���>NS�(p�0��h{������)�	X��SbOzƭ�͡����(=�h�3����W��m��Ϛ��fK����u�^���8��6�+m��t�����d���Ȑ��U�����X?e��3��E�[�j�\J�h��<s��J��u��*St6s��mS��Cg�G��k�g'Nl�7��޲6��0:D�"F�/6b O�o�&�~ʥ?�^�s�y�C��y*�
�MQe~����z{���e7�����Pr��#��-g�ўW��e�K�*3v�M۰��L�{���=�v=��.�Ʒ$l63R�)���ϻ�$�9��9�����5^�����MS�s������7��A��ܜ]-�_�y��)|�YnF���ڰ�r`��{��)��O3�W�M�U4��&�څ�H��r�h�,�&���(��v���ԃ�pZކ�W�܌���ϧgo�a4�^��TPӚ�:��f��,��C�Y$�.�J�Q�O���D�N��'�F�\!�U��m��Z�p`�����5g�,Z��� ���t-%�k�r���u֐.g{�Z�5�\�^�\�oܕ.9��nlK~pf��C��Fd`�쐊�<��/��h``�B^������Ū��?���,
	�LO���Xv9�nxrr{s�����/�,\��W�32�nK"v�}����Pn,���5�Eē��C�c06�D"���/i/���#���8�3�3����R1'A�pe�;v��͂�XaϮ6I,�_�u�[}�ۉ;���ܧC�ٌ�����L�/��/�����X��2�	0S�*B K�o��s?i_IJ��rU�d�.�*����[#����{����ڥK��Y��Ã��嫔�����\_Q% U��w! +w��W4_~�w`������P�B� P�~$!�+�],�Ed� �#����� ��h�V W�}��?��C"0x|e�7�5/�#�    IDATL����!��z?W�P)�������{t�?�7ʕ�y���U�nz��	F���p�������/�}�z|muɱv�=[� �.�,��b�*x��:
,��I�y�Nӝ�)h*Oi8my�ۗ/�G�G�G��O�����������\�����<l�f��;_��^��n���ߌ.�2�p[k�1p�YF$���E�ms�b��<��"X8�T~��"��>�R�w.JZ�pV�o�c�p�.���U��!{�\�SH�e��@��뚠jA�`����3�����~�q���B�������������˿�Kˎ�~������]G��ge
�/~���/^�+�O���B�^_�.���#"zAf+ ��9�6�H�ǧ%��Z80C.H�)��`�"_�� @�Xs���Lę��F���G�����p�q�Ƌ�+�G��@�iu��ӄbz�?[_S�o����A_)_�h��4�V�<��u��ۅ�˩t�m�f�Ǘ��_��ޭ���Ҵ����Ңf�6^��2���i���)Cf}s#�yExJ�kG�s�A�1�
y���L4��I%����ĄV%���{ɍ>"s7@v�&t�_#�^SJ��h|��.�yΈ�MV����ӣ�Y��`�d/�<�� ���R�Q��N.�l�>�	�o_��]W��<���CL9d��H^N��|i����>�c8x�?��3��˼u��J��k� g���"B�Yʫ��i��\���)i�T�RU��/"�o�IE�_*�T���P����Q��I�p��p���FNbA
�/H�� y��S��	@BNB0���<��� 5"	�GE�����Kw���!��4۟����N���	�V��,���kh K=�B[8+w�S����s�睤��U��	T�*���J-H�Q^_���q�CBZ�+���'̖�0x$�3����*~�%�@���R)���MY���h��1*`�J���C��䇓))9�b}M�2bx��4��*�DJxP+��A��8���*�J�x��X�3X�EH���?���C���)��� 0�Q^3�dFZ�h4��W_}e\�JA`��K�Z$�#L��g��3n����x�K6>��#h%�:���B��K����/��E*�B"��B��0H��|e�# :Q�~�#'y�rhNN��:���ʨ(,9���K�/�RF%`����Y�#w!����n���
B?9h�a�*�H*$�B���ɸ���oNڊ*�
��0�by80 \�]^U�by`S�.���OɁUFj�pu!���)��/B� �O�ʅ	��2��ػ��O��\�rW��U�Hl��B�D�OE	�(�e��\mA'�x�$מe��[����I��Ԗ��v"���Θ!vw��}��g��غr��ɴ�ol� 4�8i�<���*F��ʫQkA ME�PK9h�<hЖ5����"(3�9I��Y& ��������W��ds۩YwY(��/9,��coyo��@@lL[��<h=q �}'�Mҏ�d!Ӫ}e�+�Z%��B����D�@<�͈g<�]{��5vuĆO�YY����l�����+�Ws�{����f^�~g;��j,/�j��(.l/��H>}�2$��.���`��RV�����/�&�E���O�g�H�/��ڳ'��w6�o�ͷ70ㆫ�s��5 o�4��8{ᚪ�r˓E6쏷ol��$��l"��s��Xh@���͗�T�K���Rkn��ˏ`�Һ�O�R�Pw�W3�CS=��.ԗ�C��'�V���٠c�ꃃ�����'�������?��t�ywv�P��V�A=L��TLV)��[��~���<"�@lG6�(��C哲����0[M�ܨ�ɣ۱�h�K���_�Nc�0�I����ek�A��aK�������m��w���D���@3u�(_�n��=���"'�,HI���x���8���.��ť����^n���O/Y�_�^��5os2�,���<z|���g��f݃��G�=���q�	P��A�<u������pc�|#��x���@ ܅()��t�B¬zo܌l��41��f|�*J/�q�Rԥ�~Er$%Nrd�"�@�t��~˲Gڞ�(��u ��y�r��ӗR~��T߰:�"S5~�Z�1�i�^�����Ǐ;�oȍ*d�ä!-����b��,����ߜ��{��bo��M߶���(�*�m	Qq����`�p ,Te��秴���Ң@�ɳ�;��U�͉��=��h_~ק���yi"v���00�hg|	�����L�A�����gW���8��>T��
Y �+J  ��B�FJu��j�E�(��_M篿{u~����+�+�:��Y:�	B`��3��6LW7���n9y4�_?zyu3�O-T�xX�IE0���t�1�A�,
|~r�Bl�W#��dE��V�a���{=�"��r�mv5��ۯ?:��̽VN�zD��c�&��%fm፧]|j�X��J������%C\o�^\�J\Q�~Q0�"	=[���%JR�f�z��<�����-��ΖC`�xs�G�m�%��w�?�g�s�x�զu����{y� �7��T�mǝ�1!03��B��E�U#��|�o��1�L�Yw!ff\����j["$�p�uD���*8���>���̮.�������ZM0&yg<�M���`Q�Vv1^�ϳ$���=�l*��h��;�kNz/	�F�FC�<95�W�X����%'o�:������/I/�)o��T�Ȑ�z�����?������xc����"�������{�L=i�_R��UCW�dhhC�AV��g�}��_j�()�K�)v�%���&gsv{��rM�
�]F�B�M<z�MџD�~k�W��r�����`+�������z6%s��l��o�D#U��m�B�&r�Ϣ�@Q:
.����V�L���9�{���tm�f�sݗ���d)��G#1��X-t��.���>��՛�Yɵb
�QѪ��L��.��4?����D�?~�1�V�
�n����'1��������z���{�l��H�	�'�����NO��^jڼ_6�(~4icH['7o�:��V�:O4Φ�#�Y:q�0�Վ;���J���Ud_�	�]��byDa�"7X��Fk�}IZ������t�Kp�}3_��n�a�r���z��
�*��0ȅxc/U�Ĩt�:;2Pf9>�C���i��@䡶�:jͩ�y�����]�a��-�ҝ���N�}k�:���b~�^GvM;:iǚ����Gd�$s�o!ہ�7!g�R�0o����ؘ�~��M)r�A���g,&+��V	�D]� �K%޽ft�]���KJ�RM:ӝ9MK�D�;[����D��w�`o��[&����ln;(|=	�a&�#�X�b_"���0�1P8G8e��������^�?B=i-��B��:-��u����>�α׉��7��ڳ�N�ak��'�aq]49`|���)�i5t9��^��Q^���]J���Y�X�-�����̷ٸ�B�Wzi��.'D��}E]�B8ᕫ*��N2z�r��1m��n��9]�7+�]&���rDx�0r����[�<HM@:��S#XJ�������
�@�]k��iA�ۯ�z�ɧ���br�֜���c�k`�Cވ!���t�^ƵtnSK�$����&�rGX13<��y?3SY,J p8\����?��~?��+���OĈ*�Z.<w�	 Ȼ$�/�JR�+�w��)��/� 9`�Ud����l3"�j����<�J�%Q���F;�[|x28:�d�C���}#���j:>3M���o����7�~��K#�E^)x'y����c��j�]o�hB�Ỉ�$]O��M�g�䙃N���h5c��\\���|����7���?�����~����G��l����.K����K���HB�;�����]�Q�Q2v8������mHˁ<�̸�H�B-z��\�`#��~�^�!VT $��GHU�>�*;�p�&��/�W8Oe'���)U��U���SCTY�ۿ���g�5!b����ɓ'�$���o���Y5��Yq�:AN�V4%�TM���`�����\w�>(p���/ �/'��q<�xLp�
w(G�1B�B�	��W�XT����q�*|��{��Kד�vF.�ڶ,F�Vw�pt|�:ؚl\Of�>XL�B��r�Fn ��J6�|�~2z̾�)떂��z{%РD�"��&͵��]�e�6q�xf�Ϙ���W_��ѕ��W����"3�٫�z�?ÜV��)�Zg�a7��M�ư]�C�%��̳����Vù�*�EDsj�{)�R�Y�UA�#7R�( Bq�nt���FT"ޛ^�5v`��n�W��ܬ;p�^���fo���9X�AG=�Ͷn�L�c�dʆ!��E4�,��Z\fSn>�>2�>p�z�rGϵ�㭩�v7���l�'�^><�ck�!��`(�� 	J���4몢��Q�*~+h�g�w�S�CRx|{3��.�@Q0��f �?�6��D�DW,O�C�\�o5��T�Y�@�	RZ�����<
�U8T� 89�E�p���HNZ�<��%�'�6(��p�����4gh�?~B!P!�1ZŁV8��J"-�~
��J�Q�<\y���+,�D	��F�ցE�F8H���v��/���2�(>!� �*���y��E����&�I�A��:D[�|�DQe`@RV���Ss��-�h��/�(l�U�W|d �x8��UJ��$08�:U4�(`���P�J�	r��Y7��UX�  �]�z�J
���95�a�rI��4����Bk��駟"=���NQ~b�)<ɕ]Ѡ�S����h����*��+z�HE�
D��������|u.B�*9Uo �3��)�E6<���UU��Ԧ��.Dգ/��J�UY����M��]�(��;J��+��VZ����	���!��Z?�fdH����҅�b9!��A�� L��V�������Ʒ D	[a ����`�`���ԪA!<b�q���՝��+hQR�嫌T ˡ0�ʋ1��|+�*B�'�+�������C���J�#Sia.��W,���U-��U)ۗvOt�َӮc �Ŋ�Y/�{��-�#�:q]OΦx�¨�f>�����L�C��F�>�l���a2B�(��J���'���|�$�RNS"�a����W�P��<8o��v�� �hٵ��S��S�6��Qeuk�Wg��9-D��ᢸ����ǋu�M��
aU
9rU4A�B�yW�B8E�W/��d(��q<�r��������-|	v��*M��e�w=��e-{�޻\��6v��������(�sH)�A�@�0��#C��)F�⑇��Y5��dF]T C!�A���ˀu���g�����Ǭ7v����U�4s�I�-���LY��-S�5�o����Ą�m��1H%�5�����FRE5n�h�_�<� 6W^�S*���a�����B��,x{�%!��<SF6�-�a������ǟ���������,�|������K�%���
A�`�N}
q%�؅������ѯPB4dW�@���'x�U�5n]�m�{[�_e���QlK�fy�=����d�'��v� ��/�s�F\���K&�j兘*PR
��+b�I�ȫ� \0��gꁤ=���k������hI?�	%�9�g7c�;ʸaZV;��S+{��W{����ag�ό�(�N@�=󧑁R��к }b8К'�@����a�B����c8�W*=�vQv���>�;1�rY��}��ۻ4#Q�ޡn/���Aykr�̀_�D�x�g����j{쎚�1�=#9��r�k,jy!�\��(0«"�V�B��Q*�� �n�\��cc{h�Y�p@r�E�4��6�6����sB����O?��ݛ����q���b���b��-!w��
A�6p��.p� ��'$��cIr%�^���\�#�װB�D�;4�b�`hVt}�����a�jlD�*m��rY��ҙ5C�ή���tr���w ���d$G�T�%	�O���Ev}�D�T���8��ae��ܸ:u�{l����e� "@U�lT��ӥo����K�7����/w潽��5���%`0Ï��p���E��lԲ��[����;����ˊ&����$,�B�pM !������DrvР�O�Qa��%��BL��l�l�	olϥ���ۯ`����񕛿�Ҹ��

He�Z�!��nZ :�)�,�v���P~R<��:�x�e+��f���paH��w�3��-�ˀ=�!�&mAz�tl�tq��P	�w���Q4�MƄ�]w�+d��<�uK�k$�o�u��0��f��+�7��<�5�����f�x��	E$!`�T)�����	�=:�����'�,(o�Ɠuw��5S �­>]���,
[�S ΄ƪ{:8x~m� ����e^{��X'/��;O�nH2�W��pbe��Zx �8�>cu��T���	��B�m���I����E�x���uVS:��kp!�w���t8�.D��s7���{�L��B@����y����t%��/�71�!98i�bL*V8jIx)򯍠U
�D�0{H��i�h��z�~ݡ��m~%>$�%�\ٗ �m꓋7g?\�g�4��d��kR��3�d���xx�L���F��Sq�����#\�gKOi\�����]>������ɇ#/���):c�8x�b��wT��
��!�{x�����t��Sr8�|�ދ��l�K_�q5#�(�U$acj�����t�)&�R��Q�NȤ5-}u,�B��W��(���>���9s�ҥg�..:��P.1�C©D[�/ίg��!�]��V��#bYs��5*H��rA�~�H?ƾ���?��Y��5�J��"���h6�'`5�Ex����p����{���_�\�w��t�K%�X��.ڵm�(;�xBP���`*�ou�4'�|%�R5"/<�rbM����]�|�?Z][�u�<��|���V`��i��F�4�4aҷ`�I��ZPcF�BFg6����	�.��Ć-rM��;�)8:qV~?6غQ���X_�+&�J�H���tۛ��A�x�7�:��,�~K1�{�w��Δgn��wy�r����7��d,=��D�LK��M�
�d�
 <}�Դ�7 �C���L�%����D�b*�.eq{3�I�q73���@o�]/���@�3�K�Z�yN~G�)��am�,&�oOu���]|�՜,X��P��Q�m#��G�r!I����90Ud_%5�#0C�.X)4}1iS7��32Cc��-��uV���Ǝ�n���R�Gw���q3nW�����b����ab��H�A��q=�"��%��9�L�)mR��'Q�b3>+���^��9���<�@��Hꇌ�n�~\-��sg��>����5�%tV3�J�Ǫ�nm�dlFES���#~E��u��[~����\�U4�����$~JU�A��?���(����O_?�#%M�R�|94HR�$�#��p&���VB"
����o��B������U���X�G��^rmu����Ao����?9���w]
��؇�^�˫7�_���o_;��͛��l�a�#�d��0���.lӱ��DEgh���l�O����É�E/ n�8�`� I�-�U����y�����׿����v?���>����z;�C�<�"��gb_��޼w������t:k�ںW3Pj��"�gv�'��؆T/ȨzI���g��Y�R|�/���19� WU�[*]H�N���E����S*�$LxI�)k�
����툍j��Ҧ×���;Z{�p�҃Jo��щ�ߖ�����	&�`��/��/� �U�bB�����sa�	���/�K�:���I�^���%|+��VEt�6�nK)���ʩ����^��@��[*H�D�I�
���7�n�{����6�:�7;��@G� �x��X�n�,�"/R�Í�,�W    IDAT�Qs�Q{��rteT��H�^.s%�f+l�p��U܎�:��_����7_|���;q���%ϵY*���ѩUX82��6��! ��F�3�6��Ɠ09f[!�	�t�H�>��5��eL�a���5;2+:d�3�b���ͱaM�B��,wE�4
m�����hy;XLs9F;)e��t�V�޽����-�t=ny#*k���D�y$E"�A�kR�r�	�f�����ehdbA����O�9��O;,�n���_�߫����������t�M���`nr�ȫ��X!�'���,Z��~����`�䁶�HB�d�'������VFb��⒯@ �N	eW�wQ~�ݷ�Yb_?l�
�
~_ɋH��
���`�S�����;�"�r&���4"��˯%jwzG	��bJ��R�y��(0�~�'$��!ėC	?0��G!R�*���G��WZ�G*����$��Ej�����=!V_!x�Y ,C
D��p]�.D6��b��>����V�B�A�i��@���KzJ��
�h�EI�(ߚ#C��r�Ԛ��PX��Nؔ�f�KeS�,*t�B���$:]Zm �m\#g�G	ʁ);�������	&S$�s� ����a`��J�ӧO���/^�@<��J�á ��<z
�t��Z�"�X����bJU`�b�����!
�*�N6� �r��N$�#P5�X����׌�`�P/��+�#��+m%�����g�{90�|� �"��]�XԢ��'l��*!��B
�p0�������#-z|+-�"X��B��+V���UhﾅM8"�����z��hX4 ���xe-D^��� � 9�@������c �%�@*�Ɖ�R�Vq�TA�c���2�I��2=u_�-:/�_��v6��;�lt��8Ag�'�1emu�Z�:\m'�Ƀ���ɗG�/�{}V��ۖ���$���Nq@Y��W� ӊ6_�
<�Ea�뚰Rk��� )&3�C�}-��'�s��Qo��; ��ۓޞ5����p�:��&���v��mܲ�b���]L�q����(����N@��O�����r� 	f`<XID��s��e���5sד�Ѣ����/\���r�����Z<a�mt>88vs�|йo�b�ׄ1����-rD�T_U}�`��>J4IT������W�RT��<��Ԉ�* �Bw3���ah�b2�诮Xr�T|�bҙ�g�ک��91������vo퀕���'׷=��7�T�ڶ�QH�ʯ�� B<�I�~����Uj~�Y�KαъTގq���1����;��d<"�mz;�o���G��=���/'����X���,�^O��ғ\f���	>��G<̀2LPQu'h�O ��.��j`DEr,���`�M�d��cvk���Y~H���w��B�u�x�G��2m�W/��И1b��b��������l��|�Ҥi$A�i�|o4������dZ��_l�߷�Ol/�������C���<K����1�37;?�8�����?�h��󋯯G�~g��%7��4Ijά�C.a�Q�#��6�gHHQ��O�#�ci�4002ρ$�*�_'��f�#�3��V�lf�À����MlakD���SETXm���Kv�+���3�q8��p�<�͹W8�S���V.�B��)y0���W,)./+?��T۸*�&����a�I��N4s��bc mԦ�!��v���l������W_}��m&�\�ꎯ�uh5��0���,O	��.=��oZ�@"U�
%���b��
h���Q��r�-�[�����gA�;�O/�DE��&���oI|�S`|u~s6�ڍ`�K�?���  ����(�$�GDA^uQ���/*�5�ñc6�m,>>ڏ��G�c!��)a�7��Ⱥ�?����'?��/�ק��F�w��h���g�m<��[�	�F9:E)��� �x.,X*�0>��`rf̌�/q��d{�c�C���膍v']eCp.�[?���Md~�k�6~8��iI���%����{o~8E�|#W�msE�@MLl�E�Q�K*�,x�v��ʆ��������������یmԗ��'�r��;���������;�zwy|i�v�vu=�i�F*d2�s_U����5�G	���N^�gh㰸:��`J{�Y��Ha�4��2H�L��R}�G�}]��7j�B�^_�o'�EP�1S!�H��]�e�s�
�vh���|���r�eD���Si���pɷ�&1�RҎɨ�S�,����y��!t��֖��^�<�\���E�d����3���<�Hă�\d׻�����?�ܹ�?~	ے��I�
)�%��9���l��ZK���	C���������j
�2L�%Z�Ll�j��d2�%�=���0s
S�>�L�ɬ��Z38�آG���fz���ly��V0�\�f��H^��/[?1�
�����-�k�E�#>lt�����Y�H�[˳�þ=�d� ؐZ���6g���SA��`����?ܽ<��u�p��0���E]Ys�-G4hhwʼ���}u�q�c<�a`U
�
R

r���� ��T�gY�a?{���`�ӝ8\MO#��&[��9,&y����W�q�g�ˑ1w#.�:-&H[ua)a{�$��h(z*��+t��jJ�g*�I>0�XՈ����4%���F�(�I
Ւm�G{�oE�ǳ�h;1B��v�KVYv[J�WD~P�~
��/z�}R��mP,G�>mA����Ď/.���l���C�����w�9ͯ�'�ڱ�����G�#X��q������iMyϮ^~�����=�$��nw�3��j��:����H5�R�#-<^%-V#[�}��I���Om2rZJ���d��Ct?׊�E�0�ծ�`��ڹ3���m�30s��h���Y�«��`�M���_a����I�ဩ��j��3��v��3l�C�Qx�#lX!JK�fQz+ceL�z�u����������Ʒ�+���G���� c���6=�b>]R.�`��W�$m�j0�1ޣ���Q��VE~r��V�\dm� X3�ڢc;���oJ�rcz�����>c �9���%9o����u�N(�n��]�[�̡́C��K�����`x��Q�������#u�J�|�5��U_�Zl{���f�/i�6��~I�}m5�EW�t��u"^�ݹ�;g~�SX3�D�T�G3��V7l�/[׳��aAְA��[ERܫ��Q�HB���F�/'J*?�
����pQ~V��JU8� �` �D*�R�Gl!�R�qU��-0ia��gy��r��_.�`+��	��םJ�HW c��X܎�[�o|x�|4������#G��^������?�����pf�����o�nJ�[Ə������Z+2����w��o�*!��򜝤��m# '>I������mӝ-�ӳ�9�����>����O=���ttς���.�R|�,د�̍��]\G9�g�iք>^��~h�0��-�걺H��U�(j�I�1=~��MB�����ϒd� ��� 0,�r�%���2Rw��Z���C�'@=�c� .������������_����V�5�+P�t���1�~򓟈�ة��)U:�Ү�jut�@��q�x����@��Y������X�A "DI"{QX)!���ޔA��r�p1��	m�D��Ժ�p�n��c����������OX��g[xm$G"�xy*��]2dL��$m75���h�q��~���$ �Dlt�r�ͫ�y�-l^���8�/Φ���x���N³	��D��@�ir]p�����Η�D��P���d�hi"���1ꉫ�#��GT&�M@�S]+��h��\$ߚRꉶ���&9g�)���]�Ղ�E�*S͚��s���z}c�Q[�_�o��۴*��dz�R�)tlL&M���
d�#S�6Z���e��}'6�aq���Q�l,{ލwl���B������O/�����ƞ��緳���l�B��Ȓ����O�n��)j���@0~*c�j,������ |���"��B�+��T�.Q��(�T Dq��[}Q��wt
�ӗ�K����ちh�V�����"������[�B @�[�H(P.��I+�2��0����V^Egᄤ0K�h�«�p$b�ċ���
I�J�/�
��b�p��Bz͐�)��B(#:6
�4�����D�b���OY�p��,#8����v�A�Cٙ"�IV*Z���q�E8i6J�>���Ͽ��K:����A��V%V�rhC$RˠD��5�,V$��nA!����W
š��EM�B�����N��N���-ߚ�/w�;��ڻ����"Y�D�F��&�I���Yd�i�t���d�EkΐFrzaw��� T���}�����&��G���M�'���B8���r��%L�P�|9e*�|aSv%��h p���V�`'H|��֭[�p��?�)^I'b�T�OV���Y*�Y@��	�������l���HQv
��p�*���'/LWF�D0�B��P�*y�7+���*.�a��*�RIR ��3A,����.����̬�@�NENT��LJ��*�V|��0��]��K�I"SQ`���!�C��B,c�V �tb��� ��$���D���!��� e.�%�����dF~J��36Q%��I�G�y@&I�$�Ki�?�+��0-~B�e^B��/ܘC�_����eUw>_�W��q35��^Ǜ雝�h�֚�ؙ�Xz�qe~q}��.=j�7c�k��A+?��4ك����xhMh0�������T/�VcW��I4@���Ђg�-�Xr��c�1wU���۝5�!Յ� R�)�[����͆��ГUU3����φ.��!	�~{�\u��/���X�g�˝����	pF��
wLX��O]��olu�Q���,�G�m�Fla��6
kO=0z��?�w�ۓՃŪ�#����Ц�7���1J����V!h�(Z��6��[��G������.��0JVKn�5vtz�h.^�]�8�&��fjdō��n���E;b�kWmd����qwH�[�Đ�rٷk���eY�Z�l\�ON
�A�(~��}����3�1(*��U5&���QlA#����A���	�W+���ٷ�~Q}5-��5&�eL\���~c�@���s���4�6�O��(?iW;����%�	�XS�)�ܤ2�de?�����V��n1G��!�JY�=Rh��V\�n���`�����r8e^[RO���B��BQ���� i�Xd )�KEq~���
��0>Q�1�sPBG�ʮ���,qDЩhSO,���\%�.��j\h�����x�����֯��ʒΩ{΋$�e�]${��S�E����1�* �x�Tg�)a*O4�@�����Fq}��-��ŕ\�[{����a����0�[Lt�� ��q}-�&r�}��7;;p�K?��}S=�!n��P������)��m� Q�ϊ��$0%�S��v�-L�����\������щo T�a�sf��l��y����}Y*�0�1מ1�!fT����ZHֻQ:�C���<����.]�|iɼTI*x�p;%�^ ��g����m:�xT5��VT���dɫdr�u�}�\O��k�8 �%���@n*�9S�i�km�Oz�"�0a�u�P\rL����W֢8\�2�rB"��
�O���-�[�v������F�ezKWU��e���w]RO��|��:{`��+ۭ���֨W98>��N҈H�r'�9�Q��=|���%�Ȫqi��H�86�:�a�Jq.��u�Բp�ʔ��y��2o��^����v�k���zj�o�+��c�S�f�k7s�ٹ���h�M.����~T��r�R�� !��		�<�T�}���Z�C�N�ˊ�c��7��f�U�Ey��<�e2]Ԩ�7�F,��n����{����������zԊ�8ǰ�ҋLu?1�C���S	�V#؅��|��ܒ]���4J��h����K��-O�l-T�($0+�<� JF|����ˣ�W����V׻�2�G�ш��bib�����=n2@���ӓ��3�j�[��PǴ��"/Y�WS�LYR�� (��DBD����!� �0M���Bha��Cu}sscY/T�Ua�uV#@ݪ�%i�VJ��ͽ�ɋ�|8a���3Z�[��3�,SdprL�A-�`�Lt	?��Ј��۷UxsC�n�)EKI�!-H`!��<Ѕ�S�d���ƅ��^#�vi�
T�[썏뱂�LrNs�� �ݍ�^�s^b@������2��U"v�b��,�9Y�
�g$���(���d���'�E���vL��v�Uf��ؾF�t"q<���v�p�q%Yq���$��Jj�:W�oݽ{����������
��N�`!�sa6OA��}ь���}��!��{�䓒�m�gUS��>�B���ɼ��Vmի��/J�ܽw��e�9�������R[p Nl�;�d���٘��0���w�����Cc�g��`�2�k�Qg �(��C1"^L26��R,��ʔ��o��	'o��~ǈ��8_ȸ��6��DXw��5]��F
E-�Xx�s���r�t�b��|�DoV?[�}`�d�f�(I�J��C$
�8���R}<~*�XH�~K*�M�C���ZkmuWG.Cq��F�r�0.�>��������5T�\�])�ޠ2�<;�*m+������FwӋ����%80'*ņ�Y ��WxV
R���p������̢�=���jl��*5W��f�X���Z�5��1�6s�y}��r0��L�=*r����%�i�EΑy<��:JQ�0���I8+k>n��,l�8�e7O%v-��v�u��U7���g�[��p\+�*��$x63�{�f�P��Ԇ���mˆ��������ʬN?Z�[m"�}P@A�2��sڲ�x����_�����b�_z�ݓ�����Z����ܼӐ1f�sϬަ6��;��m�Zx�������㓕�.
���l�\�Q���\�=��89�E�v��6�D*�  �U8��?VK�~&2!����T!� `8���Z���y�N�#���"�:�I�Ο����(�n�Y�"xB2p��y�-^�)3�_�rr�20�&������P%�)J)�
Q"?90~�  ��*�
���K�	���?LO���2/���T\�!�W�J�gp^�iX��Qvz5�ll\�[�ڮvZ+U�]��Xq��W/����7����_y�RhX��O}`�\;1?n1d��8݀`!1@(��(f�ǣ��DNY��VЫ��~�c�6�X�q�tŤ)�����]wM�n9�Ć�_>���o~չ~�ꇟܽskgw��Rَs���-Cu"n7Bm��j(Ա��G��u	�Mـ!Z!�*��.�d5��]<D]`V�9��09� d�I5"-lZ�(�D���L ��y�C"�O!����C��D隵m�C����1ij0��Z���r�*Y�M�@?Ƀn̗_~	��K���G?��Y��iE����gq-1"�d����8�='x�%� qrR0-��CN��t�J[�"! �l3<�y��%+I����N�屃V�VV߹��#G�
c�d�?�j��RbG�+D��g`<=3c	c��c�~b�<t��j���y)�w��H0���	�^��dp3Ͼ?x����hq�����%���!�T�rks��5]���?��������m%��U�*WҐ|��S���+ο<
b##G	FN�bg�;�L9�};֤(�Y+ d�ҧR�GE��2�<����%��|�L�P����X��-�%�%�V��_Y�gdΘ��	�74Y�F�Hk����2-��,f~n'�Z�~4<M��ƽ���wd���ӿ��z}Zg����� ����?)r�I^%ߒ���/<����ژۋ��'q��g�DQ��>�d���I�o�C	�uQZ
H���JE��#m���2!�9�V�)0�ό Ѹ�$    IDATI0d�)�p830��I��x�S  p� -�%6�#IBJ(6	L��D��_L��� 3M�蔗p_�rQX�[�nݹs�b�E��u�Q x ����QpC򃥴�?��?�*��@�I��z\�xnd2G,�$V8�ʅPq2b~��ݻw�E�� ���Ǥ �����s�*u Q�"O�����e�	s����C�q�� �DB�T(ڙ	�����C��M���f��	�NG�IHrF��@�$J�gV�b*��pfb �<�D�@=�S�����	�t<2�Ȑ�� ��D�V�)��m�j�*	�ZV����d#"�9�
�[�EV=^!*i��S�p���<Q�_e�<��@Z!���'O2��X�ct
��Rl&�6=��(  @߿f��E��~,�D�`��}\ZHJ�"�L�R'B`�$͒'~�D������`	��:)��$�'=�J	b�ğ��T !���+6�� p����&�DA�/JB�v�<%0�Ij�'r�B�Bi?0�3#�xцԜ�����vpr����V�[����D�n4�l㤡�������F�[��.����^<)��Z'l��X��"#^��/#��+V�b�R!��a��TQ$Y��L��O�h�����xĢY 1�7��:�,{����ܻ�*���B̬c1$��ŕ�,G���e6ߵ֪�<=s�D�Z���m����e��T (���D��ᶒ��	�Rg- ��Pb��✨��Fav��wF����g���-�@�Q~1A�����������w�W�,�'�%ߐ��r�Sv�����rH1���CI�w:��RtH���i�
�(!*����o5V�W1�j����7���Y��"gQ@
�>�F��`]\����mq��ry��Ag'�3u6[���m^�e'߉�0��V	l�<+�����1)�A�d5���u�}����ݻ�65��n��X��mk�7S'�a�7��K�&��_����������洽ݫX�m�l����+��B�(o�Tua��G@~*։�ށG�y(a& H�I u|(�/K�����*���r����]vf�8��JD��6xbpi�7L2�S8j|l��^�io�P�E�tw,��'(
~��Ț�A�8��i�~*#Y�M�|����	�)XYb,���D���ۍM���e��b�.L_Mb�!�X>�_��ӹ���Շ�_n,�Õ��^m�bS�eض4C�sR'`/&#����HJ�DHc�RŊ�8!�27yb5�l!.�l�#L�g+���MI\�z��O�mmZ�Z�����zÊ���(
O%�_(�(�=ON'�'KgŴ�XA7����N�}�r?�0���#^��M�3���������bc�E�J�`=��s��M�V�֎yP``�0ى��L5C��O+����Z��mm���\(m�\ �>��L�}e��1�!6
!��*L�:� 
��1,������<aJ;��Z+���i��E��5i�	Ӄ{��	Fy!%��HAb�F�+Sq�a�B�������ZT����$�8�C�%pE�5�8!Y�J�0	��<	�|.r��8��s�t��ɮu��3�
Q� �\ܴ�|s=��ܪ�1��*u/_��'w~w��h�>�|����(k�Wy����A�@?�XSEi�a0��[T���(U���^��WRĲ��b�\mnz�o{gg�}~7�P)��괵�%�82���M˕'$�J�m6��?\���h��1j�PD�5Tۄ��?ɓ��[Ο�J�	�qa����P���Y<tcI���>��]4J�5�8�I��2]���z��tH�C����7֮?�<8�n}օ��0|�J%��\%��EI�yHZ��#PE�g��ʖ�lշ�7t���k9@*�G�0��|V���4;��jZ�)�U˖�=<�{��j��H�ή`����D�t(?�3FbBgT�|�?�}��š{Q��^J����o��r�=�J�~�``
�X_� ��	��<�Q�I��ݬ�vH��~�^nQ����B
���W�6uԒb�L�_���_������L���;�X�T�$�aJ y�����B��L��:�+���e$�B�����	-D��PBH(9��T/����]u�Z�r����{^Rg�*�-g�Rb��LEW�9�'���M2+��SΎw�OF��4B9K"�C[$,x�����)��L΋��oHl���t������}���]r�:�aׅz����!�c���l�xJV�ʍ�ڵ޸����'��|5�&[^oP���z44 �Ѐ����(\6���sR3��79UA�z1$6ٟ!K�$�]o�7 ��ceT���ލ�{k��P������F$�3徟�_Ў���ǅ���h6�g`9�/�j�'c2Ž���8�(L!�m�ԍY�s�TV�j�]��ͯ����m���HΨ"֒Q����CP�	���p2�Y��C�&ؕ�i�dpDT]����d2�dA���Ǘ�y �:B����m�*��F��@FXT�6�yO�؇b^T��&�	����z�S����a�;�iYz}7�Ѐ!lңCb�s|rz����Q<S�hp���K���۵a��zN9I�����O��!X��D! ~!
K�n����w�8y���h��5�NmѮj�q�Hi��Ea ].z�ɚ��Xn��������'������x�xR��)N�:UD��¦'w�:���� '/~^�|�8'�1Q!�H�^��AO�d]��O�s����Z��vC���G6w������Jhb6]� #�k���Q�1��h�4�X_;�W�R��`��B�bU��I�@0G�D%{y$��
E��������+��N0�c���:.�6[ף�����2�x3Ό��a�O�s���~��ףA��Z 1�~�`?�~LK",�Sl�H0�@r�9�
�7'�V�|��(�t�K7�\ �B��y�R_��`=p3������.l�
�|����ߟ��0؅Hx�Bm�-Z������@�I��K��+CT
ǟh�B�x_�-�b�	�y	W���L"�0&%�"�"~�az���,�I:F���'I��|ID�T h���2T��aw�}i�{u���]Z6Z_�qp{\�O_?�?���<?|�=q�lۿn��ne<n�&�	ĕ�DMv8o��8Nf�c��fP�R�:�3n(��DQ�`�}Z�3��A_��cg3��a� ����N�r��Nz�GN�?��յ��|x���ݭ�Ku��r�1 G��]�?\��;��qzt6;��{
�d�\���3��Q;J�u0�$'y�s�o� ���TD���d�B`��9a�ȟx� Ȅ�V��ϷM�������m�ɝ~c7�r�ʣG�TV����}�������^.����Hk��۷5��PBck�_���{��L�(,�-�7{�����XN��;w���1C�F��Շ�D��,vIb���(����	@�@�@(��	�R6������
����.���۳V��`<]�R��ko��@�5�]s2���vmU�Ň7��7�RI�j���6�]=8���~���e������(����c�@�+"��袇%�$"Ɨȍ--�jh�`�0$�b�U�#=Q.�R�ߗ��=�2PxF��?�H��Ą�hu������4�&B�Mօ���%��b�5���X���X�7�j�����.�j�����̣M�֚~i��W�xm@#�U�#k#�!�Q�L��nti�f�P����F�袺q�ed�U�`�5�Jk�҅���������ZQG$!���}SB��y�%x��C5G-N�����U�<���o�M��$>��L����$I :�19C�!�S���Sq�Jlf�I��f�����s� ���r��O���@^Y4�7�p� �.k��]M�Ia��|"L��iN��(cy2;��Zrd+�$�" �pNr?��X(Ih.�(Ӭ�:%jH�X�����x��ϟ[�3��|8��p��4��r�8�	|��J�9�I��B�qp���g�(M�): P�UL~0P���"Yм����o]J�#C�Dє�򂐾���h0Œ�MÀ����"G����裏�"	�O5'%Y_���GJI�G�'�|�`����Ç D!@F���j
���+y�l|��w��nc/�9rb	F��^@-ï�@���>�L^)����Jr0��P@$	W��b"Uu�WH��~]L�N?���p*�ʂ_���*FH!�?'�XQ<��_H�F��R� �`?y8�\���G�$����s~�/!`�O_?���~�FFR���GNo[�y*2��Մ��E� ���y.RA��00Q��r}��pI���4�GT��Tl��	�93��� g�9W�H'D��r��W�$���ZB����.
I���0�ȸ��)��TG��|P�y���U��n#�BH·z�%�O[�'�z5�G���c�f�ؾ��%&'Ǧɲ��xH)����<&դW��������(!��V�kJ~>~�!Z.�F0G��}�F���jc�ƽ>����-W����H�)�u��<�'�!� :z�Eo<asj�����Gnh���8�b��od2f��{���*c��/�� .��ylp�m?��U�1��l��f��t�����Z���6p˂f���g��V����|����Ѥ�Τ���f���1���P��$��pU�ܹs��[ʖ��F����9䙄ru�j�!� t�.~��?z���F�e����{��ĽR��$㮐�W0���x:w��������:k6��)��(���!k��	E@ j��L?��)�`U�>	�L����ӈ�ɕ���mY�4;b�X`��C��	���j</`�S-_�x�2�Z�=�4����f̾����.�[<D��3�}S>ic�C3@@*��Ѳ��,H��@-B����*ԺW���n�^�~��v�=�؃U���E�XR��4>�$*˹��⸘�'�}���OOKݳ��%�h�8�2��U2e���'H�Q"�#�Glr[xck(WLjV�4�k3��'۽Vy�Y�v��� f�윩��	�Zl'��vu�'�>�G/��|1:�6����A�b+��@�zD�MS��Q�Ϣ��\��t"E�8��*T��R���u�N���lX�o�7�|���ۛk�O���g&��x�k$��=�ˈT���t��z���ˇ�O^ϚN�uʎ��E#��HR�<�&��t ���X~���� <��4@z�BI�8�3[�ZcJ�M���Y=��_��B����<��]��օw�v�����0Oc��˲=>�L2�dD I/�I�rb�Y(�8a;R�8�m��[�n�bY�9��ܙ�1�Qk����o]���R7��C��(�^�7�q�F9����������G�c������X��R�Z/��=(O
AO��M�Bfg1��
�dI�����$xf�?.fgSFY�ۖ���4X0ة���"��Z��q��Ī[��o����/��E�w���R���(���Z�K!��m���xE�<TJ�'��%
Tao*�r�e�*p"����{w.]ݫWǋY�]AJ	O�>���9ھ持q��������]�6�ٝ�{qG�ފ��#�8t�=~�"�_P����`R���ԝ�tq��<���jvz`8u��J��ŉ��'a�MNl(&8�t�OA6��޽;?z��o~u���4��!�ٳ���4k��ѽ��j$%m��<�z�{-� \J�=?��B�����X�*:�<����Ȝ�Y������_����mq���C�j$.Z�rEy4Bv"fs���P����������װ�-�����ZAd�~�<����yI �B��@
��W �I	�D�c�I��^�2�Z(v���]�:�e6�L_�!heڢ�K����K[�w���Vw^��N�q�!n�(��#'G~�r���g_�j�r�$�"�6���7Q����#����h�v������`�ڕ�k۞��&%�V�~|��hJ%�҈MxbP�0|7��fg.RE��6ݱ�Yl��{��c��C&���ԍ>W�p��P�~k%��ݽ����O^,������n�y�u��g�I���N�T��9����
�R\2���޽��;{����Ѭ��u���qрu`Щt��Z.JW,���>���� �Ϭ&4G�zOB0Bx��ʂ�zy�^6�Bo�(v�Fw�Y`��E�$./���6����(���#����ۇϿ~�r�n��91)ʞ�tI?���=�O6
�����VL���	%�$��;[k�QQ�j�ۀ^Z�G�Ks5��؛���E�q�����򳞻[A9�l_�	��B���*�(�>�ODb�X��C��I�,��L�Ϝq��U��e��:�	��냓/���w߹�Ҷ
�r®;-�}����R��*W,�v<c���?��NWV	����w�7w�<T*�qof1h@�H��a&����
�����SHE�����r����g�ϔ1Yln]p2��c>5:��7��C�N3o�+g����b�i�޼�����?z�+w��>�/����vf�T��+
��#���TNj�byD	�������UX¢6uF�-z130�{@��q��n��-Ϧ+�Z/ƺ�DC����T�L���Z1�����ã�����7]K�g.��M�jF��MQ�!�4o1Ȳ�9�Ќ!�����2���wvv7���SŚ�%�*��QJzyW���Ǥ���q���-�:�j�{���O�w��|zjWj��-1=��x����ȗ4����8�؅ȴ�p�DC
9	�� 	'�O_�K��,��֥�]!�����f�ƕ���.FM��:teeR�4ʠ��]7UL���c��6���W�n0zyi\�Tb�*
O�ɊFL���b��'�ќ~�L�+� �Ho���_ ��`E敁P�.UzR�J�A+�7��0��\ZN��e�d��M�y%�p��S`����vwug{��n�Sz��zkӑwb�>}����{�����OO��ekN��
ZL0YE�Y} .HM��vI�����]��o�'�:(^t�&����(/��a&U��c�E�b`V'r��f�B:ë�vZ�'=�?y��ū�<�{{����ݸ���]_q����ݡ������	Ų~Z?�@V=�Q,��l�,�Y�ߔ��?��'���l���Y5	�K�����$����!_�P	Oy�J�p��Z����h8j��$��0i�v
�sG�I������9�#VZM�Y��
+�lBB���9�5U��?�sV�O��
r�=r�-����-�8����+ e�K��LapdS$ɒ�5�lR�d��V8��I��9���qc��[�.]��i3�T�~hub~���ؕ�;sb��4 AAE�N�V�{��Hdkgi%'o���G�&#7.��&��(깄�����g�O��/�g��9���2����a�֝)K��d#n!�����{��2�༵��4� ��ȷ��'I|�e�޺�BƁ_|�Tuj4�``(U{��PQC�
�Ə�^bg�aM䦷�p�f��x5r�C���a�G=9�V�X��i.��nԊedo���m��D�g�0�N���S1�6;.ũ�0P �4Caz۫F��ʲUi�Z��/^�r�铽މ���N���
`�f��Y��=��˂�dI1 �$0�x;�&f~+P��B�lcِ�KH��ҢMTb��p0���y|�:��j9�f�B���io�2�Ҧ*ف����X�^��˲��#$gfʓ��Ó��� 2I�H�'<��D� �����E �i��TF� d.��2�0�(���R�")(Dr�	CI�B?ygB�������F��Kf~��z�dj)��͛�iJM�`$�|�JGIkͮ�%���kלRG�,>|hǇ$�(A���g�������C�ѳ��Bh���x����H�B�`��Ph�����.g�PbY��Y)��l�N���P�������!j��Se!I�� ��L X91Y�qLqN����ba�7y�g��Hy� ��`�!�"r%���,�*�G0�E=    IDATx��(��� <�F &duC��`�N��5G�+]��$)�J�����q�WA8!�ӟI�3�\��J8?R���7s	 �E���&*0?$`x�A�	//I���r�'ZY�!�T�	�#~�N	����e�Q
Q}�~�O�Y4�iq�7�x�P�9Jt|N�D�
>��Ė� �s��¯hR	�M0��������O`Hr�Wʃ�I &�dB��1Lu�J��|��ќ�b�b�xT�?x}ri}݃��Qy\���w<0V���/�óY�\�иz��/��������w���Ɩ��0�0Ź8����+-���~\��i�%�Й��e��B�,̉�
;Q�C�3�w���S�O]>�nu�ݭ�-��ݸ��}��qd�a����H��Ũ+�N/�;L�iTL{���'�hFֲ�X¢���Q1�A���$��C>gu�PH�L������f3!Á�;����.��R>�8ۨ�̲Fme�V���d�U&��f�j��ƍ����O��p���Q�q|���Ռ��ڨ:�D����Z�LD)R<pX,S˨��RA��I6%��M)�$��A�~�<|��?��������G�SL�,�V�����3�4"���\{��^?�=;����˶�Ϋ*���u��i-4�.ɐ)
D�҃�<Q"�h��#�'�{� �j�!3'_�~�ui�b�.�q��5��5k�2s�޷_o5�k7v~�������Y���^��\�׆n��AammW?����R�i_�&�Բp�x�ѡM�R(�j
�z(JXAh��Է�ٌ�l.�\�x��.Oַǃ��?��{q�:?]��*#��5Pw3�<�xUU�:v���Io|������J/UK�l���ҝ|F6��K��
9�����F���(�c�dH�%"<�硭�q�?�2
�X���֌4f�F�1�W�J�H���n��?���_��x0.V�OV�.�[�����#m�ny:Ar6�X=�[Ɍ!%�b>�8lD*O��t�ڂ�/<t���
0��\��6�r��n߿�ϴ��S"��n�*Z鏸c9NTgؿ���3��/��(:��ݜ$�bLx匍HE$&㭟ʅB����2J�� �x5��1C(l%��S,;-����:�u������4cK�IUL��{(������4�ٹ~�G���W���N_�|2ۅd2MxOԉۑ*��R�Ы
'�2�C)�܈.;Fh���
������1�N�"[[VH;������ڌ�z-�Ln3Gx����{����g��d���	v�|��0�1�8z<qpy2:#�ʹw��������k]GE�Tӆ�1W�4,����j����%#VqR�|A�OE�.�(��K�{G�VKE�ժY<��#����l�_�UYj��V�Y�����z��OϾ��n^}=*;Y�`�p0�n�-2�~�*S.�hCUf̓$҂��[1�!�I�X�\¸Q�6F����֊{́�����ˈ�[;Wnܽ����D�k�#4S�ֲ-��xaNQ� )r�~�������7a�C���x����=_TX��UYhV"0�8��ƌ��dxt����j��q�ߚf��h{��tc0�����MF(a����x�;j��+t���ϟLz�|)uGM'"�͎�i�ꄺ�<��pZ���ګ����(dq�!
QG�u���{���� �P\��B�b�D�£��C�+�h��_�u��/>io�/Kc;m���m}Hk�i�>n���tS*����؛b+����:n��<Q�\zQY!��r�F�$� ȏK����.F�!Qf�uK3���_�4x��H������$�&m ���~�A����/���t���ٿ��W�յ���jw���VFd?�(�|��؜}Pz�Q�Z @�*�B�aZ+��V�s��^+�&�����Nd����F}u8���7?~����PcD�p���^4���l�ZlV#���^�>k���uon����q��jZ8ԁ�l��C��5�I�D!�}q�TNK�p��p�R�yp�.6����V�[u�#��w�^��uՕ5�kJ1u�$��o� �	�f{�r����|���|��h�|�!�r���z\#ɬ5�>��J5�$��b�y1�a��#�&ÍX"mXZb��F�T�T��[mwh`�v+�b�ɲIs]�@4�,���o�|�w��2d9Y��j�Q�ѷ��ը�A�v��浃׏�<|e��S���G������8A��%��S��D��H#�A$ܩ*RHz�YŇI�/�>[w�R}3�v��*l�Tn�U)�Mw�,W���N�Vmu�:>p h0lP�g���]r{��f���!DE�)����!I``��(j5EE�����(ro����_�Քǽ��nB��~��|�v�65ʳ^�2����Z�k��/+� �9jeQ�J1�LG��Vn�t*�����JM%��.jz�BE�WB�� J�����)�y8�ʢP��S� �xȮ- G��M�/&N<a�4����ia�D�$����؍V}���{޺󫃾�â��V;�;�y<�f\�N �K�:AY��'8��X��Q�	��cob��2�
+���Q���X.5$ũ����ns}�Y��\��������EJ$�`��DKgQ��i:U?_�:zy6��E��Ӷ��uG�u�1j�>њ�T�F�$�ʂ��s���d���������-s��Wqr�:�MY,cSS-�ٌ*qݠ/L֡X�<��r%ƪF��f��{�������~������l5(�O~�X]��%��3�X��P��f����@���C��jѝڰ	�n��˭�˷nl^�!U��cwn|7<�����l�|�PìṜ6���؞2s��]F�[��f�^Fr�
Y�*<�P޺r�I� ��/0�<9�s�E���"LQ�QL��������W������#�C<IC"�#-<�R94� ��H8c$�u�c��@7�mt/o���4��vw�	������/������o��|��8��*�)$'�$���]fҋ�+�O��q��X�|3����b	%�����J&��`�L���-z��Q��RHHŹv�&���|����g���=tp���z���KT�gW�K�kk+��Zcu���18<�Z.-o���x�S��	��%���}1��dx�)�O!R�6Q�735���L�~r�0$��D�t)~jMp�	 i�ť헬
�|a���g`��o�����7�m�h�:�����ǩ ~eI�/	ϭ[�j���y@�������B��4�@���+o߾�Vl�0��"�}ʠ<�R!1=��Q��:�Ci�gWNy��h���E��Fw�l詨� N�����8��{�4T[,$�����4�ُ�8��.V�L��.����zN�˚��W��/{/N�Ǔ��`99���k�1M�V�HXL�$�
vP�<�L����YF�Ac֍�.	���%��"?�g��tB
���7i�f}I!���Pa#�����mL��QJ��T
[�4�)�n�I<e!�L�}ɘ�8ݖ���+XT3&5W<�^��(�!4t����l�-��b��k���be�>o�8�o\z���˳�XO?u�T����=q���0K�<�8?��9�g?�s�2�?���V�2bW����)<�$�@.=�~N���	�i&�I��3��׌a�vhd�`�O`T�)r�F���q��|!�M�,��@N.��&f!��.�?,�&J��\!��M@u�P`�b3���ʹ<�Y.��&�bh	��v_x`�x MDYn|��!l����(�G��g^�U75'hU ��ݻ6U ��o~��!�c�u5x�<�.��˗jc"1L��N��d���h�Y�+��2/+���H�XHx��&�)0���ի�*�l}�R�"�BT藯%I��\u(5n #���c+	0��"Rv�b�rU���PQj��`�����D�2���p��<a��҆��F���KqP�L�)$�#	Δ@ HRX,B-'\1���	ڛ7o�*�: �N���d���`�7�KST`�?<�xԵ��E��Q��R�  ��=�*5��Y���#-v),����'c����\�p�g�̺(��
X:0�f��}�(�~r<I�"IR���2|���Txf�I2���/Pl��!�?!�!��~�D�L.���D-��jI`ȯ$�����?�@�x ��<ɍL��8Yg$d��(a�#!~�MR����_ZDJ��)�
���8:���X�gǯ�;0,��e� ��Y��Y�rn�%ʵ�Jccn���ν_���o��[W^����mw7.]�rp���T�5��j^!���Uj���3��B%�� ���`��	��m���-�W��;��|����]���a\̥��2x�z�"�,����!��������ǯ�����bV��d�,�2
���e�Uk��T�9kM ��\���YQ)a��G�����p[U���Yݰ�u��@B��φ�ʸ�n5K�����_}�r���W�Aur6:��}�m,���D����<��0~E��6
��ࡊE��QN�7�q@��*��)��U�����j����K�/>sʥ�8-���,�i��(KLI�7s;^YV	���>�'�^{ɪ��\H̓��C��31��*ɐ5
q�7K�0��	 ���ω��
���+�X$��#`���h�w�}d.��h���h����0U툟��&{�y��kw^>�?����_M�c�Ng��nk3p:D��<ɚN�59�3I�;��Q���: �a�46���B��Go �Y�;�����T�v��Z�YN��L��$qu/V�^�.�Ib�oq|���l�Άg��j�����ISJHv�#2��ʴ<���`�L��	���oD&�7Kt[���s��0�8U�{���4���
���P�3`�:׫������/����a���h�ǋ>dþ��*���_k4[��+���$I�ͺȲ(0�m��<]�VP�6'�*ϭ�3%{6>��?��S���ЮrL��4��K�B���d���rY��h�O��c۝ˇ���,N�O��⹣����=�d/N������(��Exqq?gp1�%��xtvr���;���c��� �����:s���k��!��4;�;?��/<�7�>m�y�KjF��1��;X�'��NF�o�����B'
�Z큍A�Ѵ�����qZs�8&��59��:,jƱ�ŴS�u;��n\�~�j{�]�V#�Tb:�Iȣ���)�Q�&b�,�,G�����Qc��i�9���ƉR��9Jx�T����&{���3��(N!����Wr�oTw�ء;�����0��@Qٶ���ą:&w�-�F�T�n�bu�Ng��x��6ʍ�q
��w:td�Mog����HJ|�=<�ϳh؎#@Q�G����y��ґm+U�ͨ�����b8[��Wk��[����y���K���MD�5ե�5^�O1��XEMG�Ў�D=9���k�rA��f
�á�/���-�)�s��Q�����"��wVe�/S��W/��.lv;[��� �a*Nd�!<�w�ڷi�QۼVYm\���_����֨��T=��7z6Oφ&�rT-��K�,�X�#���IDI)!�O
�T�!
���;=Ӥ�D�+��ʥ����l��X�U�;?��w�9�F��e�T��P9��#t�!޼V��XPp�o�B���+����3>�}�!�3�<�)BD���3ً���  �9�,��-���!�W����|]��H�
3d�k���Z��m�j�n����>��j�dyq|6�c���"�t��V���`��$ ���P���`����I�P8�
�[��)ƙ�e�~��?���~aS{dHqͫ	��0�P��)~����O2�0>��������i���=5�*���F��Ӳ��?��6�`T�£�J��Dx8�$�
pVSxTr��'S��N�Ŏ����]�������l����St.E/�!���p1N:��E}�r���?���Ç��g{��Jk����ς��K;H3�4��:�D�٥y���!�֐��Z���	���4۵��^b�&PX�	�g��ճ����a��y��d}�ֻ�߇! �S�#�{$�[��r>��f�;r��d�1uM�W/O�#�L+�8Q(�΢m��4$��U��E6�ˡ���
�Ph_<�j�����c�}�I�(�l� ���=� C�!36=$Ű�徱�y����io���Y�
��vXK�#���d�ɈD�./3��'E�bу��	9G�x���Bt��U�w@N^f�E�kگ:�v��?����R�S���/�):�����j+�l1rԪ�Zq_ %m���غg>h�R����&{��o�8��)���	+D,�}9	E	����:ڥĿ~m��ƨ���]���@K��Z�L�Ҧңuh���\\ں��On=��Ѿ���&c��V�Fi�����Ea�Ɏ�}�d �d� ^,nKi_��	�S_F�5vi/��ر{4�ĩ���I9Ez����������0n$]Y���~��|'�X*ex�+���&ߝ.�ܕn�
�l�4m!��7��¥��"�Y$!y�B�F�oX�k�V����fGǯ�'-l��`.��a�܌w�7��U�Ͷ;��پq�_�軕�W/����1��lE͂'�Z$\X�����4�@r��HB�?M�U�����V)!�=@h@j���DSz�W�[;�Oݷ4�׶ow�}v��\/�]��z6q>֘��B���5��Ȕ>��m����^� ��a9�S��aY�d8��E-�(T��>�������
T5$*!a�,ң��` #�[�0̙�(�_�"&��8$��L(&�$O¤IYY���b#R�tB&K^\�Z�씺;��h����W?������������tJiƷ�>d�;�r����J�WB@f�s�����-��ޘ�����u���ȥ���Pio��'�b��#.�Ȟ������]}}vz6~����N?����z�f���n��k+u;h=Qa���A�7�j"�me��-/&��U������ P�y8���ee`��A�[>�^R4I ��������K�+%��T��(ȉ�/�����h` ��׿f��Di���`�2H�(�y��7Hd*�x��@8��R�֬HO��
��۷og��{e�HB?��@�$K`y(��!�?ّœ��b���6�R^	��e`g�Ѭ	{ރ��n�xw�^�Y�]M��i�!*ö�b�77'� dA�OYf��(Ԃ����1�7I�`0:"`�>�zt{�Z����3�/�d\��f������І��F��!��hR��XRpTv��h�
.Ӭ9~�&�UQ B���?��	����ňr�_�¸��6�����4+�ı�.����:`v.�&ඤ�C\#c�G�����4]�jiI�a�7[�Vd���(�V��&�e�g���P*�ʪ�U5�}�*Z9+϶�n���K���6��U�I�ӛ���4�����.9ᔗ���2`A�%O�O�qb�����3���'�g�:�~3�z�%���x�s���e^~&�?s�r`H&����B'6�KTJ���� ���0t�Q�M�� �&�y��grI O"L�I0 �����
�����'���$Z�  �(���xR�Q&�#퇰(�Ǐ�������r�\��g�EC'��QUF�V�d���o  �K�i�w�}��7�|c�P�(-Ƞ���i@q�PZ���d-P*���Pֆ� �D
맥j�_��B�P� c)��I7oޔ0��R�9HR p�L�J2+�v��L�[�J.
� ���V��
�,SԂϚU3:`
�pi�!A����e�a�<��!��2�,��d�v�ܹ��FH,�?��Ð��)6kO�C����O�b ��+vA"��*Kv<`P��Q.'���~B@����Yv�` �d$G]���O��?99& T��;�p~��M    IDAT�FT"��0�E��%I:����G����a�,�L�~"@<�gF~
#��$[13!��� ��J�y�6s�X� ^*����TI Ȕ���'�H>��I	��Q��?�(ɴr	�RT��M @f�*��L�� �=��$	H�.
��A	��	M(m�6L����Ɍ�ǽk����bh��Ϝ-��Za�o�%�c�¸�XY��d����_�����k=���ƺq&�ڋ�d����F�*NS�4��D�G��Oe�G]PD��	^B!�$��[5�u�º��}�`���~�����ڲ4b�v�Rl�]�m�ir
D_��e���w�������f��`�\���1�uIY2-x,Mf���љ�EUJ���ȴbg�G�1��V���ĩ��v�ppR�[np5� )@ֿ�@�d�RI�%�������楽Fg���w_=Y�n�x8��r�q��컱픒��֗� �`�0I-��5�B$�P��J.�� `5u��ިC��`v�ee��{���ݬze|vV���T]P�|C����l��^$:q��Á�V&�'/O���y�Ie�Z�<��AXQYk
1@0��ik�R���LR��Y��ԝ��
X* �,JxV�8�M���������n3č�j��͵�{J鍝�[���s�y�ۿ��,%7[��͞g��zȠ+d�H�eJ��t�Z���=�#��jev,�,�R$@Jn7 Cjah�;K-"���������_�i��--����]�a~*z��نZ#ڎ�9���hԪ$�ޫS{�_W��c,���U�t���A��S���[�@Q`�2<�fr�?y�H�Q�HvM
c�dF���e
��ǪO�x���aZ]Fە�w��.���/��O߿~1l�-W5QGO;#���A��d�Z�b���"��)a@�R��oTq��Ø#ː�%�y�����������O?��?�����V&�M�h�q��鷂�-Th���_0��C��Y�]_�{E�by����]�Y��F�[��p�x��<Y��~
�.�a��IE�x+U�����jg�;\�٧t��q�PW[c+��3L�L�.�]�.Uo��{�ӯ������W}�e�٣Kd�L.�?\k{�1��h�#�@?����8�8)ۢ�h�J+�����7��prU��5�ig����ܹt����mm��J[,��,��e�䘝��FjT6r[N�Q5[�������F<n��*��?�a(�p!�8��$'�WL���V'B_0�`c	�>��_��^�i�ƳVyѶHuĒ����Y���*�n8�h��Ə>���ۛ������ZZ���n�no�O�O��,�?�?����@��d���!�J��!=�,(D'�-�0�EA\�
����9�Ҝ:k��._i�\���;�۫�v$iVz��k�
�H�,�45H�aF��1��{�&'�amA�%�q�c�l�'+�">�Of�V^_���?6^k_�;Lܘ[���p��Ž��Ǌ�}�?�
c�����5�k��7�Jޙ�|w�������2n�O�l�1���%vHF&xk�@,sx�B�����m��lWAH��:*K���$w���r`���F&�.����Z���y�ɼꠏq#	��."w�6�χqD�Ϸ�8���%	�hQ��8���@�@E��<��3� �����9��'������!�xڲ�Zi��=�b0s[o�`���>��˗����'�^���~o�Y�S��m}�gRpưA�<��#kTe]��dY�Y8�8!D�O=)"3ф�k��ر�:�T��Y�4l�[�vͬ_�y����V˖���(MFN*�J��>F�.�S���ܚ?�j�[��x2���
tP��"��t�J�����"s��\Y4`Y��0ᴕz���U�7��S��`Ȋ�8��f�"���GBk��uc~H��n�)������w��w����|���z|J\��3ww�-�Qi��]
��� ���B�3y�^��p��Zii!C#AZ��TY�UsYrdZ���D�mͱ���K��ɏ�����A;OJ���ߋMB1����
���+^��h' ���W�O�����r�͘?�S�D�Ix��p�"�8��g7dN��(	^AR~�W*��&_MÀ�w��Ȱ{:m���V<�U�q�q1��e��ptJk�nQ�ݾ}���wG��9�uK����fc�be��P����5dG3� �T�ʕ+hC���Մ��$dv��ی�;E8?9���\3�v��������^gc3���P�j�r�?�A�8���	^P�.�����H�5~
S�ux�P��x���9Ñ���S��&�X��B�W�2�o�d#�vP*�x��8CQ7�U�zǸ(������Uˎߑ�7jvgY�]vo�����������,���hk�z臸�'�ݠC��%�0%PYb�Xf�''�S)	o�b�rT�KRr�m1���W��C����_�du�e���5�sc�X�d��%�#�:tAL��qlI��mv|�l�^Y@l��|��h���]�t�0�Q���A6��?=Ec+�NT��_Z�k#�o�ꦀ��xhc�jg�k�L+��(6ƙW��P�i�%��]�T�vWv�޺��/<�ܵr��;�K�уd�R7l�-��9�^2�����bA�񡆖0�9�y� =qZ�ٮW�E=;95��i�n^�������މmU���x0�[�p��C%���2��;�
�<�.���L�9w��3�xc$A���b8?�S��?y������!PI�h��+�HY8 p����`0)��K��(?��f�
u�Y$�b�TEv	�+V8H����	L@�/I1D�}�����#�v.vw/l���'�����������SC�Cx/�&�H2d0��eAȩo�ȍ���7Ժ�v(:���K�"�3�`.�Z�Wx�L0_8�t�JYp�D���j���h�1��~��d��a5XĆp�f�T?��O���t�ݻk���m���r\b~�� ���Пn����?���)�~d��D�d���L?:�MV��(!���!������=˛QPe� !�/`�))Il�F�jI�^C]khFA6$}��.S��iW'�$յ��͛7=|�9���#��Ň��* ��SJ�׾��9Ag@#thՙ�23y+��A~�F�m#���C��d	%��x��d�������2�y+��p�k�q���^�\�,�ˡ�n͘(潶z��֎W���QHR�1Z��,�1c)D2��Yx�k�5�.1u�{ԛ��#S��ыg'�_����S�s�4c:�6�oR���t"?�JA���6��ȱpYv?y�%�)^8�#6�3�i	�H�%d� ƟlL ?m��
-2�b.��F�����<��_�p1xw[�6�fQDa��6�OJ&\��O1)F�vN�Wu̶`2Xv�8q226i�0TY�b�pAR̅=��_�̝��Ɖ���Y�ZX+��Fg������w�=�j�Ӷ�*u�09�����C��s��_F�E�<2a�uBU

���L��
|����@��g&$�JVJ��yZ!� �/� |SS �H���S,�\��	C����sH����hzH3jQl�%�*!����$U aCCf!�$I r�  E	�Ɍ���X�?1KB7%�b��,��/-M�ZG���\D	�V�!2:�`���TZ#	����$����+Z�j�<`&�Z0EDk�����Sd�a4�ܕș������?���ݻ�~�+t�)Gc��^���J%��XyA�B��J����6�K� �1�@"�W) �sx����|k��:��O�0;K�R<x ��і�"�����Q,�rhC�p��L���]X$/������1T?�� ��(%&����'~�� P�����7�(�$"9�c�
���`�A-�`@��\��_�Rk���e n�Pd$N� ���9e�D�RG�b¦:2�G94�r �EB�j?C���+�XI�G�ّ
�q�O�b%���!TF�
���V �<X!$ᅜc�@Y'f�����q����琢�T�BMeI+��9!(�*	K>��;�,ñ�$����;�{I�~���bq�\��ݗ�������ؚ�`ـ�?� �9��0��'ۀ��{FR��V��-�4��g�n$/yI�^u�SU��� J�扌������3��7��Lї$��?SL |�I�d śt !���s�|�L8N8?!cI(x�����nXn��^*�Y����������e�L�g`S�1�X��)A� ���>�v���Ʉ;�|����/��7&������KG���е�{�`kǮ�YLS2Tș_��C�P�7A������Ȕy6����v;͵�ld���"�����ￌ�Η��.�p���+�^Ҳ\���"��	^�.MF����^�f��Z�{���N��������f�xz���39�,>D�("/��G�~��T]�6�������jq���g��.��r�h��n���������?������C�6�_d����Z�c��"I�2��C��\2���@��T�q}9h�'�F����l�[m;�V���ն/_�7j\��/&C��.��ҭ�F����3W��� �͜�=��˽G�+�D������_�sV��j8Nt�%�TZ��&9��|	ʯ|���e6�44�S����#�����7w���Un9I��5yg5Mc�L),��]��9��>���ΕW�_]:9^���F��Fi�6c���A�ݣ�dN�Y�t�_��a~��s
ÎD��`�=J�Da�b�؜5�',���y��Wo�v��:wq���Y\�[j��Ĺ�+��cn��������rt�q~MV�f-0�+��2$��R��h���/!�	�ƚ��'�]Y��G������||rr�si�j��D���� f��>Ŏ��i<gt����G/���4�n~���W{'��um��Q�j0Q*���VdFg.�).Ge.X	"M�M&F�U@���5I�z����n&,v�ؐi��M^���ݕ���z��M����Ҵo��OK(�2�7(�(Y��0�j��tqv<t������3�=�IL$��բ��ybI�Ӕa�OG��K<x y�L��C�E�r�d�\����j�ǃ��h�3Y)�cV+F�؍E�-�&����|ظ�L��n����?���������V�&��9qH�1���f�4p��o��O����#����m���zv�I�u�s�7t��Y3M���O�n���Ѽt��ݎ�Z�ø䍄�"��hU]���7�C�Ȅ���������6ТE��� M���i��H�許�l��O��)Xh���X�<ṕơ�FsfE�����\�Z)�]�^�CQ���� 6��Z���nu��՗�W���ś�ˋ��g�k��j�����I�����,#��F��S�=�dO"<x�k�4ݢ�k�ϱ:������q�lj����qg����x�՗K��/N��Gg��*izi�,�ٍ�Tj���f:��?|����4�j6a�R�!u.�)4_Z�,�Qm�܉(�����U�㺿�t������X��Cr��Q�������ٮ�~H~���y��F��߿���V����dK�QQ��C���֢�qrptH�k+�8a��u���<��b��1l�/��;�r���,��9>�ߨκ�Du{������\.�U[3&��"Qَ�E�v�?�{��I46���t�ppr�7wn�@Jn��Bz�D��-f@�`�a�a>��+)���j�ɊhRAP�N1����m�gM%`HԈ0SŮ�X\�g�3�s6����~p���w���:���8I�HK9ŧ�_�����ӣ��eG�tLLg�~f�D�2��>��Ő)�Zil�����'?��o��K�oч�b)���J!�e�zh�mɄ�-�U+������ހ����zE;j���2�?�H&eNup��'�ª/�|A�rIO�Y���DWw}�W��c��Xn<:�=8�t���J�q�i�y�vĘ ����>�qϧ��b�s���O?y�/���Ѥq����|r:�F�+mu����� �ĳ�!��X2)�1Z<����ܹ��(�̋���4��s��\c�u��;/ٍ����ٸI�����d�� �Q\�Y8Md�V��G\��:%Ӂm
���5{h,�������脆1~tD��&ik���O�~��3�f}���>ӽ�����P�AOb�L����<jh�U\�y�c}��˟�W���vx���vz��V6�Y�"�3��B���!<!�����}�?ك���tb����������ʤ��^����+������^y����B���=vjlL�Иs���F;g_����������ܖSgkj��hϦ.�aO�I{!�btI�4~�6R���8��ŭ<.�2��%�h�aܻ�ծջ����)M����l{�Ҟx���NK�����H:�����wۿ��W�/�\�o��|6�O�'��6D!-b�`�@�ɐS��������am�� r���A��b��D�Dw1��J�U[�t����;o�]*�#;*�N�G�pa�RU�X�g֣��t��1X�f�?�|aGά5�y����q)r]��c":���6ͻ�GZ����~_qՊXVU#��`Q�Tc�T����M�PS�0O���Jn��I�G)鮆�TW�>�]�s��o�+��a\<aw65 rH)R$7de�f��
'�n�i'��˪E�/�4̑����:���ڶIVr���.].7���z��7_x�53�sw��l�w,�MwJwLD�Wd��:��~�{0|�hw8�Fv��̲�O�~r<K�xc=�B�)�%xb�.A~B���Y��E��	�@8���$�aI�?c-�⁏�e�~B�5A�3R��E�{ʶ�3X؟0e�:���Z�ҕ��v����f�69���������_}}�I߽[U ��qM�:j�C��Y'!�d)3�~��q*?*�/�DN����r�$���\$8��_��1Z�i��z4$�
tFsJ��R��(v��l��m�D��W��7O�N�w_���"��cT�����V�b2��uܟ�\�]��W4�c+�ƅ��]�0x��ņ�"W�i�9s�,q?�E���g!�g"B���Na|e\�AN:<E`�aR ����;8�L�id�o
:�)���ZI=�����o��2Yup�X��&Ֆ_O�I*S�\ėC�,YI}\)�����L2ڭw�}W��'p��EL1IUXIA��3�	�R-|e�(`K)�A	�̺�e,�7�^������:b�b�Rlաo��S$Э�4�r��G/#v�ǴȳV�� �}$ᱦ���C�<����������x���d�hv���& �?��OFG)I�p�����42(�6dA�26�̯�%<�<3�,�%$�)[\h�OL�t��i�s�	I�/�¯B�U�ol?D-��!�	Ɗ�<��PH�bS �SΆ�����4�K�n�_ ����̋���+�b�Aѿ����ϱ��x�7vC`"�2)�D��Ȥ�d:������Y�v��+ߍ���݊+ 4��M�yI�I�~�KQ�K-!�� ߔF�����!�˥<��+?U-�
��5-���
�}E�2mWM2_���� ţ9����!�M�e��<SE�T�"ȓ���3�P�q%E4}E�A � �(�B!A�A�{�P�L>}Q�X釉l&$b��8�x|�Bf|%�'4��f`�F�-�����#�f�c[��׮��ŏ&j�컮��<?"�� ����,����e�l�0?�~��}���v��K/�dM���L�D�i�0eW��)�c� ��ɰ/�@�_�.i�����Q��y��!4y���\s�����o�mm��$me���jR��7?R���%�>�弃�ȁ�@P�)~�D-�T�DɸF�e����/��2RX�,���V�������� ��E,f_�������_h0 Ҕ@��I���
Q@x�ȚF�Z2 d���+�
P)��D�y	qp��BA_Ĥ�+!�Y���� �g�""����ŗC��J��K�s)p�~�C�A�˟(�$π��DP�,�H.1�Q�L&�k�e�    IDAT�c�����$ ����q	�I����'��d	W����D��!(R��P���M�$"�P?��ɡ���%?8�ɏa�|��`�JDr�<�sx
?=���}S8`�֠����q��{�t��Gg˷�7���hF��02.�m�ѻ<�?>.��$.��h^o����δ�����J��99Ѩ��'3�{��x�E��PZ��s�������#AzVXU�R3��nf�:�g;�L)�M�{/�����]�1��ȣ2��3�M���w��/GE����4�)+ٲxp��G�bw�Mv�J��,Y.��,�I���%4˂������:�ʜ��A��$n#���:��}l��ؗ��[��/Q�*̙��iy�~�q����j�䬴1�I�JӫA�Mn�V�xf�����,�'���6`�J©�6���b�:c�ĵ��x0��iu՞u�ޛ�q�żz���nc�z�bU��p������k��<y�m�_�{�T+��C�l��F_��8���ɓ�&�[B|I��ee��K�C�AsS�TuL��Y����+,��z�f]l���W,�ؿ�p����]����I�׬�\����G�Mw�_}y��>��\���h>��Z��D3��Ql��4&9c����f��6d@�$2!c�ex�@4X$�#�s~�x�+7��������%�a�'W���X �SL4ʚ�E��ųab����xx��x�{�,u�aE��Z9�o��$?��!�%�	_v����Q���3qa>�ӎ[�7�ǻ��������0�`���<�rE[�u��#�g�ѩ�N�v�yڶU�x덿�Ӎ�zr���o�FJ��KKB'.�O��;��=+V�K�7D�
@򾲶T���ؖ)g��ɼ�e6o�vj�:0����;�|��.���!��ᮁ@���Ӈ7��g��k?7g3r���dt<�}���ƴ��1W�*'�gʹ0�N	c 3r$��oV��p��̈��N�"_�.���,ĖmS�������Vkvsĭ.1��_�9c(��v�x�Z�R���k/���{�_�f
��������+{��q�t	�Ʋ�R�W4���C�M���q�mt�L�gcK��~g%�>���ɭ+[����p��}��?`(�/�j.ř�������Ise�/[
�pM������v��&$�������e�pd�I����' 2O����y���D$a�8� _� �9�=$���E�t.zݎ"�V�`�	͍���je�̬钃�����}�şN�{���7��rd��uܡ�ϻHI�xy��d��<���S>iÄ&�,L�˝4��a�.��6�k^LX۾v��w��W(�WԊy<�
��?f�A&s[f�s���$�yN���۵�߅����T��RT�x���!=�)d�\���� YD@Q�ß8D�pX�mc�͂���ho��625Zkq:W��̕u?��ä�P�gZ�K��b���Wo�9?=������Z�S���G�:Sup������-��E��-i2�I��WK�PN.�-Ԝ/V�\&���Z�{�=������*��a��?��)�k��vU1��c�1�s�Ş�����Ⱦ2�-Az(!<@�ғ�O��-%@�C��K|?�_q�q��픻���8�m�M�����D�8j	����A�b�>!�*�j�Um�s�������_���z˲���9��܍�p�����JŒ�i�/ny�Oh�q�[b\�h��K�|���jɣ��]�XY�t㣟���K�FÜ�Ǒ�MB�q Ӡ��KSv�>C�#�ΒR==8�w߽�Fg���G���v�@�V��<c&%��Pr�?���2
�������5�Q�V�F����ڝ���|R�?Xou��y�X͑ig���R/�Ѝ�v��z���r�J��������ݿ��tu8=am�huYV)FB��Wc��%�����9�0���n����xI�O� �j��<DP�{z���^����R���S�esO�Ӆ��6z�Y)'��T�(9���n�&�Yߊ��k�V��ԹL����p����$��@NQ�.�+�������{��@�ś�3�_(����@j�X��h&�� G��V�^4/W{�߹v:��ųJ%�ު�W���H+ӥ�Ά$WrA��Oȓ��s�dr#a8YY�N�����j��k�;�ժG�o6.m����J]g��=���t�6�8�v&L��*���E�],B�F�`��7�G��aJeS	��8���\BH W�� d�z,e��<��/�� Ţ�N���h[�8�>��6:�"co{oXB�����}$ǖ���9������㣓����כ�����t>Yw���疁0�G*�0Vc8W�^��1��%�=I�P��&p���F��B=��L���Ԥ�+��|���*�x�Y��;�l��N�Q��z�P�������g+�c���;�۟���A0��֊4�$]L2��Y��VEv��X�|�C9"g�̠�m�̔/�˱m��=ڀ�/װ��z��Ͷ��j�j����������!�e	c�\���V���+���Ov������#2��}u�D_
W6_����Y7��Q&&�Ψq��.�)|Q ��c�.��Y���j֮l\��ҭw�S�^�����ٻTm���=)6'�b��E@VXu�fco�Y�r�G����CY/u K��Mu��U�MI
�;9pt��B��爠����H�r��Y~�I��CB�"�CA.�~��u
NJL�q	ɸ��.���$L�
��D�V�BU>�ڍ��ƥK�KW7/]�j�f��'����g��/<�2�,<����j��h#�P���1:&;��h;�5e�rN��fNy�Uh\BxR�Y���Q&�R��l�-�眗��� E���=��}�dpҞej2���[�l޸����a�j�__h�i�kO��$l�rφ�N��0z�5�B�il�jYj>&a��I>3%
�J�
ৈ�R8�IG��x��@E�����
���
�!f�R�1��{�a��?�3�b2TH?*���x���U�8���j8:&��Z�.b0a��XA����޽{�$�̀�{߳a��̛�e�}1-.:�[~8��_(���̟�ǵ;�%��Y�~Ֆ��*���hx�x߬iv��Űf��s�&+vpP�h��eѢE/���J��X�x�a���ɩ��O�>�K�C�����i��Ey�A�yJ$t]5������'�������#�	H�.ˉ ��ʔ����/��D2
|�j)�Gf���X�]ݬgX�����=v"j)4�Bc8�L�?Z���I��r{�S`��h��Qߊ��=�h����Κ�6�!%��6�(B�$d��B���[0�F���=<�r-N����κ#�k�Y�+8�<�jr2O[8��ߖF�x|��%�"�a�9~�ğt�2��Q�8?�4����T�D�Iʾ"J��C�pD"ɂ�e��^����E)V2cA �����lB˚	~:�f��~��7�K� �2]A�$���5܂�r~&�t;�%3����P%�(bG��q��&�IT�Ba�e��:Kb�1���A6g���-����lm	5+�U1�HHe��/-��c.�����C+j�,�o�a8*.']@h)|YCԾ��+�H��Zd%��7�|��_0I;����N��yEgO7A#H6�/#�gE�K��aZyd܂��ݔ"�$*&4A�Cܰ��>�e� ߺ)fn߾M\�,���2��ǰ�,0#�9qe��/�d��d�(:	d�d�,td��Û�kf�e��o�ɸ����Z)~����X����,$)]�P��$ʈ�(�*�G(�t�Mr���H)�̲�� y@$�#:fD�J�<��%���#	��"%?I�� �'�DKjb�sI����r+���"���xdGB�	�O�|q�3˄�%�H�9��)_�@&� q}�A Ʉ�~J@(�o�&]�Iė?9��\&���OQ2V%�O?��`��<dI$Bƒ=�Ƃ$����,0<���^��7g�㋦�+����<k������E���n��hA��j����������.77㕸����Y˵��8�K�%�LU��x�^j;�_Ri�~���9j�|9tc�ۭU/��ݜ�s��g?�p��{#K�����Di�����4:�6xJb��eV���j߂����d�b�r�۞��x��/"E����"cO(2I"Y�/�����в������k����㝞'S<;�[gE3�-�Sr�KuƩܟU�}Tk퍋�Gw���q�����ǭ��k���Co;.v��`9"��[W1	?��b �}���&����~
�@<�M�U�u���|8�-jo}���?�ض�8�����3���Ǫ��:����Wiy�,��ǧ���{����4�X,�J/Lp����4��%�`�6�;4@��H���gb�s���mW������Fŉ�k���+�L��Z�}V���E^��,3�1_X|�/�����x��_}q|Q�/j�L��;< =2�dHo%�<��ƛ�n�a�}�\��'��b�:2���ű9��<�������;���?,5עӯ7yf[�=���{R��`���mH���ǻ�1��2�L�;K�H���O�c)C<�TyRti������)�&�%�=̳�I��s��NO���_U�5M�\[)�5��]�h���A2q��X����`��Ƭ�hR�f�����?���R���w����]Z���J;��h	���h����dH��J�M�Q�2������{]I��
�1����t{c��o~��:�U?�˧ǖ�r��Cå8C\��;Z���s������h���Qy�0
0sgf�t:9/�_�������� 1��DH��/}������p�S��R0�<�D�ώ�����vG3�m�6�츺2Rpb�(́����d�������|����������1-����a_� ���"J���w�sY !p�L��$� �e#���6���(�Mk�M�Y�/Y ���w:�^����?y���m3�W�k�N�T2��:����K!�N[ch�ȁ�����{G�ʧX�Sq�)lZ�Ǘ?������_���<�|���/.��%���b'#����������+��b��©��a,��^e��4��]���M3Q�/Jww>�O��_V���1\}�h�y�UݔDtVYl?��.Q�<r&�( �l;SBE���J�0�g�<)�;���nnw��ٰ��~�y�N�����k,��L+c0���T��-��ztr<x�?9����cJ&�q ��2c3)Lp�����s0Ӫ$�$j���u$i0%<>�>ٻzmg2՟��55�n��k�-��`/PK�%�|p��vWW���E����[۸��W�\T;ͯ��7�dȔz�Z5l�����X�t.����tb^�3��e��ʂ�K�9�ͧ�MӃ�;֊�����ӿ�A��@�U��bp��!U���pq�WWY��[�CɈ�eltt2>��6�V;��m֡�d�_l(h_*�O��C�<��~��������������26~��kv��<5��g�:�O�TM]����䫰V�[j�dX�t++w���f����ف��{�*���>k�H�`'8����=a,���﫯H)KThzQ���z��vu�]Y[��J����'�����]��ݸCb<pѕ���'ŬX1�lI�
���� 7f��K]+�S\�.�=�..�{�j)O/%)T��_��b)����z~�dK��M\��h� ��Z>w�{�_��nþ4�O�(5�>�dE�;�Y��8 <�k��z��?�3�'O����˃N�n5�C^% 7��lD9wc����0M�T�z���V &��B	+�^k�9�/n\��v���K�N�D7������\D��ejM�ib��Vd�n,���4'n���=������	H ���a�Ң�3$�aO��F%�ėk
(;F�^`�����?4ῳa͙�b'����ȣ���O��+��z����`{��������:�v�lv��ӑ�4+��t�҃�n�_��sb�N
����2w���x�a6����mwVi�tq˼����Zݸ�֋ͭ&�K��ɱ!��3���c@���M�"��6`s�1cr���wǃ���H�a!]lK�db2ϴ4(.��sj�/�8�P�R
)�2�/�"���N;+�Ϗv��n�\��7,M���`,��u˝q��2�W���o�5��ҝ;��^y���|�F�T�Ԃ�V�	TS�N�49K��3B���ePfYy�_�]���o�N��z�Ľ���˷��������zy�G^��gƚ0S���q6<�]CCc�2�O�ѣov�u�e�K/6ٹ�6(R����F\ó/?ƨ��rm7t9⨺�f��m)y~�
;��
��#W���U�b�g�������WY{�R�a�xf~2����qī�~�5��������x��}62��0�Q��&D�(ٴ�Ì�M���E�2�?k��в�G���϶:�+�ŵ�^wc���l��-�2��O��2X��v���^��b o�l<���Ɠ��ӡ��d/	��RVxH�����V5� � ��J%��2�,�K�o��gF��g��&��ѓ>N���&�?�<�~�d�r�8:>H�����"M�E��n_۾~�}�����Z�~~����G�/~��G�G��qT�"za?4;�x69"�S�~�3	X$�l	��$�����`��t�I���b_5 ���2(��R���FX�pa�b��A�BSlS��J���S�=Vt��|gGO���Oʳ�f�ܵ�������������^<�W3�v�I��]��MX�b�@�xK���IT��=Idls��̸ A�IGDJ8��]ѝ˄�!I!ş�E�(:+����fI����R_N%M:&��G�-z��o��G��	��?��o�����k<��!.�x�N�`�Z|Й����w�v��.kQfL�F�K�@�p�&)�ťX),�~�V�v6�\��]��(�#5��
��0e�ac#G�<o����ƥ��
�j0�;R���E�����
�1C#r2��J��`��t��w%S�����I�����N�B�^z�`���P�EUe=��T9�|e��L.���w_y�Q@Ȁ�)���4C&�N,8K�Ip*J,���5j��7�S�
��|L�ĭS�E���WIN�ͣ���)�3����y�P�j���o5c��V[���~k��Ν� �+��!)��@E��؆&s���L.�V���N��|�8_齰�n˿}r8>�u���PJFb(�d"n�x�w�e?e
~���,�$2xz_&=�T�?i
�����p"�g݃�:%)MϲPDLj�YtDD	�+�'I-��aVeҢ@���Q��N�u��s�;�Pc�&���L5~p��D�U�tI�q~�If�LT~&�/j�� YKdt��|�f+�h�"޹sG\��|���_#"Zrļ",� }#ev��Bv��PfK�L!��Է��l"����?����#���w���c�&��8VN)#bP
�Kj٭��s��ʗ�29��,\I��4(�8�@�e��(AO"��8$:Ԍ"�S~�H)I���c��!l�/e�I�K�p \�v3R��I��Q����3'!����䀓o�����b�9N�8AW��q?D�_���V:lH�(� L�/������HB��X�0R�dV%A��)X���B�H����HQ��@�K\4$m8���IdQ8@I��RȂ �E��$��!���T<H��P�O|�$ôN6Q�/
��R�,]�L�qD ��oJC,bL|ЄBK��B��.:�E�t���b�������'fP�D��"˃O�:�������p-C��d��T2�(Ⱦt.#B3# ��O�RDB�7�?o0`½�����5���9i�U,����`����Kf.5ʦ���n��c_U�W�|���������>���d�m6��\a����Ŵx�ڗ�S�t�H��W�c8~��'{��    IDAT�0����n��!/֮l�_���kＱu����J��щ�Ν:,�q��BQ��2��X�q��:�:���y���x�ƱF�l2.=��QP�� Ǔj���Hc� ��'d	��
��?.��Y�?����o�\��j׮�t7]�_�b�Q�E����cG&W�����o���o��o�;���k�ͣ�Jɩ��S�!4	�X~%M�)d]X,��K�@��)쥝�̯>��U7��}���K/~���Kv�"���'�@�^F��.�����K�8M|�kU�^�q���d�dwvd�V��9��{t�=EUS�0e+���wVإ�1b-����S�D�3�RQ�N�?`,'��x�����N��h�J�Xn(��-�1v����x�/4��nή�Z�|����O����/k�OZ�擧S
���u�I &@ٿ��0?�`�H	�
Y!���Q-�<�d��w��ꕗ^y�ǿ����M�����#{�m�5�/VL�R'AN�X���Ι�����efO<�<��F^Bh��^�y�_��#�s�Db ����$�'��-L.���Ga[�X��x�%V+_Gf<�޻��/'��Eg�1��CԚ[�۔F�	c�H̫3;�cߥ�o�n[o7.���,�������_}1�ٟ��+��j�[hfM��{�����A_M���Bzx���b`�ļ�_��Tv��&�u�����J�r}���r������ǝ�mU'��9rK�1�)��B>1\��)�I�i�
����Y�����a���-��Ѽ4�x��m��Jy#~hB�Q��\4ʂ�?s�yY pq�e������>1.N�?魽�k76��^֢^X[��BIfv��=m[�t=�l}�{��g?�϶��m�Z�G����M�)&Z�%�*�9�qRg"��1��eh�8����Rq�,�3N�gu�-J��nM�_���nv�ܼ��>jo_1�n�^!�����F��6�(V�#2Uhd�e:0�;������`~�d��t�t���h�'1��-��p���B�~~�p��̟�(�˩������V-6xa�[�q+����z�)��Q�qCRTI���j�Ŵ\iyP�Ə� k+�+?���99�㳿>�ы�}pqh�8�&�����%c��TZ���'����E�ؾ��
��x��'��ꥍ�+���#ۛ��G[w^�+�J�Q�Yd3��`�뀇y�ؙ�?��@��<4w:�=<��Ye����LK���-HJ��[:r�,~�g|r�s��PN���x��tD1�`=rw�hsu��v]� [R��_��_�KɎ���=uL���ʋ�ή��K���+㓋q��'��`7����d�=�!P�F�x[�V�Rm���Ō�޵s�m��y�<�0\�������L�$J�ݸ`Y�_X�������S�+vלO���jyr:9:��c�01�3�l8��+�,h"H�
?]�Rc�f�9K*=�#�
Ko��M�uݒ�I��7O����B\K�F*e֢��h�X�3��,Oz�kѩ4���Z�����=���?�u<�=.����g�s��?�#u~� �ߠ^��d�H�٠ ��uj��LZ9^���<u��	�ܺ���_}�ǿ�Xl���8Y8�X�tケ�>��6O�{�(�����'&OwT���o�<��u'+�'���i=�TK<�����ud6	�sX�- ����.�2/���������S�ͺ�]sI�������j����T�:P=�O�łDI�à�O_��GߧB����?�}<:y�����7�]�V#��%Њ�B���$�X�ã�"���#w����1,���J�Fe�fq{jVxgk筍���7m�C���XԜ:�9��Xi�F�hh�8I�)�u��G��Ƕ:s��W�Ј+�9�U8?�!%�[�C��I�Q8�D��W(ળL�$��6p�W|��Jyg}�u����z1uqf�J�3w����t^ﲃv,���v�*��7n��i��j�޶5r���̂�pHtR�p�l)����s\������C�k�E�-w6W�������?y���o/+�+��j�cGA��h�����Le��Eq͎�>��b$�]���Gg��VuE;�Ұ�lB�-A�8G�褜y�l&#�{���%RMV}!�Li�M�y\�d�O������ac��џV���U
G�C�X���kQ��H��"V�˕��߽���g�W����i�i�ޏ>��tő&:�72AsVK���S%H�RM�C�8Q�b���j���7��W����|����.D�ly����j�S���3G�!je̮���F:������F�ӭ��힊�|b��̭��k%Ը$�87(c	�a_��#Ss��>�������nas;C��8Y_��}��`������fVw��!D�����9)p�͌�M�^P1:�ܙ��ի����q���E���Ɲ5OC�s����%��F��/�㙄����A=w
��]�(HJ�8�������+*�{?����G�t�������\�8�ֶ�χ�V��̅mL��BkYr��s����tj#�.���0@��6�)6���\q0��A�8�U^B�7E(���(	�S(�Ȣ����%&�/|���SrR���q�0,9�K�A
>�G��������^������V/�m�3b����_�?�����'qR�<r���D��"�7E	>�a����0v(����g=�<��%8f�'?���, ��o���/!鉩�ظ�lՊ�L㏪�BK:R��h�=u+�x�ֽQ������_�����߼���x��������|y�����_���wt��u%��tSC�%�.G����D��5�O� Y|bZ�%N�"@R�2b3�,:N8����c,`�A������<�F�EWmM}믪��u���S$�9KN\�Uxb�1�*a"�����o��9`t����C$RL�^2_������!�3�E�O	:a"�E�n�йn�Vnܹv�F�uѿ8=��'�j]eu���/<B�36$s��1IP,g
۔Q��)���ړёK��.�C�G�㽣ž3{<??��Of%��J�j=�q7k�JnB�XMn�N(�.�Ɠ�,T|���@�O~��⇙�%&R����$��@ $��=��2���AYZ&�B��%�@�� aړ�6�J��Pj�dU#�)t+�RRpq� .��w��t��eu�-�ڋ�g�Ìr���"��B9�F��Z�r�X��j�*������p<l��P]~}/�!b?γ��<�Ϫ�ܥ��a�ӺH$�m~�fW�?!�X_d)�W�ȅ�
�E�)|_Q�M���"]h�
�^D8�I�7�}Q^"d,l�9���%���� &�K8� �?9�	�e�Á�d2��2�Op_��,��HZ�t_�EMr�E��*gtq3Jz�Zo@G���[����\�=cy,s�J�(?
�B��?��?����a� �B{��g-M�,��F��(Y3V��#m�ܿ_B��ܽ{W�#��o�M��Y�4�"�2�n��Ώl'S�r"���¹��)QND�J���)=������hZ/�Y���$�&W~���+MB_|������MUT
R��YWN@�.u-��ɏs9�;Ԑ���<��B�<��-8�i]D!I`���'ES�Ił�kf�Ռ٢���ѡ ����۷�_�N�p0�2!�y'��IW�RVА\���)��8�-�*VğA$����.?G��q�_��E�/ �����&~8�AA'�)X�"BFe��'�$G�����E�����~��$��LK^�A8�<)�DD�.��P����s�Mh�St���?���)���ɉ..���Z�v*��DN:��&"��%3�$iJ��ob*�����z�%�����/W]b쒙檫�bf�1��fV�~kt���Jop�;���6�UM\�tm�۸��fO�&=u/u_�v�����7��긤q�|%���5~����"T6!S�Nu��vy���o�l\���{o_�qۼ�R<�>��]�`J�b��n���x�$�S䵻����ټz:��{x����M��W�qR�,|�$�I��0�'�(K?�,�2��]#>p@��`1�a������V(:����e��Y�}�Sd����ssU^ ��j�,����V��6^�}�w2zX;�ދ#{����1KBz��C~y$M��V}�d�O�~fA��)��?�TgM��K�W�z��k���a��I�?>s�J��p��X
Z�ݜ����a���?|}��'g��J��:��)��x�%%��})=�d~b\����V� p���Ș���-ϧ�qxO9tڮ/2x!7J��z`R�[D�Q�ѹw8u�ΓU��7�WΎ�X�Z9�=�ìe�C�t[�X�4x�3/�$��mB�q��pȀ\I"3���B���������{���n�����b��zrd��wC}�{����躨�Wb���D�Ո#g�{ӯ�\T�N�s���$����3}N~�~R�BdaRR1�r�	'���.s+�Cd2�#ܶ4�P�k�q���}�Z���l��x�n�m�FW׬�y�J�]klUw7on���z~����f�������4� ��r(����OrN?��+;N�Ry�d�׹��~����K7?��O7��j�F�2(�ʃ=6$��������Q�r2(�x�a{x�hx��t���/L��+��p��_���azE%��a������L��9�o�_,Ȃ8��P匒:֨֝���p��i��*��T��zl�7�ù�b -�FP]�sU��[�;wn^����{����!��.����z����zڊ4�W<�E����>���ig>j\���j�i);��N�fW��jo�Q[)�<r��?����R��8q��x>8^L\ I�cci�1�uy.�q=��xC���F��������F�r�ӝY9��S"�~xp�&r~~:�$�hěR��q�\ mM�G���B�1H�u'���H�5g�c'��#���2z�敋��n���6Qj�bw�f��]��]y�uMjE�-g��6K�H1Ïm���*>�B��!8pq뭦!�s������7w.]�����o�~��ri�%���h%�Ma���?�d`+���#c����ӓ�p��w����o��ǣaT]S�zϏ�H�0��r%c��)p�gq�㓃��a��}a����B�d�\��
��W�ӣU�Q%f'4�}�̵�U�X1d3�ջ{�R�ڸ�}y����G����ڊ����&.[�b3ӌ!�I�Xix<�eÏP��Ϻ�TDJ�G8r�Ź� �������7���~�Z}��3XO+���r�1�XY�	��@b(��k��������������C�{�%��Q:�1l��1ɥ�H�~�69Dc��AB��O5�O2�- a��8g�`i��<k�ſ��fqx�۲�5�D��b.?;�ٴ���T�-�ymsۣ��.���;K�Bt��68L]%C*M��$s<D~���y�;���,��� lj�as1^U�?k������ѧ���t�A����?�]Ln�v�}͹+�8���V�;��CG�m�?x�����g��fqOG�p0@�D��\�I\t c�LA<�i��/EM����U�L�GI[b}��w�v����0/�q��ʷ�j����iŚ1����=qq@��5Gǈ�q�ʥr�n�Fy�zv|������ƖV��h�D��-Ηj�C�H��^�쐼m�F��a;��y�n�R��V9��}��]���+�������R��(�g�󓃊ӱF7����j3fr]n����٩Y+g�<z0�ˇ��fŁG�b�&�U:����,D�������q��%����e̎[���\��j(�,pz�|�����.��	'S��+�v&(F;�E刣I���j5�Z�f}��r���;W��y�r}��p|V�烡mw��9l+@�q8!alc^[�U�!�Rjӑu!M���	���YL\1k�̼�Jo���>~����m�'�����.�������!d��/P�]12���xa\)�ZԓG�U�n��ڶY�3��o޼�1ϳ�X(�5�f�xj���/��R���H�9XHm�M�/��p0]>8��vV�Q(�鯦�	V�l���r�8���S�R�[�]xJ+c6V���%����7/�k�'��a<<bpډW�9FS�a�7�!R�Ďp_�
�O
����R�{̀���l�[/_���˷>��G��Q�r�.��-��\]��Q-�:43Dg��S9V�=�in�Ƀ݇�����ݶ������Y��~e�ݱb[\TB��1xư��mF+sDyp����Dr2�˱#�l�V䦐A_���	��H#��䦷um-��kαEׯPE�s˺m��u�]�V=���E�"���tb��Ec���0�͍MC}����C�iυ�������Ȳ�!���{�Łye!S:����z�z��ݹ���{���Gl9��������E���#�bu-�~���f�m�n���h�BZ�ʮ[X���r�I|�:hr����ZH�����g=@2 ���'M���!h�����&"�oI���&�D�C��MM���_?ӯ�W��)��/�r׷��a�{W�^z�����ޥ���'�|����?�՗ONOt�3>w;Qg��.����u�yaY
H�/LJ�o9�����v��ϥ�"Z�!=��)4󧯸b��g�y $�.O� ��U�$X��6�E�m���Yֵe�9��w������ys������5:�i�jh��diݓT�6���T&�����Ğ;~��沼��p����I;/>�(�.��� 8�'����0ñc�	UO6@�5�pme�k��\���_�����׿��/~a�Y{�*싦�믿���W��8���
��;�QQ̪� ��@��IR\~ڙ��EJn��!d�Rbp�����(Yri��^6��t��.�ym{�7/���9[�Ą�R�Za;1�oT\��M�L�nG<��0��W��M>(�dtl���xt<d������㋡��f�����x1q=���N�.t��*PxV۱)/�OOf���T��@�<yOO�dN�j�(�7���N�t �"p��6�a��Ҥ=t�-�.��Q�6�JX�(m��*Re�^���2���jZ��C]������PvӕA��U��1��>t�-�G�<d�&� D�}�t�(� ���X��8�~T`�`d	{T3=��ž�ip�F�#�� ���;���PV��B����-�*�24%����W�Z8ȩ�j�X��a4��"��)w�Dqi>��2��ӏ8�Z�EL:�~�2:�i2�g?�3h����E�P�dr�R*"=k�@e*�Y+}E�Lq��_�D�!�L+���M�
J|��/b	_@8��dZ=�I�����%p���R�h��$I9Ձ`�X4�(G� l�X�L�tY$� 0v�J��Q��Y�YZ�{��5��E����:��Kf0q,�K�߽{��L;+k�H��-ED>|�1p� 1@N*b%e@�Lk:'N���b�`�3�2%:�bީG�
(-VA�՛�q���_|{ ��&u傔Pb������(��D~����9��0YBDZ~�@��E�de>6$��+��
�d����](�%|l+t T�Q.� ��!���_��8����0��q�_|a�A��|H/E���[?S�������eQ��'��B%'� D'VF�	��f����J$]� �/�t$�O��iRHN�۝���F��Ab׹��b���\ѿ�V��FWZ<�"��O6��+
LHW����)� rX�˟����ɀ�B��<~
�-���7�O
����_�I
|,eh0ZL�&e~Q�L�O��� �2���nS�2���0��\ѹ�8\���U���8vh:d`
��DX�ʢ��}�`��+^�t}�����%w�XZ9��<}�G��O�*�WrygG�aH�p�T�8�%�9�7V���Z�3}�6�+��(�JSϰ�t�?�s���>��ҕ;�_��V�e�Ȍ�~����q�v�����bҟF���`�7������y��Nκ��g@D)�r~AR�J�<\�P��/�*(%,H����׵O�>S��Ή3v�2/    IDAT�W;+��톙D���a4.��'�H�0�k��s��j�O��|�_��W��VՓ~�83_��ڝǢ��i&�����$}]̕�w[&J��K�?�BO2_�j�V�l5�h�Ι�Krc����������WO�M_{��}�5c��~T����o1M���Ƞ���������O����ٮ-���AI:�����qF��"�&+���Z~q��M���lE�3��y���DgZ�	�iΔ�żؽC��\����w11."题,��Rc�a_RV��r�V�ҝkW����E��QXqQS����ţ3�[�[kk�����	L��Ql2�`�m�3�t�$SA����4�/5���+���J��|���~V�:�i��ay��t��49)F��^����1��kOycS�	2����?���a�ͤ�]
��L���/~t�ȋ֥�T���\s�
M˦�R����шh�4d�Ibf<�^����h,f�q�1)���k�j���SQp:Va2 ��Jm�/&�4����7W^�<��m�>�cùZsSΧ�9z6v�ɦ�#.F$��]KS����hȐt;+��"��)�j�8�UW7ێP^[뭵����/���?^��R1�5(Ϗ���/��.�6���8��|X�uO''֜�8uL�����ǕS7ܚw���tVO�݋6��%CJ���"X~S��2�.�dA!�¼+�M��$�5㺥?5��o;��Ҫ��͓n�f������qZ�b2�I�Ҹl�Rں�hM������I��Ƽ|��^��^��Z]鵩�BluL����;�w<�K�����E,�Ы^��Ѷ<nǽ��T8�O�s{_�^�,9�K)Ϳo����׫�[6[��ӧ�M]��L@d[6Q���N�q�j�6T�yr��g�x�1:��#j��Iq�����H[�&Z��XL�&<�)q���pqSڑ�`-6X��u�n����j}e���#�*Z�3�-���Rh\��P��c����jo�ͷ�^o��lo�o�yLΔ��2fjVXE�+�:���k�[l��J���}l�'Ե5BĠ��s���_��{�׺7�����Ƶ��v��K��d���5���W��C�4��kd<�a�N�^�?:�������I8���3�N�����������Á�It��<��A~���m4�CR�P4�Y� :��m��=�Z�t;��Y+���k�1�/��:��9��{������F���h����G5�w� E�6d{c��i��U��s�����Uϕ�������F�Ȍc(C��閃���O��6����O��OZk��1Y���%Kv��l,�!���T5����'�l�U�?=��^��މ7fs]��e�m�K�J�09�|IoٻN}�@�r$�����1�Pt�B�_th~*(`������bks#F+aݛ8���]hL��t�^��b�Eą�p����nC��;���Ί�D�]W;2DU��IҨN�5�c�l�.���Cյ8�Շ�X�,y���/��4ڊutX��ۨWz������O�|�w���Tz��e�/�l����t�G��nI�"ғ����<GG�������}�wow2�4��XPL�d_���V�_&
�$����ϔ�����6#�18z\Ve�O��>�3'�k�����-�ƨ.�G�����f[]�ĄF�cH�N����H��j�����nw�b�[5�U�֋N���[#j�RW�L�D��k��=�T��J�Ŏ8�m�rW��Ak���͇��;woޭ5Wl����~P_�^�g��Kþ�TQ�{u]5,���}.��D9zd:��ˁ�G'���W/f��Z�j���S7B9���T
E��� aL�1�+p�3J"_q�S�r�޷Ǉ�V����w�-�럨z����́='i�2�lkAzL;J�xQ	J�J;���_���Z{�S��t�nbWb�@������(061���@���F�� ��_��<��VY��K��-�V�X6�G���������G�ƭ�>�O�w�NNI㺁F���M�>���~cG�J�ư?��7��%�ja����[?6H6�Q�䐘̤�������!g������#����)[���'48�GLm�K��Dq+��t�>G���[S��a�ծ��]��8��8ZY�Y�kn �c�J�������4[�(��7u.���l����:=�bb�S+X�f��r���@��j�
�c�þ�0�##��z�|c������o�������z7�wa+���}�0:�3�`H�G������Q��IbS�:���3/Q�.�}s����x��z���j���qm���U-�yvm��I!@�ݔ�Eͯ����#�,7�-F�a�!s����<�A�{but����2ѡ]�, ��9�k]'*�N˽��0��]����2z�r�#V�ս}�}�%4z+���f�J51Ba�4y�:bRhQ/�_*�>�U��-
J���6�#��=�[�y��҇�����������۟}�槟.J`�X�<z89�w�����0M�[�dGp���7�q���p������c�1u��fEU��|N��C�(g��H���6s��~��� ���
��LȡɅ�gP!�P
����ADP���'�PpQ�}A��/"i����G�TAI!q�+_��AP@͗�2��\]�,�M:}�K��^�^�y|��?��_�鯾:�*eXb��L�ALn���N�������'Z2 ¥(��d� ��Cn�~�'dA��\�-��er<�@����0�$"�@)���z�-Xuv3Hi˧��9>n��Y+u{�߰w͸b��o�85�����{�5\1�;��!d��ӯ���\()a�P�D��O[!��_�)=�Y�t���0!,�I�,�%P��2����t8�3�f���"�%7�M�z��m��k�|��9Oř�E�Ν;��E����l�NL�eN:3U*F�\������iBY(�̤ 2Ϩc�W���d �C4�BcU�Hu$,���e��5�7n]�rI�1�&�{��ؚf��k��i<ʶ۴b��b�����a�5��O\�1L�{����ۺL��O�G������lp6��nrSk��Vqʰ�aei���������It��%~��\ʝ~�В��	N�I
$)$ܗ������B�S�����Q U��	C$
�����/���I��D��zE��H����_�miQR�n�ι�H{[�a���Ъ��d�Ib�K��_ԈȦ��c���<.O��z�n��|z<=}0>�8<r?����&^(��4(���K9�@:�I��)t)����IA�&�/��ίJ����A�)*|�3uL.#���trYy@D���h&)h(���� h�d�t�vf2�A���D�K>ŒP�7q@2�'J�p����f*ʑGP�?I�w���d�� q)�r�R�&�ĘqE�t}�04l�NZX"M�%C�9�&��\���S�~BF��N��x�� �b�b���2{� lE�VWGA	���PZ�!y$�Xr�2��e��U�Sܯ������/�s�0�yTV֑u_]}M_s_�;;����rI-%Ҷ�'����'����o�l?��E�Ej�{��=}Vw�yߙ��7��kL�w�@    *�Z����+�ܕ��L0��ʪ���TPA˓{�����E�&U��H�\��$~�(�Ig�B,�Mh0P)���&M�ZM	�ԃ��0�H֪&�S0'�<x���`�
GF䑅�ìlʐÌv���X�ol�1���
��e�J�/�gu��b �g�GsdɕV�*%�${O�MM�D���-(V5%����Wր��M��}�D��
,[��
$b�G?:s 8i9	a��XN���Q���2��2���,�}}}��s�Cmm+&k�8-�L
f��M��t���,[zP)�%
f%�܀�g��W�,�/�R�൵$	�g~��?�s�X ��?�
E/^F��(���(�0�xD	��&����r���'r_~�`DP���q�@�Kq�	՞��=��Ao�Lg=�<���U*ҳ�����f�r}��pwk��j7Oϼ_�j��P�ѻ}����[��~i�U�I�J`x�K����b��4�ޛY_�4�\{�̷���Χ?����(�-���ϟ9��V�dt��ŉ4{@�[��YX5��yf�������Y��A*��z"N��Q��?�En�I�sEjQW����m��G Q�O.���;4��zdq��$A�f%ft���\�Yug��zi���v㣷�O��+Ʃ��L<�l#a��̱2����aG_��I��vh�l:zk
C���Z��R/{�q�¸;���|��~���?,׷�v�f��|�n��k,2�(��L�;���bn9���ݳcӖ˗�G�.��3���MZ�<����"x���M��������'�rQ��Ŀ��	�>�~�
'�L�Y"���?0�5�EI�5���d\�kIS]���*6�
���U\�8_�<l�t��pt��͖�o{s�������%F����7��B�S�G�̚B}f�DQ��j�n����ii{c�O��_����l�Q:�R��w������7���)�8���**h*f-ض�Tr{���o��|�rު����3*N��L�Ĉ�%7&q �#"$K_�wRO�$���\��IV�L3`܋v��o�m&��EX�Q괚�7�&�\H���>��Ss�r頼��qX*���+!\�2���-��C:&ɍ�Ճk�ۻ[�I��lS�Q���6��ӿ����1�k�]�7��?���᳟|��?����/�0?�w)Л&�QE4��B��X �r����.S}��֋'�_��9F�X��vT�lX��X�p|�PI�`�׮�R�J��l?�k.��/<{OR[�m�uf��R][_3Z��8�K|TGlU��A~�I����4��CJ����޿�ƽ����O�ۍ��=���l@/�6L��R�{mc+�+mH�8Ǯb��5�������Y^����T�:���W㑎�����~������2�]vR�ܙ6OK��������=�aS����*ʵ1}W���������_x$9`�Z4����*Ȓ�hI�$���u%I�ɐ�� I�ډ'��d�|Nm=��"�7�P/��/��~��.j$�*FK,D)i��a�e��N�x��-�[;����p��jKr�V�e��=$�������ģӃ�(ve��0�	t)��������ȶ����;�}r㽏�e'~���lM�����R��Ĉo�S��Qgҷ�y�vg㋳G/Z�w�b	x�n�le�Œ,h��@��3�ILtKb�r~��jW���aE�$�l#��V���h;da%NN�9�?�e��y��l!J�Ph�.5*�YN�(-�Ｗ{c}�wܨ�]�R�e���U{�tg�Q�V��(�&�e�j�Ω2W_k��6��Ȏ�~�������<�bӿܭ�������/~UY����Ԝ�l՟L;�25ֹ5.�x�FpG!Ã�7�2:쟜]~����������=~F�+9�tC|�I�~&ђ� ��W���$U�4q�&��"8�B�3e�|4[i�z}���L�N9n;��4̄���N*�kU{'ΩT-��77�M6=[��*I������f$=��*������ыWh"J?��J� ���X_]��F˳�Fu�Z�m/Wi�|�����F?�]閧�%s�N;�;���[w�e&$����q��ީ��i��㯾�x9 �\j��f&���'�D�h��%�#�_�܋c����J��J�SH@H�C���c��(jc^Sb�2�_3^?��n��b�/��ckj�a� X}�	����ڃ����𙍤���i�I`x�.S>�����j/e�L�J��T0|w��0^X��m��r_��vaԼ��8��dSq���O��'���l�,�r�>��<g��A>"7C���d,�ʕ�$�7/�/���|s>�v���s���B�r�P�M��ʉ�z�52Kܴ����10�"5���de����f�~q~��ʲ�Ftn�7v����F��7,��>N��I@� /��&Ʃͽw�߸^�v�Ӷ�D�#%�[�V����#�z|t�ٜ$'���	��ɸ؉s��VĪ>����i[sa>jW������������?[^{SѦe~�&ôĶ=�L�֧6��2�{$�}c��B�y�P]���ˇ��[��/�7�<T[[qN��!��JI1SD�f���@�g�\�+���h�B��͞RP;�'G;�!���}[�,��"�y��ԄՎ~p���!�Q��M���EvT���+3�/��W��g�q�9l�0����~l��9;o�O) �%O\�ӿ�0�[u�~��7�~�I��Ӓ�-KΥٵ�����~��?�y�����:ȼ<�v��_�zq��K~�+�IB�7r�r�M��L��Q���O����ڢ��FP�6�0��ݿ�ws}����Ha�6�׳gϒ���������9�l#ėJl$���ݺr�ڤ��{8q������C̲51M�$��:�zP�>������9�\Y���?[v\��BbУˋ���k:��+4���B	�i__�e��*-�~�O�1�K/�7OX��M]�L�KF��ћ7���q��_���V��P�ȕMO���A�<��c����{�!* k��و�"����e�ut:��b�#-lmፊ�]�8b�'
T��p)�𣓺#�`hȡ�@T�1QH���(/-�t��ӣQ�+��/����A����b�{ ?3�T	/d^e�%O`�Y������#����m��O���7�Vo�v��[�����������Ƴ��
�'$�bi��'r�me]1�$E}c�)j'6C�
�EΥ Ze5�H�Q�}��J�)b�|f�L�s���')@��Z/���R��)�]l��,uR�F��ț�{���HX�9<��l�����{R" iC/����Y�Nh�,�o�G�v�6UA.g	�	�5�$����IFi����Wp�[�g^���:��@���#H�0�lO����֭[���R��Jy=-��Z��D��f*9�� �駟���;�	�y`TET>�U�QQ<� �K{���E«�9��j�����E��7�l���Nj�������`��l*#��T���{-����������A{64P����!p����d��|�58��@(h��wTY�[4��idp!'G_��Ŏ�M�l��0WN,����X4J�2@#�O_�Jl��e�Z er_�>??�&yEG0�}C�R�:�хעZu,Ic��P�mC �N樨hpPj�6�mvD&&1Q�|�Bʀ%f��a7d#S��(2���`���Љ��x�S��mS�~յ�Zyxq�b�U�]��V��
�<ئ(~P�WG��[A���u.�(*�Z��G*Q���?&B3�"���B��Y���Y:����/	��� ��WHf�&��2|&����E�̒�XfC���W�D��Wx���<��M���,�Z��rY��H��@0�Cd�B��/���<r��+�Y$~�1M'.�-��6����Z"�$�-+N�8��ƓBSy�F�@J+����́����8؄ge�	,P1$��2���ӧ�%�G f�2 I7�l��Ñ7
'/��D�
�*�I�:ܼySy��$�z��]Q~*?`�Q��B��+�p��A���J%	��p��$�
�3�6j+$�*%9�b�lk��\9M1���*_	@Byq�! ePc�ʁ!��d! ��.��`6<~*0M��I��l�9�Sy��(,G��{Vߠ�� d�`Y�	�@�I���2�Z"�V��:P~Q��%3�@?3JC����FɅd�2_y���s����0Y�	g�C��f8�@`H�	3#��U�EO���	զ���k�{Α3�)`�g�,[�Je���;Ze���\26?�%d�!a|�`�X(R�de(����ÉJ0�d�����$i�[H$ŸJ�2Se�2\1x�p�!���T����b����Qڸ�0��o�2�F�ɪgP��NcW�w�,'����L�a\HV�xp�����۟^[��mFɗg+�������     IDAT��E�����_��[���TKʶ�X�\k��VY���'����dwmyo�~�����w띏>��OW��elE�˭�A{���0�M�rQuo�fMr�.r��o�ձCm���ر[%(��p��Ip=�j��h�DɊ���Us$�Lf~J�z=NO&�O��x�%B��*�r04)����V����G@h�lZ����V��U��Xښ֫{�{��R�tlsk8�����ð7��uz�u���j��}bl��L������%*���G���tǛY���������~����ev����*���ɓ񠧶1�dZk�c�[1�3����>����y��V�M�~5~�������`���\�V耀j�n��w�L���8`�P!�|�d`���F�"l�HX�G@�
R?=rT��(��e~�.���`�����LӲ�ܩVn� @��w��ܺ���9}1	u���Fc�`smݹ&��N��!��\Ǭ��38���*��v5S[
GB����Zc��[�������7F.����MG���fy��D�B�qX�,R�CS�B�1x<	�V��ŋ��/͎�˥�U���CI�Eg�{ɫ�g�-�Q&�	�� ��/�O�S����/?�H��'JUL��ybh'�v|�7�����th�\:FByQj
jC:���K/������li���kw�7���:�6��\^����Z[]�;�'��=~rz�n1s�8���tS�`�u���zݭ���fe�2��y��������OJ�uƙ���ټ{Y����cq�Mq��8�Fg��O��龱�hx����ѳѷ��٧��I�Q7�V��H�%|9���ѧx�O���C��u�+ڢy:a<B���#D����!�����ƶˆWќ��uł2*�6�d�ܞ��(0��nߙ4v�����~ya��n�W�I�b{8�x�:}܋���Նc�:"�,zcum��6Ʒ�jm�jMY�-d\:�Y[].ׇ��ޭ�?��/n��ii�ܤ<;���w��m��0����g�� _��������i�g��/G�]��9pɏtGr��BF�Gt@F��8�W��&��9��
�& ���a���ba#�D��HW��m03�x���)Qܳ��(�F�a���XO:�wˍ��;�ww��l$�����Q�n��L��e�����!]����GVb�Ŗ�Թ�qd�)�',�'Vj���ˣ�p���}���u㣒k"���J�GbMۙ����x=u'O&��dh���}�9=o=~���Y�kK*X�сC�+��Z��|(̏:	&D��Iy~Nl�P��_S����(O���a�6$\ Ƭ��k�W]m�Ϟ;ZG/�b�M����.Q��y?�%U'�������Z��+]6ۗG�L��M:\�L6a8o���z��9�7�ea�bNID�V$v�H 7*�s��ꬷ0��������7����u��K�����;��.
Ɂ7���JG��n�|���h�ˋ��cO/�_?m?;�� ���!�߰kR#	�W��! @�x�	�G�fr؂��'�	��<�!�Dvk�*��m��7=�8ne��E��mv�e�T6j�`��3��F�Ǧ�[�(B���7W�H�1�?���mmo4�6�Ĩ�c�D�_��|qd�͢���I}��v���7n�'���ӳ���|˥����_��?}痟��>�h$���y��o��w������7И�<�!�Bn�L�Ν��.^�|��E��Q�����u��x:���;!BS�X�����\<��s"	�Z0:g	,*�lr�˟<��� �:��؍	�Vs�5S4�$�A�̃�	��'`�Bb�[l U��U��`v��훥����'ϙ!7���,RZ��{>WHhf>�4�֖q�S��@�3��`���]�1�4�ͳ}���;�k�7�����g�ŷ� �lZ�~5u,oԏ�aM.� <A�*�����V�Ֆ}��Ͽ��������jLӘl+�Ӽ[�[� 4�C��
��0��ܺ�ɓ'4 ��H��%6��u	RK�,� 99ye�Ġj��$e}m�Z�S�1ğ�@D�Uc�ʤÓ.��4�u�Q���w:��՝����5��GD��ɥ=��yrC�Q�q̽�.�Z�Bgl���Y�ľ��:-9bHg�KDz��2�Y�����7n~���l}���>+�0^O�&q������Y˩H�W��S����;6�t�23��������Y~S�B����i 2Fű�VՒV� R?{�����&e�j&��U%�3eu���WHv��楻�cJ��O&�4�7V�n��0^�M�e'A4T�g��
0(5w���.�0���G+�o���)��ꤵ���^˚���u���@똳�!kT1P�������G��{�_ͲH+όV���j�p{���ֵ��?|��/����ɜ��@Ԣ�jr�±����q�GB�'Ǽ�y��b��Xt��C���}�����x�ԑ��`2�(׽�r����õ��Մ'$�䂓�����g��.��x�EU�&�9��T��V�脶�������Z#"�/�9��lY��ʘ��C�k��&Yu.�\���I���5\�7��~�u��?��m`轍n�Qb+}�Q��7�(~��aR�w;-+Rƨę��4�YY�n,�bO��ܾ\�����n�|��~�?�|�q���lH��Q���}v<�\�S��;	��F]�"kE�x;7��T��xtq�p+�5��>��h����b�$rJ t#(�+ϟ?���F�6?&��J�~f��T<I�������B�?ȫ����H�EcFs�  ��e'�)����	� �0�O`>���ZY[*mm�@n������r����w�����3�j.kc0S��iK?s$���n������gI�J9��~0\��O?�
W 
�Qbe!�*$�FM
M&�e[ �X!�WT凍^�`�a�:�d�`�� d&c��s�<�:��뗖7�7Jk�4W�ض&������
��5�E�BY��V�x�S�5P�����%�R�O,��@��X�{]ࠒ��*+���)	x?9�8�B�;x�h��<W�δ̈́I�CE���sHRB�b
v��b}�>4�袉����E��r�ۖY�w�ܱ�i$Hź�\ʡpP�^~%���?��@~r�(�̉YY,w�
�ݽ��<mۊ3f"�@��1J��������q���\ ��*F)�R�U����=�he\��q:}�쟍g^�ڿ�9�W/س��aJ&c
f�2��=J��W���h�+D,O~Ց)|9M�_�)ֵ"r#E6�p	��g�	�)V `�X?��O�X�&:U}�c��n�D#�:���P
�n���F#o���Y��8���#&�.8g�w$���,��h�P��9%�a�]�M"��ʬ�b���U,��n���<;{r:�m����^�8Z�cd�sAvU��
O
Q_ I~N,���O!�$�\8�Ds[2X�*X�;~Fv��(-����x��:~�/�)D�<BL>x�CZ�ON�W��e�aK� 8��rf|�D��EU�y|��G!��y6Y�T��d�H��|��xE&�F��N�W�9�&9M��L�K٦2q��V�$�$��L�+GG.XZr~�J��4�V~!�A>K@ID�u�{�.$���A����"�r/0e�E�� ~NIJ�	O<2��D=�ϣ����4-�̏>|����֚De�G^���*�o���(�4EB��OV$�,S!��
��	zE���]���#P�i8ᨑ$M	.��v���b�$����9\�B�C���"�B*ڪ�,���������_?z�(7&��_Btȴj-��7>�裛7o��Q ԎCy!E��'�5�(�ƈep�V�(�����c�y�'=�@��	�jB���o_f�0��H���"��T�O�6����SNN�������J�p?3a"IH���-��L���P��}�Ղ��-a2	?H	9e�O:g��P�f�Z�A��x��Y����Лè5���	 �f���KFF��(?EI�%�bd���B�pz|��'���j$!��"�sUq�����Q��������pY ����< ���i3a�W���K��/��D!<��ґ��)4ױ`_6�Z�,?��\a�%��=X\�jR��t�)�
&7\j����J㍛ח^.�{��N�����Fmrz��٦Kdye���\�n����Fc�6�L�����E�߼\�Mnl���=����v�?���w��������R���f��ԅ"�(;=}�-���_2-��֥��ڳ�boPz����4G��`&J���dWBC~4I�φ(HM�!ү�
�E�r�|%�j>~�29-�eB�C��yl7j�x�X��=mQ�h���˙�a#��*�1l�äͭM�>]���k��{+�ι��l�QɰR7��l���]��o�X6贩W4�t�m�� t0��q�`�p{����������_����wے�&�T�TzG�n�b�9�<)�=����b�DC�0�°�qo�:���/��/z�����X�S��{���
�P�:/z�h����\Ѵ�U�S�L.<��G��x $�y�e����X���/�ҷjγ��ōhB�ʹ����偊�q3�x�Ѕ��񱷲�y�?�FeD����V�.;;n����*rpp�7o�PP��?iY��:&kNC��H߃Z����B���o���}��/�cĬ�Ԫ�N��cG�h�u1�ukR�P,�g�X��0���S�.0N<�x�e�Q��r�_c��z��ZI4�RIQ&��z��>��LZ�����T	�x�D��� a�6!���E�|�M豨�Fq��]�1;;�8Щ������BX�rj��8�����b�m�Tj�Uݺ��5}���n�l~�[�B�;��!�F�����񿱝w���O�({;�v�ٓǥA��7W\1{�^�?�}�������׶TJK�Y*_�G�J���T��1!wOJ��c�';���8���]m��E���f�d�>S~���+���w�5��RATB�$>�q8�K����<rDL?y���eT6��
QFbo�78�F������P����%���)���B�.nUf�����Op���{͍����r������	c|�©������ܱBW�.7�=$����V�h�V{`�Z�:�UƮ/�-�������o~�8�OX��e��P,��c�4���clx��ݫ��KO�{�N.�lPbE��J��QI��D�dc}���^�U�TxF	OJj#�`���%/��[�o"���\��6�b뗡H-�x'�D�X@9��Ԙ�ɍ�B�r�]���du��x��k�}�f�Ӽd���W�޹s��:�}5A�єd�#e3�J�[;;�k�~sҺ<X��^]�v����'��O?�����&$�+TK�6�~1u�DEV'x�v2E8f�=�����]���c�.�f��Naoބ�Q#��j_���S>_�Kݓb��
B '�3a��V�Ur!W��F�ӭ�U-��ʲ�ě���q�{���Hw�bk�a&*�_����&�F��:�ܩl2�~g�f㝛˛�˵�x}a�p	��5n!:;�𢉢[8�]?�ޢ?
����ͭ�w�X�WZ�Ϫ.��o:�3�o.~��?~\��hV�&+����ܽ��fG6豦DO�+��I��hw�×�z_>jz��Y'����AT�R�Pe��I�~r���%?�����O`�_T�
�⢤
S���64�!��&;�F),�#��ՉZ��*3E�O�,T��d<��)�������'��a�f#p9n���	�Jef*�������Ε�IP���n�`�vc>[�v�����=���/����������W��G����y1v��;��Ā��C�ew�	��E2�]z��u�dyz���Փ����+�dߤ��0K��`d��;��$��tɥ�g��I= <�V��մ(��p��<����4�6mz�;Z��u�6��˱�f�a���7��H7D%��ڌP���4��wo��o�i�+.Ag;6>}�����ᦫ_z�aw��iq�e�KCĄ9�3��X����g�U+m.N��=9\ׯ����v㇟�J�Z:���N��I�Ͳ¾&)D��e�,��� g�#��Y�������^>o�/��e!�}ƹ�K�g�n��I�>ɮx�D���ѣG��V��9���)䭈-�9?9D�` �H�J'bF�j^*��F]J !��[��}���33�ݳ�g��;����B�c�]l$��.������;��q��XcJ���*@�g�鱙�������$�y����l���f��K�����_w׫K�����~���������f�Kd�&/�'f�u��$&|6���яb4@FJ�A7$��ȗ���O.�����Ql'.���j���q��L��s���>��>�J��� ;�O�sV4��R�Eg�t��4T��и� ]猟\��d4C(�F�e,0��P���ٵ\��� 3�W�̃ ���l������jyx�4n�o4Jm���Fk���VÕӃ~���Q�۹0�wNv��+����u�Mχ������zc}{�rc����O~�ٍ�>]�nz$b��?�z�:_�q#uu�x��RU@�\�0	F��[�O�O�Ǘ��Wrcs��/Y��9Z����������&N�d'QY��Z)��`���%b�T7΢0��N!�wt�1"7�h��8]�F���I�7�q-;玩�����r�Hl͚f��̿�w}3����7�՚c2�X,�n��\����9�W��;e%����}�`sg�,�|��v���x�}X+�І�)�[���n�����Wӓޭ�����7�g������V,V�lߎ�'��s^��1��;NMc ,��A_H\Zְ����磶*���BVX��⡋�7�olƑ3�B=B�7�M���'F��� $0_�)42�@���)	 ���S���M��dK	�e`͙u���$�$Bx@�8��Wy��b��Q,�����/��V���/�rx{��z���������oO/�]*a�1{�aDGRl� N����Ŝ�C�8��*��(��r�fB`+
�oV9�$|~�vK_?3�Zp9Q�Z�9��rT 	}�b���,���df�F�3u�[Yh�(���mk�[&��ݰ�eA8�(��� PQ�g�)e�D0�%�S֜T*�������!�i#P��T �j��4b��BN7׬&f��}�W� 9>�9�I��O���nq͡ܭ�EUc��ե�t�9-�T����O<x@;M��``�H'�I��7�(�;���葥�Ar�iPl�����]ZUX�3� �������o!�
N6���7�h�B�[g��&��2KK/���=f㵼���%K��(����[ϵY�oe�j?;�hN��W�܊P�3��S�+��0�B`�Kb�U��BˣRj�����Q�?�!� SM�����G �l���+J�/<�����!ᮀE�I��O�I�g��0�$��<2�RQf�m�U�C5c.o��M>�5c׋�WG�m��em9Y3�0~��]�`�Q{F|�ad�8huy����BY�[���(�uׄ�,�V�k���s����7�g}�W��Ų�@�P��	̜��"QB�(I$I��/ N��P���+�1X��;��S�$	���U��?�� z�F� dy Y� ��M��6?3/_N�@�rY��-���_8`���2��7���&#�b�Z��'XB55��וV_}���{%�<����C.0p��*��e�bdI��U�� C�A��0R�Y��D	�I��ߦxʙ���S#��.~�-)� 7���f+N�,T�]5Ⲏ���Y�>}j�R��(k%	`�e$ep�]����h	�ͪ<��
Oy(�;w���G�L� ����!��	�U��U��=�IL�	�b�)r*?�طSDS�\r�*|�{�RZ�̚���<�T�/�@��|��&���/�n���AT��+\	�0?̨�Qʀ\� S�|95�dk�!Tk��RME�/
 Ûo��b�%�j��GF�d�`�0�A(J�m|�|r����x��/;i��ƍp�~�����H��(Jߌ�.by�	���@���Xh�<��'Hd{    IDAT��B������@m�`���+�5�E%s5Xq�!��S��+����0�gv�g�q ��3i+�&���D���e���uA!��GZ��� �H.m������X���(0��s�R#��OO�ha��?�x�/'��З�L�N�Q�S����N�_Z��.7���#(��Q��P�][�j ���p���x��U���Tw��V�t�2_����w���_ϟ^|���Gk���k�w�6�Mݥ�9k�L��c6A�[�v����]_�ؿ����?X�vӦs��CG������t[Q�x)!F�8.Šك�,B�����V�KF����֫֐�ݹ��1�$kǰ��ł���틼1)��I��j DK.���#<i+���B^�~��-X5�"��O�q�8XY��Y)�G��,:Rl8i�|�C�g��J�����"�R������?�<��~�չ�d�&/��rҚM���]fn���.�0�5ww/�������������Fcs��ڭ[��]�z3��-�KYO=�8پf�4��|N�N�F-�7;h���u��������֯�-�=՗�[X����vM�9�z�P	K��%
e8N ��ɺُ��5'<� �3�(���!��������[��Y.����
���t��@�G,xqc��	���M�樭��)v\+�{�W��/���y2���iw\oF�H��8��՘�����N@��1Vz_�䮶\���yk{��`�ڭ��w�nŝQkb�2h���l�C�l�X���w���d�7c�J'�ح�:�����oڿ~�;�����K���7+�&I�B%�@d?9Qp%�2��I&��'�L�@Q�������L?��U*���S��	��t	p!ic1���֎� 1���RgJ7K5-�V�*ͷ�7�U�f�����x�ͫ�������Y}o�O*+��w��i�jq�p{ԎC��A�t�.qy���>z���}��[�{o��V�)���7g�U'b�O�C��Mc���p��\q��h2��8:>?>{�yy>iO�u���������~U�/H(��&aQ��@tF+��4����~^���E����ϫ(�䐐vd�yD�R5����b��\�IB�`�2�-�C��S�_;u�ƺ����3�Υʏ*+������/�C�Z�X/Zs��w�����Y�vF:�h3*-�����jy�s���~=}���P��;wo�������K�w�x����ͳ��6*����jul�kPr$v����%��9{����G�xL��xLc�`&X�q�Ȃ(�E�L���~
W_�R�B>�L�T����~C �%���8���T�������1K��L�P�*t���U�W����٢gW��U^1���������Og��_�����a�=l��k��Z��wH�����`܏�3�ذ�x�2k�������޵M6�{;��~����V~h3GI�(Y]��v@�Sb����F��E9��2���ՙ�4'G���^�0a�N/�*B���O�MVDR?�a�.���r��XD�(� ��(!�*P� �k��g���9wz�:���^/���8� ��@aK�bC3���*<:�l뭴�/�m��Wv�J���?\�����!f�'���I�;���ɚ���8�b���Tb��x�h[ܺ�������ֽ�w�&孷\"��[JG�N�2�Z*[ț�Q��&���T$N��QnSI��g��G�o^\\ci@l����D���\��P^ ���<~_�(�i�t+a������b�M:�j�l#_HT���f9=gJ;ذ�ܨ�V��D�C�l�����P��
��w���ә�֐����jm���D�kn������_鵍/�l����ޭ�no(�zc-�$nk�+N\���F���F���XY�,��޹���?y��so>�F,�FD���{����7t�`�9��I�@hp&-��
���0	��dS��j=�����/����ϻ�Ő4����1�=gj���8cd��?ɎVȘLΏ��{�m���K�����Z-R)��Z�bk[�Y�mn[��ݞ�3		v�f�:���o�"����d��jo�� /��+^�����?����_.���gg�M7ѕzk�0z��KS��6T���"ӓT�.]ފ4����#���+�����{s���1C�K��	֜���׆��3��t�>(R%HC56������˳���I{VZY��0�	5�����m-�ъ�.��v2d.NI�l4�A�\�,�S$NBD�:�E��ށU��ٙkJ`����s7i,��<��5�f��.w���`�6w"��uD��Kו���mK�^� ��|�����o=9د��?�Ft8r����|6<��C��6Lu&Ӷ�_��[o1�gB� �@1l�v.�[�m��ώ�>����ƍ��ݾRu'5O�f��m��:�nFB��hQ>��^�^j���;������/�@[vݮMM����;Gg��x;��h���\�˹���	�0L�7��Չ�s��a ��`�<Z�oSY�:��ka�ҫ��ʳ�d�V߲;j:�mp�B1ђ���n�m8O.�����he0Yk�-���/Wfk�������w������[7����}ٯ;�w��T/;΄�+=[����bi{}^��{]Ox��Dk1dW�����oo��Vy��]p��1�N���<��u�,�5B��|�~�ut�g;�Y��D��l6G�9��26�1�Y�B�M�B��4���h��(��I�l_4��Ԛ,�G�fK���n�SL���<P|�߹py>u���i�/N.7{t�8Z/rAO�>��":֌5�lR��G��Z�Ԅܳ�1>�ޝ?�{kwm}g�7���2FX�6V�k�Y��TdR���;r�B�^�k^��,��V�V/�Z+�����n\۹���x�����kff&���[�S~e	k{bM�1���=����l]/�«��W)��1ףM7��LGe�*fq��EP�ۤ&�<Cp,O�O�K��X ���R�K'\� �K��D�Sd�����V�!�w����_*Q�f\!�L�(�\ɦ�=�Ѫ����Vm}��}�=��N~�w�����i���}C����a��� �y,��%K��}�ė�,^K	��9�����̗X&�櫾WQ��
d�DA�O�q�U[$�+�E^r7·�2�0$�G�2骦F�I��*��G_"`uu�|������=Ã���W����ۼ�J!GJ^n���%WdQ}�J�Ǖ�2�j,���Wr��@D��O�$i���hP.YB,��_*_� |)<q2���rI�]'�@S>rXH�V�� �����Җ7�"���u�*�T�|�.���A�L�}���}��L]`��H��`8�S ��6��p��j.<)��%Q`�]1΢�
��������V����K3 �I സ����6��� %݌�C5[ ��r�Z)no��.{ͣN���ag����O]G���˾�m�ά�A��t�����S5���w=A���M�D@(�$pT�p(�� ��\~f T�^g��!k8�	@r��y�ER	}�J���K.Ip�{E�l$Mj'!c�iC�7�[��GH<�]�E�3-�8=�4���E����Y�4�|�ɤGlhq���a�(F!bR(�8OA�ᝨ/3Q�1"�
�be�zy��eQ�O��sZ�iw"�T��˓���l0<b�z�2�W��2�R4O��1�(���p8�~"uvK�B�vE?��Yg*�W*`M��R`yq�������/$�90�\���)v�^���+ ~�E�L��d��kGǤ��&Sr5���i_��m�J[r]�g�(J^R��~?�f�3*��M)$�"Tf
�����_�����8�V 	Y�Q���L��'$�H�ܟ��7y�#�Y�Qq%၇�l�ט��";M���_à2"U�}�Ȁ#�9�bbBE�V���*9�i���C������EjY+�D��&��HT\e�U)��4�$f� ���Z9e�u# �(~B%�j"�*'���X\�8���`ɩ�L�	�tq~�d�%NE��{���ܰTUIbC
ŀ�SY�~�Z-��o�F[(@����.�'����d�a����O�5�)H5�V*��X`�TH�ȫ��Qr�2�W�*��c��S�+�6+�����x8�|��H���W���x`�F�������B�V�ĚŇN���hb�XZ���9�Yh�yAU�`�0#r2��Eq��|Ul�H&� �������}�W��ډ�'���@�����8�$�sBf����`%�����ϡXd��`�K��'��x +�Hl&X]M�������J����Ъe2^cG9a٤�s��c�vd���`���R��xo�L��Sy�Z����o��ϯ����s��ٷG�������zimc���l�,�ee2_,/5��8p��{������Yy�l%��i_���qupQ�'��fG��M<A92Y�;�Ӂ���gLڼ!��<k���s[��U&�+q4���$)$Nb�
�g�")��$OA��>�{�B4��H�ai9l�-�U�����Elf�+9�^�<�쬿l/��'kӍ�t��WyRS�
2V��NL�����p?�&�5�L�B�Fi�����d��<<�?K����������Q]�,��`_��.������݉��$[���l}ž���6��w�+��Q�A�_X�V،_�݆��/���T0N�����q�mT5���L��Y�~{��E��ւ���)漑������/r8"���~w;䁶`T_`�><H}E�L %�Tr_�֩�LJ���O��
e��_v�7�m�����]�F����1"썻Kj^��5�h�JgV]�ꍳ�����~�Ώ6nw���/�O=y�sr�kl��3o0ڏv�ř��j}s�ِeV�[n޸s�p��ny�Յ���ԛP�S�T��y����<Ԕۈ�-&�N��7���v���~�uO7�<�0��ٲ���4��%�IY��d	�g�/?�j�"�`J��d�l`�U 2��̨�]{�o�v��{�٫�ՍU��ٖM�5�=2�$�vV\��؛0���E��/lo,�]z��y���X�^���ӳ�?��vgp���(/��Xc>x|>�����-Z�����ʵ��͝���>���շnͫ�b�!&���N{���n6+eH�<D�M��R��y!*Q-������&����W���ǭii}S���9E�����d�^9[tN� &QF��B��F����R���g���«pIh�b@NQn+������<�jc�F��'R�8E$�Б��Y��{��M�L�B����k�~�/���>����^V֦/��qۑd�Fl��8]m�q֏����v���[v/<�T[ڻ~���?}������~Y�v*6�lWƭ�1ұ�1[
X��v�$�z�V�uѼ`�?{����昆�f�N'�R�`�$�6E��b Nr%a3�@F@!�������%!g�A�G�@ ��?�-z��P��,h..Ύ�W�Wk.�+mO�1+���HvRW�?l��m��Ѥ�К,�Sp�^q9s�؝r�����z���7����?}v>���_X:�t·�Fc�7{�N�s��$��Z��u��������w�]{���ʵචl�<m�XH���Uə�eN���G;w
/61c�O���Vs��e��i��կ�Z�ֵYht���J
�(!�ARF0�I�@^�be�\WĦ͓�R��+<�LpB���ú��]��u��Ǜ���u�4�	^���8�[�����f#&Mò�+�޴���X��*����Un��q���G�w���7��\\���'��>YX����q���eZ/!��w7W?���7޽��V����qW٥��Aez:o�V}� �"���%b�=:ړ�!`��:9�m��^��|�yr6k:Cg����I��a�cQ�p�A��ɜI��U1ə~��d�J��+���w�rZ$�À�'�F���0pFo8o�u.N����F�ν
��F~r�R1R��Mܭ��)�f�m�FJ����������_}������o��A݋�x�49��z�BibD(�M�ｾ����ؼvx���҃���]W��d��r��ּ}Fp��p0r�B�y��L��8��K�f+�x�Tw秽R��������?���P�����q�$�I�D���Uq)zZ��L�8Ĵj��� �r��:Ѳ�z��Mߎ��׼|���Z���R[�X�s��m3��KaCЇC7{��*qE1��Ϝ�W�;��Vu���?۹�'�;����>y<�]O�:a^������9XX^$r��BX)�+c;��x�l/i��;�7�߫��~N�s�Z��}��+Ọ�F��ǁ
�׈8,J�"&�*�ޝf�����Kzw�	ɸ8t��Fmi�Ν{���e��� �l�K�+��Raq��W�@�Mn�3蜤N�Ko���4��QIE��^�,��6mO�֖��K�%+QM$�	>{@��0�#0���D)d�ds��X-���4ʵO�{���凿��7����'�:�]���v1d�]o��P{�WGp!x{���+fڴ��1��x����m���xs^�|�5����Y�rpv����T��Y�`M�p�R!�=q����v��ٳ��@�vc4�w�h��ƍ��{����P2��'Q~,M]�!�%�O�L���ix$�bJ	 ŀ�"�֤�x��Υ��|�Q�8],�o�/�g�e�&ew@W������	J��b�ʤ4�=�1�6*{+KĈ�d�fi��������?�����S揳���Y�rz�r1^�6�Í��W��F=��&�-B�7��x����o�Vގ�a�&v�,�G��r�$!e���%�'z��Dj�j"d�A�s�>m��n��rx֚��tX������K˫�w��޻o��;��֓����\��Ș$́zBD!;'/��Mm�:e;����{{���_5i��y�۶���T��΂V�u�	����yk�d725���doRq�=���׷�,|H��Ə7u�goݹ����õ��}�eg����ۚ�O�='v�����;A�mo�,����|zq��Zsu���[w��xpk��&�n��E�[�<쵎�6)�
PO�hk��[�:�R��Nǽ:::y5i��-�j�0�	k~Λ9�/�DI�F�$):cB��'R'y�꛲Z��	,�C5�XiEi�ae!0��w�˘]ȬEe�<��`��T�� `��&�Xȳ0�����4N�Y������W�6*^����<�O�͓�s5d����!�(��׊�>����s�*���g�6�~�^H���\���꧐��+�\ p<�$�^Hf�_Qr�T�\���?,;?�A�mc~mzU���i�t��s1�==�uq����K���޹����v9`�7��[nz� Mh��G)0+japV�˓~�l�ȬX#��=���mr_�` �K&�	"�g+���~��%*��!�Q���Q5�iHU ���5D*?�M8Ӗ�O��?�#*_#l,!���]P$��%��VV吽�Ċ4�W�aI*�yUh��LԕS��B���[�����-zB7�[t,,YY!HP��a�M���ī��CO2�6�`FEhx�(;Z���m5�Y�N�H�굏���yw`�|�����{3�7�3�(v�$���2��Z�@� �*T y�7<�U�OI2J��	�˄�{o��&� �'* ���Q��`K��j~M��M�<��R϶�iS����6퐛��mb�p1C��i<�9#Q�h@E+}�I@Ŝm��=��"d�p�7¼L�Q�;�G6ST3ʺ���h�8TU��.�4ȶ5��,������{�/�Y}:Զق�M��`CU$*�TM�@�8�#B��tW �0�,��V �e��E����
L���*Y�_a�B	a��e�ʌ$�U����?K�'��H�O	��"���W�<P�J��9M�~������#�I`�� ��᫨��h��aD��L�:0��,�֢� Y�+H�P����%��5$@
�&    IDAT�a˹��h��*�1�  x`�c,W�Q�Nl�P`<�W�W�NR���f�H����^5m���~!�0��C�L�i��
#w9f3ـ$OU6�����P���-�|!���ܣG�$�y�T�ڈI�B"#tV��#����`�FDA��rׂI�'O�@��Y;��M*�PePI�r~N��UG�Ϳ�R�$I�B�`
�%o� -V�V�9 �Q<��|b�[{��j��X��'	�i�߿���?��	�*��֊���+�,�|X�u
a���W��B��P����DI���ˊ�S�e����$B�
K�oQ��6쓞�a�	�g�X����L?�H��1!�S��\�x҉���S��3	�0p
�I���d�T*�e0ţ�p�1�,�"�4Nɍ|Je!�w�����&f��)� ň\_�_�)�!L�bC"kI�,��,sb�箪 @�IԹ�9xi���~0	��'0��YhČ%��'�e���f8̒C�%)U�y�gbV� E��U�8s4��:5��Yo������6p�����%�qQ�-��z�y:i��[���B�GGe�[�^�>�pZ�Q����|�=Yr�D���}Ujv&Mj��]�������8w�d����N�
Ft�#Q�Ig�~�ֿԩ�~s�y�Bǁ�8q�Nk��3ŹR�TË��Bzg����G�i�;JE�ԏ		�I�%-d�tCx�������BĊJbf�f��?�#����I���1���9|{���N��˰�Ǹ���rmR+yä+���/�i�j*;iM{��՝���n,���|k~��k��x��-wZ��m6���F�ް����/�\ʵ�Q����ۻ�Fiw��f ��r�/#'���`v�l�MT2vz�X�8�ݯ/(�a[(O��3o)9wۺ=�|9m�K+��x+N_4*x%85�G~�9T0�p�W����%cA^NZ!������q�b��������O^��Kf
������tu�ڠ/�R�i�)����9n�b�6헺�n�:�T=���[Xި��J��������޻���K���gk�l_L�o��K��M�׽Z����W��s����d"n"W*{���o1��@ϲ��g��A�TP�&�-�q�/�����[QOF����ls7���bkY�U���5��T����3<�T�QI8 �F�F4�~����">�l`\�D��H�o�Π���r�q�z��^YR��� c��eHm�m<�]�J���u�ܻY��ֶmn�CX��Z�b~��y��ŭA��t��ɬ��{�<��0�}VjN�l�ͷ�5έ�0�Tӕi�f��lN;�S�T�;I�`�2��(��SY���ܨ���X�¶3댖�3����+1=�C8�y��SU�����br�K�T�D(YH-$�Wt����'C2*aC&Ԃ�ϗ+��]��t;�<z��Χ�ܩ��Zu�t�� |������t6;m�y�i�菎��jl-���Ye�L�sP����7+g�V��Y�l��`���ni�Sz���e��6O;�ӕ�zcaRe ~9�Yپ����>�`����{ߟ�w-~�ݪW6g]�\;�K�ƘJM�W͂��� z9j�����9}z<��o�[T\�~���zĸ���p(�t$mVq&�� �MR�^���/��& �A�V*M���� |�e����ݬ���*۶w������5N�4�5�@Bjh;	��
�qe�&9�CU�iB�Qj�Q��w?~��ٷ������j���2V�&ɿ�������g	��v����ܜ/^/�	0w�����<+��}�6�!ې����,����ҡ��	�Q�������O_����֓�6U��Сx�<�NV�A��Q!"��OQ(��!�����d&��殢x '<?H ��k,_������قK���~�xǣk�*E8ݴ'��MGbˍ����K�F�yk�S�{�\�,�ښw�<�3��q������w���ي�u3m�s,���p=�ǩwJ;��r��w(���؜�������ic#�!X�.`�{DS
(�m?5���������Y}�*���x�jPg˅���x�A�=yЇC�Ir�)6�L����7	F�Ռ�e�T8Y^�[ۆ���ٽ��J�Z��}w�����4��		gpfզ]�gINڳ�U��5���*i)^�8̨�}�γN��닷�,�8�}�`���E�ܛ��
V�pw��,��]ujp�Zym��l�g��E��1)擋R��� ���l�PXO����-�t)ZO7��	�/�=��:��G��u^5g��Zi�v'^���cg7yЭV��b�^��Pɺɮ��'�
�re,%����Ȉ���H+��j&pt�<��"��g�������+q�5q�Tggi�ܴo�n�e� ��v���Q�Y�b:��Zo�땲�����O��?{��/���_�_���\�+:]�P;X\�k�N�+t�Օ����'��7�\/�;+�y�Z��4��lМw;�q�qo�G�##7fm^$�_S!�d*�yԥ3���^6�ώ]�d[�����8 >�Zz_�6��Y4��F���7��j�8������ B]`-�樭�� -rEv��.���Vs-���_<��M�{{tx+�+DÖٞ�p�c�ԥOҜ�g�t����Κ$ϑ�ǑW�YwUWu�13=��Fr_d�W����Q��G��fk�y�����=�ut]��w�}G���И���D ���p �K_���,j���ެ�XTG��V����/������ٿ�/t�{y9��]���´��ԥ�Hc{b��e��)�Z��_��{�~��u���ɜ��u�;\��bk~e��,ۮ�ݩ?ZY�f6,#t4� �+��+��ոb@�}�s!P:�sx`5+&�4*m����F$��L��* �����Dh���'����:R������H�]���������Я����d�8���C
є��aQE{gu��]��k����kkU;��
cán��ڃ��{��M�|y�n�4�����ͳ�����1��-����)�U�1=�����GG����c�^���U�I��r��z�C7*�4�*�-C�Z�/{w��Y<N��g�$�=^qy=99��[�^3��/�j&׾���o~�����9�V����O�9ֆ����F?�a
?���^����|�xKU��xm�>EG6����6�?CX���N�v��!�^lS��_�j���(��wý���W}�?\�!��������?����?����˯�t�o�o�W�񖧧'�=[V\hҍ�M��J����vu��w���y������޷�U�}Y�>u�D�ak��3��������ʀ�`meo�@D�y%�Ķw;��m�V�k�݃��n܍2�����H�x��%3�J>;簔ff�bFK�NM��~r`��#J��TD�/J)h/՗��i-�����aL��'0�<��r�3V.��L'�����3$�����DǢ�#�qՆa[��vU��;�v`�m��?�����o|5�䫻n���jۘ��S�����!��`q��J6���0
�!8��(�$5=�$6?�Đ�K8V�
�p	/*s�(!2$O��,h	��E%�	/�Je��b�c�uJ~�������w�y����[\q|�<���Ղj�Io����AO�ɞ�'����z��%%Z("�r!	���Mi�N�D`R�)c�Y��&����g��
<`�8�4�(<`�rY���E��㏔�������i����o�[C\�� �,tq-���/�3��d/_��u���I��(x��P�'6!��#P�,�@xp�zw��5�F�UF�J�Ni������!�1���9���X����V�AL|�s���G�;��;�����m��F�<��Qc׹����٬I�H]��h��Ѧ �+�ȫ,em����z��X���c�b�d�(��J�����!��ʡXՓ1EEXx@Odg3&~��E�`��'%�����K�yB�q�e F8�s7�)v�~�/�����B�؋78>�XMWc��^���+�vǵF��[ִ�88 �f�����ۻ�.�F�u�����uz.��QG���icQw�|e�]�w;[Տ�a���(�UIq�,!r���.��X?Ee,���
l|-v��&N��:�څE�%� 燁Ye�p�B ���z�-� <�K'!$�p��I�pH����/��0��T~
L��T��v?��O�kj�J,� �Z�����IYPY.�a�
��UD���L�'N߹j^!������C	ɔ]b@�,Rb-���"|�q��-�l�53�Y����spZ� �Tg��Hqᆎ���|a�U/R%1r��Z9�.+�J���l��V��\��H¯f�r&9lU/W�� /u7�ʂ�/^��@i�K�!� n�XTrOF+<��P�rL�(G0��Z~��Ы_L{���]��kB%_�q�/��/����B��qIZ$�����Q��*�ɱ�"��WR����"XB�J"w��
 ��oPn�ղ�,Ѓ�r�\F�_���2"������<�@�lY��x �<�`�Th B���B!r� �� L��Y@�*0p�$H�y 姴�0�drQ�K�^M�H�L�Q�J�`�&�"�qt(��S��+bW�3x��6�T��d.s�!<��+w����B�B�*�?2�ǃ��#C�/�qa�X!~�,69 O"�$+�'��p`8i7,J�ə�O�$Ɍx$���+kH2?3�X���s�~B��±�[5��X-t��"���w��g�NXV���\�J6.�q=�|����d�b��M�z{�>P���^Zr"ʤ��噒���J��#L��W���X;o
�"8v���.�Ẋ[�^m�%�!#���ځ��i�	����|7�'�L�a�����f~ɀ�����ŭ+������h=:�C��h�Q:�,�\��lKx��fUq��a2�X�T��Ĭ6��Z�AE�vsu���R��L��}:������i6�rf�q+0��*n7�\-���ݕm��!����{����l~T����j�Iς�2����g�*J��"�?CC��ڡ�_���SbG�K��ƺ��1�d�ţ��~z��zҽ\o/Go�\����,�ͽ;��q;�<��W�0�;���1�)��+�Qɴ�d�-ϱ�$�r��RA�����j"��X�Oat�
�D�Dj0��W�_܋=��i�&2Wl�f5n�Ա��b���9ކ�nѫub�]Y�G��G�wt�`.����ť��B��X���
a�"K]��-����T{�2^X3U���ӴJ�1#�muU�o�6�"��ioz�ގz׋��݈zx\��c�H���:`�PV8�aBxp �ǃ��� K�/���G`�\x!�*�o��H��03\t�y�;d&Ӹ�sǁMOvڭX�Ĕ���C���.G�P�D�k���5lTF�v�q�ӚD��A��h�^V[ak�V���"0��I�3��$�(��ilWuN�6�,���+ g� d�R�q���mCpW�z�v��*�=Y�Z,���m��z2�D�w�'/o��s����5��'��[�fU���D�sd�g�J�W,�i��7?7�-���I�20%9xe.�j�ʾE��v�������P���g�-�U��{���DuJ�L���T>f^���+��N�m�+k�z�����j_|��-׃�����*'WW���p�xʭ��ك���c��m��;8�۪�}��������U�u܆zV׋��o����ѓ��#)�vb�u�<6qӭ=W�W�ή{�ZQz#�HMb����A�]T��p�$� �R��1��o��ME����-D]̟��jSS�p�$\,�D�zݞyu3h���eU�N��;�3�L{��{?a�3��,����P����{�{ԙ������(�����T����YU�����}؊����t������������=d@��z����*^�6��=��cL��ص8po�n�)L �⚅�����sS�O�/O���t����a��CXj`��[�L�l�6Y���0�OI���s�p}LH��0�JM.��:_���'3������]o�zMk�N�D3�]R��㸭�^sW�#%������孫�k�C���m�����Ie�9V4��`a�:�K����^�ܭY����W��_�r�۾ث,o��XNz�ɘ	�k֪���Lom�BW)�l�]e^Ж����I�~�b�sխ��N/��X�뷱0���	D�O���R_�/�01<LTpQ� ��v�-U���I��?'��m�׋�T�­5��I7.6�!�B�[Dno��*�1�eѨ:g3۲�:ZL+"n4���I�3�r�ݪ!	�;���\�W߾��V_TN���EZ��kǚ�C�c4;0�M��V�*��#���֡��V<1�c����q�����mk��n	�L`�K��n�{}{>��~��r9 ���ĵ�ۭ�=��P�^F\�F�훲!���\x��,�Hx�e�S�}8&��1��̆�1��t6I��
¬ ;�;����^��{����ƃ����'N�4j�sʸ����h�����Q���[�ո5m�v������Vk�`d�z7�R������O���O����6�Ϋ�N��kg``GE�q;1���$\��p��E\���z�T��bh��4/fPٶǐ�n�3�x�m\��.5��7���ӷg?���b��]�͐�	���GfƏ�Y�aRJC6>+��yf2�%��N_ xK��-[3_�i��Ȋ�<���xU�囦YE�No��g;�;w�f�.S�1��A];7b��4�  �.^�O*A�Cm'�5�ۻ^lV���jT�X|y�?�E�])����iupk��dD-ε�v�m���kwV>[��|�9�R�8�g�қ�a1!3��X��24.cv��IK��K
.|�.l���g�˛�ٕ�s�{;M�&V��Aϻ�0�HX�K
��Bt1���{$#�gԕ��H���s܆�� �m!aRY�IYNTG�es�R�͛n�����\0�N�)���Ћ�_��5�;�n����^kbkϮ�d���QJ�Z��ړo;O,ѓǛ��]uԛ��M��y��Zg��ש��e�Wt��
U$��vW,l0�u�p�-o.Ď�~�تۨk���V��dM�SK����Ӌ���V:7g�����*��|��/iKe����?Clb�E����JN�[�ē�y���5��S�Ybq���������mz�c8a�q�E�� �<�@�u�&h�&.X�p���V����|��n�覘eO'}7���8G���~����z���u�f�=��:{}��r����R3
��m��U7	�?��Y���γ�U�>ts�锉bЬ��D��������x��6<���aC��ӰRŬ ���:ٻ:�p>sw�=c��p;�i�>}��_���o~�����Tq�%?5¤�ėĴ�lzC,,0(,$[D�e�T��S�<`��?�#v��N߄ᇄX��4��}nt��f�R��5�D�Q�)m�l�Eh tv�wI��TM��|�_���������W/n�0�ѭb؋n"i.K�������Y@m<c��"�n �u��f�o&�$~rl`��ɴYƌ�Q< 9����Rσ <�Bb��`����+���YѮ���f��R��/��}�g?����Yk��n�tdf�p8=��v�in1�-���G.�J��r##�pYw��"���M���-Ř��!�r����XrC�pY�l2#��ᄐ��W 3�,�m��t�����
^�~�����Q�_�rq�0�
X����_[�;iGf��f�����V���@�Ql�I��,�/����ODK��႞�I�9��&����αGS���a����t�797|N�|��R}�?]�[�+�:JQD����3m�m`����jp�f,3�[,F3��mG�<�$X3�j��)N�+����W\6c��b�%�3sVjbH�����7�jEr��G*5 c�dvh(Jr�� �R&��P�b&D�JD�/	 &N{�؎tb�C����e�%�.e^Y M�5W������������Mwot|w��[g}2� ��Y��[�    IDAT��������J��+Kˉ�{��2��s�RL���%���M>�&�������.>�=�\�^��?���ذl�����YeL�( ?n��?Y!�O�����yl���֜��!k�.+y�J�̃� }���`� �	�sÅ�.QI+!�!��$ 1`��Y !I3`~�?os �ԪzM����ڹEf�� ���	-O�7���PKq�p�t��GX&W^~�`�  *���g����B29�����<��q��`�$� ��/ ��W@���1oЗ��7��\�9�(��rN^ҢS]�e:�Ͳ@@�"�6���ӧO���?����䘯,�P���I�"��1�ߪ���%%H�_��$p��������@f# �3 g�K#[��/�CK�t�t:�ɽ�^�(A^�HAhvD��zr̚��/t���);|VRH��)"QB�'0��.��f�(THd�pW���޽{�lI�C��Bl/^��J��B��Q�,cITm���Q����e*�@8����I2�\���*�O�+�$�#k�e-;`�����BY �G��p I�o�grT���O��.�~r0C�#h�2�`�O��t�:m`�'�V�i�s�&�^Y���JC?���r�V�}�LTVV�Yz�1��q߸,BϹ��l�����g��43�����#�?kK�tB�aC�@.����+jS�Y�B���1���&;��`��x@fBΤ�<$`���gb��'�g����%� ���< ��v<����?={�ř]R�1wV�c��٘�V&!��嘦cvp#�b4������Yﵶw���|�1���؉�^�6�t�F1y�nd�Ukj�#K��CL\4gj�8�:�Eho�jBNff4�lK7�ؾ��Z�7�뗷�w��ެ�&}󾝎I�V���Q�Af����-�WBI)!�����R`��܅�Ĵ��(��>1��`���Thz�*h�%�xcj���W<��ò�б�<z�k�4CtMpXXʔ����1Wzx�j`�0�wo�,i�[�N+��1���ېf����4zJKAU\hV\�L+�aè�|�KD%&�c�r>q803:�bZ�4e*�qFV���u�����7v���o&�yu�=|N�����9m��\q�<S��9�J�C���9���k�����&=*(���gS�Ο����Ė|]�GqG�u	�o�Q�0�&qk q�j�\E�Ԙb���sk9T�����Xrc���̰�%����,K���tXi���b2XMG��¢�,��ͦ�f���ڈ�*�%{����=+Nj���'�������junp��کO��IZl���bچ~
�(Q��6`~�H�T��ă�<�sЃ��M�gq�,,�t��u�������n�}l�J�E	�-�(��|hu�aiݜR��Ȁj�!w�4�!CO�p��j�;��klA*�M��C��C�(��6��ӵ�4&��l����"�8p�y�4X�\e�2�a,�_�n�v�Y�<Cf���M��؛����ʫ�j�α��j��[�[3tR��5�#��係$�R��_8~�s�š� �Q�:��<g=�8؜�!��&c���\�	C�چW�ʣf���D�Dc�%�q�`-�R���:N��clYk��׵��Z�js�mnk;@*� *���j�W���Xyֽ_��Yt-�٧�,Uۖ���r�����I~o�T����*�}Zt�u�\�-�M�(P٭9���^�.n��ƿ����Q\�f���-�Vp�Sv|cd&��x�{Bp/��(��X�\M\���!�e��T\ֈ؄� �*.]�'@no�֋W���|�u˭�������6�DB�E0�VC�.��
�6�z�΢2s��v�H̄U�e�[9�Μu�W=+X������؋�$���P&��$�s'�����L��li�m0�/�[#�iK�OܪǆH�/��pۻ��^^�Oo�//G��wb� f�s�|i���O�h�J����/=�K�b�{�OPbZ�4ؾ�آ0\����p�H�:`�9ن��I|+�7g^��g}:p������جcqTb\�I�c��^��9���8���0���֑[�u�^+�d����z�	r�c�Va�'��e���ye|����A���b��w ձ�"H�[��f3���֟8��t,σ����G'W�ߟtߞ�owZF�\ě�KbB2sx������ȣh�c�$�5�� �qc!(-�K�$*��H�Q�sVciCOT�����9־E�N�{eu%�Z�a`Cz��f�Pk	_�F�+s7�Y�1!ڭ�;���[�+y��p��7�0sS( (7���(����8�i�+�H��)��&b�Z�_�A9\4Ǧ���p`�<��}x}~�q��b~j}�$5;<,�[1�����+n|��^fr��;}M*�`�ozR8�%�ۄ1��[L?��6�9� ��a"i�;�OON��!
Ƥ����i�ݸ{�c�L'j��Rb���~K��wF��D�7n;�]�xM�+r^�r�g�XZ�c��֮"�]W�T��0�LV�d�����۬�����#�v���V+ѺFc$��x9�n�>Ga�v��34����u��Շ�o^�ړ���u��G��;:�stl���J�,�y)�2������c�aC|�T�OE�M�ɑY-$�|!/܎'!-�]^_L�#�(F�]�����{.��5!^�v����[{[�ȻIָE�bl����$���!r9����B�m����ā`�mԷ���_T��x�v�I6ٱ�� �V���i��9N3�{k]��ô�s��o����/�qƦ�C�#�ޯ8��<��kbe�=��J�v�xys1]m�u��_�V�"�Ͽ|j�Edg�%瓟d������⧨d]Jo�D8[�&�&&���S�l��Ev�vY1�����ߺ:�=��X�s��\66�}SlN��A̻�����T�ب���uÿf2j\������6]Ŗ�������������~:1E�?�tHKh,YD�k�=�.����v>��Pz2�45cb
TY�2�w��@�Lh�R/'#;R��hb�������7oƊ��k;��f��ѷ_?|r׏z��L~<�m�ZQ/M�I,Vs��Q>�=pb�/H�(����� �}�մ�;ۭ}O���Nb#���Lv�=X�/�˾1m6]
��ń&zF&�ʮ�я*^a����w]_s�X޷א}��!n�V��}�:��3<X|���+�I���3�Ӷ�����J3�ɍ�!��q��N�4nW]��C�.=�<�@���)�d���ܢ�l.M-^%�`�e�?ϫ�'��u����	��<���/����q�t��ȷh�M![���]���̕���K?��ɯ����G�l��+*��3�2?ղpnӬ�U�$`�V����ό��h *\��\�9�s�Ͱ�~sq����o~���QHJJ�/k�e㑚���Z�d�}e$0�E	N�@_���7I��B�o"#a�<��(`�i�N��`�S��Ó��y8��'y���y�_��dX�"4uIvC�C�K(�kKzg���?~�3����x���tx|<�zZ}��"0;*<\��k1b���R�B�� �rG? Q`��,9�Ԋ��b�%$� �s�%*Zz�4��bS~��O	3�B�+hY�M�VO��B���_;�b�*f�vn�e9u#9S����N�:A����a)�Yá���իW�B�4+|R/<�FV�S��, �鲨&��M-��,��c�����ШmEz�߸�$F=q�LHX��h��BM��v�`��b�e^�>l�	�i���f�	����=�:R�q�LY+�{:��Y[8!R�tJ!�y�LZX��J�,2 �7��b�����`�%.S%[ �%32"��@��1���ONB0T�[`�K���?���r��f]���cI�p�nie-SvL��Rf����aǝ��D��-<�e���o{���߱�ȫ��rYLw�������§���mF�#À5��Y��b����FGo�s,��1Z���Pֆ�`[2��[�B�����՞퓫�[�5�xf5�TџM�J�%����a�b���ğMp@ �7x�) �'``B ��=k�(�(08����%�\V��l�	.SI�?�J�'��0��%��u-6�����A���H�"\����DT���R~��E�"S"Br��L�<9 yR%���Z�) �s
A�rTD $X&�|�NQڑ��%�hf�P�o64<�vN�V�$��()�Z�J�$������:�-�A乎?��T��bY	�vj�e?i�DH�-���,�$T�p B��\B3��
TF�x(D��#f��/���<ɣt 0r8aF!(X���
:�2�l�����E�fI;�����C&T
�rɕ�d *������>?���$䈙�#��ZS��*H�+��@<x_�(��d�*��$�`�P�X�}��AeA�2
Q|g HY�9�K�	z����P���4�B��7r+p�?z��$ Ԉ/'Pr?A�ɏ��ȅ'���á@r�i�B`Q+\l"kzf�b⡀���<tJ��rX���^���H��z��Φ�z��n��㎝�x����ۦǔlX�%]����R�5j���P_Y
D&��L"��L"��W�+@*�T�9��D%p�4$|����݄��$%���@����fZ�$,��V	� �Iœ!%G�-����z�j���K{tn���aG{�ٶ{j�8�}�Val�n��.6��i��9��3�5�/���D;�Jv�l���m�)�9QW�8n2fx�i}e1ai@dp�k�K;<�.�+]gX3�˚-��#F,1���
Dw��{l�r;�_�L�=/�Ǥ�_-(f�.��
��W����)*�@��j$�P� L.~&�䰟YM ��,]���۴��7��7�u��Tj;�����n��9�B�X�1��� p]0�S�F��x#O�Um�b'�^`�U��=fݱ��NmV�őD7�N���8F�ag͊˸ԇ񇎙 b���*c�S(f��Y|u��������l����[���2�5'QX��O?5g���G,�0�_H�PT�?�i ��%�W�g8�)�-k��Đ��31rµ�<���X��rח)w,�żh�0(�KP�l�]v^צ#\O��e�~v+�Ԭ�8GR�V���JsRjǘ2.�"qE$٦:²�n�X3�K_��l�r��渑^�Ki���ٽ.�?�^��Vz;���Q������xi����E����pX��a�*�ū�W�9!	�+J��,�\ǡ������N�f.�'���"�mo8��R>�>6Ҭ<>ܩW�X��\O��Ym�S���1*f,!�=��95��\Z��G%�Tje�{=$���3B�ǳȪ8��˙S(�c�w����kf�/��X3)��4*ȡt5aa0��OF���nz7�ˏ�߾�/jG9�[�nJ�fR'�1�M.�	�\��O�_<�_��M�{���[�����v�0����Gϕ�$r�鑊Mh=��}��K�v�w��(^(fd�\#�HZ�t^�wi_&�!�[^r�y�t:��^���!��⻛<��Ռ�4��� Du�FUY
�[﬎��fc�~�7���O�}*y���CasE�=�� jꮽ�U��fqr1s��yo<D�V<S�?kf%UF?���%��(�Mq�jQ\&��d쟋.�L"�����7� �f�l���������k{��ʱ�z�K��K�¦h��^u(Ha��*���(>��zefU?�ʽ��Z9<\eƢ�c�BP��o,��$Tw�f՜��O�:�r���PXr0��g�ȸ�2��xi]�p�<9}b��������r��|������ۭ�,`g蛭�6�?1U�� ,ǜF�(��M����T����dB_~x�#~��(o�	��G'P��m�4\�߽}{����t���!4����m1&�Ǝ��l�&�**�DŲ��g���p54�PW��'De�I>1����x���&b	�9D����	1�'CJ�����AE�T/Q+�aD��9�M�����������/<=u_d���y�x 'FȒ'�ëL�`#Hu�:���_`dZ��~�W7'd��?3���$�)�Y>X��/(�������^�����B�I�ܪ�N�|�<��ff�"bXk���%���8rVo��K�8��c��ߔeR{c��0�ihaQ�LXҶ��X1x�PT�,ԇ�ftU���Jg�$˦��T~����OX:��x}�{;���YH��HB��Ir�)�R��Ţ�M4��7�c�3�'�F�q ����3�-�^H i5�M�����߾|%+�P/t}y����ړ����ј]�swͺ��-)��ki��-�-�䏱O�7Ml�/�#��l�a9�c��u���gnc��`���DF����U��Y�쨐0����j�e�E���˒fغ$�f���]\�.��[[(�Q�9(vc`l���^�rx�3�I�`����ԛ���W�o�T��ST�w6���d5 Nu 0k>992C�~�)�]k8�p�����*���[un8�چb��B�ʘ\���˗qrᘞeecg�vZ�֪<;��\�{�w��O�v�Ѓ��0/�[�i܎0��͈�T$�+�;�ea'����t��h��Qz��qߠ�X{���!�l�"������8W�ٙK�i�bg���Vܕ���#��'�?꺨k��O_-����I	�OV'��U�3,�\p[mf�/^Z��&���{��������U���W�ġk�Qy�գ�c��X9�A�v{9��rH�#D�0�t�W�n�Q���Ǝ�b]�>���XhE��ƞ���"�چ#�T1��$��eQѧF����i�.�\]O箫f���r<���>�~w9�.jzy/׎����}�����cd��I �\���i�����>���W��L���$���7j�Ԥ����/~���G����q��������;��ڛֲ� :�hY�k��7��kyqEm��b/N�#�K�F����b4�M�����j��M�5�g\�7����7^��)�a����j<$��ދ�r�����j1,�#v�Sb�D�W&�eu��S4��ȥյ֚$�C�vN��{�:�M���s��?y�ݯ��Ϟ�ZG��|�R�����I�kM vK�� �Nb��� �����D�F�
�a��&�O87!��-����s:0 � ��6ؒ��;�,�
7H�g�N�v4*m������߾<��F���MN�;�m���.�(H�A�x�!��b���c�H]BDq%y��$1�����T<���*������ff$���U	��&V��~B��>)��$җé�i�Ϩ���W�͏�����G�O��Ys��Z��w�o��UG�U�%�R�A��Nj�Γ9*EƓ�I�,VڤA+�3� ԯo:	Ar(Lx�^e��/�ra�K�P�̼0���,�I�h�����^*0,��u��t�en�|����FO�w�w�hT�����C	%��mZ	3�JR0~_�� $�	��
J�NV�a�ӟ�b��i�=��t�6����ILute�3j��Gr���`P���T<e�<vXyk��X� ӛ��ҝO���h0\l,}|�g�oX8�Q�B6��;b�R��X�M�@�N ;��l����Ab.�aK.��cN����&-��6x'��
T�)������6�$~�`H�P����B��I�137ը5�@�K��٨{��;�a�A��b���F?x�8g�'c�����n��^��r�$���#��Hl��h�2b�c�ta"7��'��6⠶��z��Q��q�F�yg��_<y~�T�~�L�Q!�y	om[,�Dx�����@�yh�}n�Y��X���3x����0ց�YT�ז��i9!�ғ���2�}�qpf��(K�à�|��W8���?��nGSJ�����xԡY��t�A!Ҋ�<�$%�E^�C� ����O��%r`\2DT���`��%�?��Ͻ�H&AJ�~Y�rH0�����f��%�p"�D����B8�Ϟ=��h!ZI,m��ȂH�VF����L���#C�a���ׯ�%m�_��>~�%9    IDAT������1�޼yc{C�PT=)N����B�5LN��ݠ��`!<�39�6yrk��}��WrA'

B��ŐZDJk������T i9˙/^�0R�A�*cs=XBP����qj�O�T49�T*H\�0��Zd@�6˽�PA"P���S��$W��QU����ϟ��/�0�" s �}E��Y�e����'��Q�H�
���2�'� ��1\ZÓҞB���P�T�<$�����+/5£8Qa�{	,!���~<��"_�_����ܦ�%�$	!�@��@�m��$]�8j�nU��=��W����N�nr`l8pQ�j�2�4��8�㰁5���v}Ȝ����m��a�JP�ྸ&�d���K�*�h����g�|�~�B�X!��~?��d]�$�X9B��O 0\�'�"0�SI�
O I8Y�������3 $@ۿ_?aH�dyK�W '$	)?9Ӌп6�v*6�ذ�?�"��qmѩ�5�nof��9ͺ����m���d9�����<�Ȥݘ8�ݡ�n��[��6������2�5GUg��dk�C�Ʉk���\a���2׳'�q�7.�UAͰ������Ewyz=�x����]�*���,5>���2~������)�'d�!�L�K������JƦT�s
#b��p�u����Y�_�!�n�WO�{���K�4V�UR	�0Ri �(U&3M/�X,��*�81��9H��cUsr۱ݶi��N�j�`�<3ĠX��qǥyn����l�H�]�+r9�>������ztcqs��w:\wa�z�v��L��! '��+兙�A.f�[��ٕ��
��j!�M &C�7�H`�B��� �T��T��م���J������yF/�n鋆`�d�F��q�,n��*F����مlb`+!~z���-/�WƐ�R�Tei������rH�4�Jc�!����RŖ�8��cu��`9\{����������?t�y���~kood��ir%W���@�ɚC� �N2S\E%s@
ɟ	)$=S�y8���f��ⲙd��3�ˈ�Yƭ���}�����;�����VD3�;���q��kx���i���ɍq�e��q�>�X����I_5���&5��FE`��u��L� �Q�*!���2�,��Ʊ�D�����fx�E�Y�%og��?q�Wo�FL��R�~�_��;p�.�̲�(��F��3O!a0��6�''$
��J��%I`���$3�B!n�/�7�W`O�|z�mK����D1��B<��f~��PI��ł�?����Ǳ����lmB��l�����O_��Hf*�i�Ҟ�J,gZ�7��(U�n��Z��ݰ�2�|7�x�����ګl���'�������,f2-EOxy�����E��IO2O"�!����	O�
�����J(I2�_�Ҩ.x��c�6\P�i>q��Ŝ4OԬb����d2�����1���hwl��}:�aW�(-UL5Y������`�I�:#0���g�VTWȌ����{lm�mQ��/��ʀ���::y?��t�o�����>]�F�Ƅ��c�T�#��a�x��Afqb��E��O��hc!�j��s��d�X]3��^���11o�g�����B@�i��Ƒ8�Ӹ�fEAHk�c������M,�P��~�B2�L�7�U�$�I��j��U�G��%Z.���O~�,�Gp(<q�sY�#ձF���|?H�D�"��pzu9���|�\�p�{syKs��;�G��'�ؑp;#�"����oz; C��0"��'��I���U

T,x_N $�A ?9���
��5����~�����݇w���&���ub�Hl��d�E(q�1*���8"����d�ض�p2<�g�%��� 6���l,w�8x�^�	����B]n-(�7C�
��U�ug��?�3�F���-�ehf�����Yu���i���v��.k�N���_���¢Z�"��A�g�9$�- �������Z0$�ę�|u9F�������dvs�q��ݎn���=������aڱ�+q��\�x���YH��WN���X+2,�c�8m5"r�Jy�c�f�(�SUM���|���Fyb�h�~���Q�	o��h��,��Ԁ��2)6dܑ�8��U�ϢB2�?q��ʛ���ǲ�"��!E���5�Q����"��<nccJ�)����Y5�i� 鏂��;q�7#Ήj��`J8��ê֌� ��zX�Aj{L�/��1j���{ڳ�5M*���M�.��D���3��:|ػ!�%.��+�\�GF�f��V㠶�#؆llQC�����>)~��A^�P�����!�QBl��I��k�xP@{���"ۓ�ۡ��oN�7úi&+s�Ԛ�� �,	l9��"�"�7��"?�޽3�CX�4�+C;EN�U.?��^|U�%�0�ҏ����
�2�.d�$������_�n�憽����n�֬ĝ��FlI5�����ҤؘRٞ6�mJp�MMby���Vgklh@�:QUf1����t
��ua�)�Q��)�Lyh%���JT�"�<�8��ѣA�Y�ƩX�Yw=|����7��ɺI�:-ð����s����Ön�.G�]}i��+p�Z89q��^�u!:9��AyY��y�/<N`}��\TJ�f:ϱl�3S�K���}����}Ϡu�EE*;�D�ƒd�J�&�ax���C�8�m&NW&�6�6[��m�f����1h��|"�*y'G,�Ţ���Za�݁Ŵ��ؐ񙣮�L���Ͱ�S��ڎ͢[���evw"�m`�wͲ�������R��w���H��s������gσ���/C�Ga��1�W�^��������o�y4��b���ȘSH�(_-����B?���˅'Q�y�	Uf�?�6C�U"ԡD.6$�Ί�H�<�s���iUۮsڪ���|��7�Al���;��iv�U�h�75����UJ��`�x�t�$%~�*XB}��OTq~��'ś����["�6���O�ɜ�<J6�����Z�\�� ��L7EH~��$b%���'V�%���@�����W��������_�S�Щ�.֖�*��'V��ƨ�MrT�ʳ���:�������0#������CT!pPU�-���|�������7%A�0�O �|�@{i������CV\0�,p2�HwiT�L����z���o
�tJJb�b��%�i"f�XT�J� ߨ�RmY�,�?������-%��!�����F�v[l[3$��ơ�6M�J{� ���ʈ��
OX�����6t���6v�P�6��t�������v��μ��&Z��	q�����AY��P) �D�Ys�K�*�.0�R�	=T ��2��w�~�����&����sX^�0���@���� �;�U�'�2;I�lBdam@v ��g����m�T}<��F-{����no��p���s�إ*��k�Q	ՖY�Ke����<�Gw&��Y{9�O��0�U�*�$#LU���v*��a�('9���3��1����}����.�u$;mT:���nk�Eƙ  �!`�;��DhiZʕ��=ҥ��rW�lZ)�B���`�y��c�����p~!�.��Y_�G,��X8sl *H � �^RZDA%����l��	�p~}�$�<�<�\�<� N��D2Q�L�Q��TF�����HL��xP�+Jr�����:_�)-��[����)����B�r�!0�w^�۱�es�_,RFY}�kG2�-�RN�C��H�e���,82/k?�E@��Ƀ0m�ŋ�o��|9@��
�0 FB�(x�7$��(M������B?�)�,0"���������2��jP^XD](�1tj] *�$ʈ~�V��~ 8�Z�a�i�H܃�C ��'�$%�ie�:�����_���Tr�Y�3R�c#�ϟ?םX����.v)~VHI�]v&'��ʮeLRT�?x�K��\`�QLd�t��O�3��
 ��H�B� ����2`�V��M`0b9ha�I��T�C�������P���HlDKZ�B�`)�Z<��^�mˆۤ&��ۛ����mw2�O��d�2����^�����ݻ�����j���Mc�dp�E�\b
Yx��rG���l0B�!~&�f���Q:_0��	Ox_���Q�G.�E		����y2I��Iq�(l�$pB���J�&�B�&1I6�j������`tzz�X�c]��0����[$\�	>.w��f�wjm+h��>e3���]�.ro�|�\Nt+v �M}:P��aa��ld@�sˍ4�H\�����9Z��2s� <���To�7�y�g�<w�~wtv=�����{w��x���2���>+�,�l�$��[����{�7QX'�7��3�)0�*ʐ�'�H�|V" E+�#8��rzrƞ��g����jwѪ�;�9��頱_а�Ԧ��������SҠ���A�,�\4S4�P7�,/�$�/a���iT��V��6��43��u�h�4y��]��iwpu���Y�����O�o����V�<oS���D)�b�3�%LH��(ȁ�F�R�`0}���OS���6����K[�C�"?,[A�x8�8y7p��gO����%e�9����VQF֘n�-�?�.�q0�+m��e�5d8#ec�ϰΘ����2�	�I,Ї);L�1"4�
ۊJ`�ňX�1Ld�q%�3n����~���p����o/��ڑ�����F~��<T.N�+چu��-DF�qs�����2��$I�(?�g`&�%���#;`<��e�Ix��QXl�'��������$'!>n޻�>��T���Ŷ�I�?�)��f�ȈR`̀�dċ)[,�1�V!-eU'�c�-��9U�[-�v�k�_����^�b��mJ"a1̏� 4�q;���Wf;���tt1oVm�'0����T����|V�
�BX
�ȽH/O
!�eդ4�����~�����%���Rk\&'� Ax'����f�Xl�m�E�v+�$�d�;8]
�l!{�ײ8yը�;��C$��O����9�Yg\�N���2��eNJX@��)&2���z
�ΫcFאn���)�	%�����̙�������>��׳��sV����`%�ѨS�_y9?�|��bX�#*٢�* vm��Hx�x�]��J�aU&�9cA�G��]	�q�Q�x4x��e�z�����n��s�:G- �j���+M�۳s�m��-$�*���<,���N�X�Е��0�����/M��%q68X�(E�cs��&TS�/,��6ڒ!���I��{}r��M�������>�֞?݆�5\�(˞�Ģ�/2p�۱:y(J�!r���	��9,f���vn�C��(�_}�L6�T/�[v�]^��4�j�+���ri�ű�q�8���-$����IIz�#���0m����}}ZgQj�;���Wqj��$T&!��!D ���x|��䥣�nVj��r�' =�sb��̻�>o�?~�x{v^����F�rg�1����l�����?��e
�_��ȴ���"??�A��`���\�^ C A�T����a�U7��1��������Q�� �桧#ߠ$�JW���=hm)�tC�#�gż���9e˚q׽=��a��ś���{��2�#5�Y��.L�V�x�����B�n����ӛ�����{���F��E�A��ßE�]��' ,RȒ{���3�\Ԏ@����#������N�daH<R��D��4[im��_]����(ظ�t:��K�T5.�?n�띶�@\K'#C�� ��[pU�}��U������{�1�6ȕ|��ib�c�EcbH�2��%���4��BB�ʠub{[�<�ANT��vmi.G��>=K6������z����IwX��k�7�����tv?�"f�t,JЖ��Y�)�Fw�޽�I?�h �0`/x.��W�_ܖĄ�t5J��p��$���wog���������M�=y}~���io],�ѐh�E_�7��hX����A ��Q�#fBK�����BÏv7!IqP�Y��=6Z5�i�+��·pJ��T�(y-��YNԿ�t�g�7����梚GY��u+��Iwԟ]�\W[��U�oW�Ø5;;�O�V]!���K9#q89��jJ������!�b�I ��~J�����9$��������1J�˿�˵� �PVa�;��7��O�5��v�1��s�\�!{�Dݴ]֡9��6�
z($TC�i�U��	E�z�\��2�aqKˋ�\������0����<&�:�������N�4j�bB�C��4Z����m�z.E��^���xi�k�c	پ�\�ᖜ{���#���ΧoG����L���7Mָ���"4(^r�_����)��H�v0YA��-� ۱E�����v���`�G62�(���ͪ�li�ڶ���	+!��I75k&o��N�Է�ub �����#��Xl�L�آ���1!�Q[��	M5wI��u��ދ���H��F^4+���j��b$�vH� ��{�͖�k�e��U�=�ݮm��n���g����KBBcfk�U�)�D1�1F��^
's��L~�fK����Ղo¤&�$�=�� ��I�k�� ��I��$���%I��_*  ��J�y�p�fk�m;���{��#ו��F������k!�h�.hP��{f9����8��$�����Y��3iK ��K�8��$�R�J�B��a�$��%R���N*y�LxH�p��\F8Y�%_�,I����B���H�$F�L`�i���R��kl�[�V����G���_�����������;03� ~�P֬�"[F��e'+x�XN�m~&x�H�ĖQY
8��I d�N`I*0��]���_�̫W�dMϨ,Q�.� <��;�b̏��?����'������F?~L����
�a/|�^Y�Y~d���3@����E'���P��~{�Iv/��_:VH��v�o.똨Q�1��q�*���-&�ѳ�6g���1^�Y�+�\7�v�����2�Y��ojU��\�8?F�
�!�W�y�~d��
�%��c0��$Ė(`i3X9�P����\b��H��3������`aR $����j}�WN�É����42d��8>������,�˓sVB���<~�wo��3�Y�����x�Z�Nn�����h�;~x��tl6�\��t{���{,C�r�L\Iڡ�j�z�&�qgQ�Xs�h� m+�w��ؿ������v36#��j�}u��Q���Bk�3�8�$_ ~��	�ğ���­0�ͯX��rA_�f������F���<�XU�D%BB� �,�p!<Re^
��&sN�,�ؔ���rW��cz`�|CB@
��,x2h9��i��K���d�/~Jp��c�B_�}�6� ��_*�?2	F�ї�
O�2�D�B����Z,�	�:|��O[(�����P��oN;B0 ��5"k!���$�R����Lc��S���"�!U��5��g�B�	�EnH�� �8z�᧲K�x8�MZx ���S` &J�R� %�(�F�P,���M�`0GB`��=B�0 䲎Dr_Yc�X�hCUR����L!�=��V������'� �P�Q�,�&�R6d��/����PwT�Hk�Y  �WY�����w�N���Qm©��@���ƣ\b9���=�RA-�fw���P�(���PE+;��s$�_*��@��ٜ�� ���O`�E�( @r���`2�T���!=	��x0,��e�a��1��곭9��ON///�g��ko�0���䨱��j��p88��?��'�F�`o�H�k�.&�;oT��])X��@n!8iH�"#���$���*x`%u��W̬HH�t~?��� �0 ��&*Ib��a�� 'r~ �X�g.���I�	��(��gfj�-��J��0�}L����i����d������gУ�    IDATa�ihm� �i��K�j���2�� nPn��N�Lxw�S�nzb(�9N̬LB��,��N-+*���������e����
�3'��3��q�7:���^t��7��d������E�������Z����"�p���7?``�g����G ���*��Lބ�Q�8s����(��I��(�..�I��;����q�ξb�ו���8ۋ��B��q"��L�t��/Y�z`�&�v��im�rA��}��8|����:�#VF�[n2�`���Ic�Se[	뼥�x������ݛ����z����|���n{ϋl�w�D��F2�6LH:��E����� ��	�_��I�lP�Gx"�*�!D_ZN �̬%Hz N� �1��*^�^}�Ǘ��W�����p�Yq�)3᧑���#�dː4��O���<ͶŒsl���غ,�.su5a\Wb����#sP�$V�q�$D=5,���A��e������y��i��\��b�~�U?�Ӳ_��H�R�T2}P4Ghl�I��	��ϊ^H~� �侜T��O"Ϛݤ�@�%�OQ�a�XF&�g'0-�6W��-.8�ZO
T-xm�nFJ�5q�Jy,�Yk��_�ܼ&�)^W���hde�;<�z:,�%C�p��I0d!�JfbS'�DGA�gn��W'�7u���Ӌ����1_�PG��� <�J� H,�z�6}��c"3S.�P8x_I���A4?�ˏ�����O�J�p��|���KĘ����%��q�����=}|��p�`�+t.;���iV�y��?6)˟��v0��&�0�	o���A��kRT��F�W0��×��JO��Yob+�$Am1�h)Xd+�d��/>:08zw:����M1`���ss���J0K��dJ���7�cK`.�\v� 0'�	 `�3��
��@l��0ځY�(���|!d;Å$�Uw �?#�ً�?��ݮG����Evϛ9B@��tAo�F�,0X"�!.�3� #'�F}K�[z��W��8'��Wj#=�M=�H�bT�mZ�c�n�\Tn)�^��o�|����7]7*��цBOV�ڇ�[��s����ȣ̛0M�SQ K�e���(���OI�u$��߰T�-b��+�O	����5[6Y��֭�a��nY�m�r�Be�1�� ;Χ���"pQ���dD&umx�EI���X ��c�9z�X�/2��`��pqBT�t�GJ�z�%���"����<۳��^�b����f�����ٙe�]��Q_�P,
N�)�J�i�M�dh#I����u�/��̲g�̴�g��8���%P]H���qX�Q�'��Ft��xt�B�w�Br�*��O�ϱ2�4$j�V8��V��$�5Ƅ��`{���5���q�z����^���x��z���l�n��r�g�:I�֑(�Y��	6��l�c(hy�m��������X�<���L�f�q�D\�s3���@HW�Lr���QX�$�1$�%?Ӂ�J����,u?�\���: I����&y��d����G�9��*��f<�{�@������?}(������x2Mn�hY�_í�
�i�?v��#wKZ7b������7���8ZJ7��)�u�m!�Pgo��J��e�~=��"�<* �0��t\w1��{�u���.�ڵC��:���j�84r�y:���4�&C`���8<L9�XZ��  8{7 YG�@`���9,���eɈ�Lf�	�w�K��m��򽾾�i:�׽�x�Z<rZ�=.YP"Ff��ܸ$��(�5��5�=딑���)IF���j]ԋm�W���S6R�p�i�����#� )e'�yVX�3cބ F\��j�e�ª�1y��z7{x�������p~�h�4�V���Ɗ'O�0���E8��ʃɘƶ���	�`A^�'��R �S*v�(@1�Qb��
���L:9����&IВab:?�.���l�vy2FR$�A��&��=�� �2�W�� 
��"�&�'Ew\Y��pzĠ&��&KO_u9���eq�l�p�ɰ�6"M�g�gn���Fr��V�-�M�ǯ>�gN3F�ߤ��O���ւa����n{��ò����@����cK�s��2�҉E$ړ� � H �f�b�`���`��/�X�d�e��\�}|�e���Z�B/ÑJ��Xm�3Z_t��0�����W�2������M'8�n2�	��8�%�A'N���>#.��Z ��t�u,�فG�����!�cXY$�0G��e�U�bH7�Ia7�5V��������I���݇Ͽ������[����s�g��ďu��!4�@��7*CmHOْ %�O�K&W�eF*x��1$!}�J(Jݥ�$�$�a#/�[&�I���|�$�@?���Y$N�co���jCsϻ�f~��c��f�~x��O��}Cp#E;��T$��`+���%����%�� �����K�L�t9��.��ob ����p�!�I3+#�+\�(`t�^O�}92;`�W ��RrOH����~B~!(�M�@����c��a��V樓���������#��?�F���{���6���e\tt���DG//d(�,�@�EW4��F=
�P"��X_?���ƅ�O�#^�������1
00!��~fg'�w��%��=���5����r��Çj�Z������ۣ�������;_�5P�h��W����Qʙ�G�I
f	�t��f���hUk��-o+R�>��r��E�ל���I��|�5�ST^��d��&�,�3r¤�V-���Vo����p���_�]�rʰ�"�a������q�7��G���/���j�^�ZQgx $,�	�J���=!F?X�L�g�����d�g��Ir'��Z��R3-�g8Kb9���{A�~R~�����Qώ��.�]��:3"3CdD�{~nU�}�����0777777��^K#o��-�@@���΃>�$Y����_{�E �y�%H�`��p����^��zM=}��g���no�+e��ZCk�������K�{䃆�;���yw|{ϔ���t�"+h�CbL�kDʎ�d�!T�;�A66��WdN,�MJ�M69��7���k;�k�V�{3����c��HF�I�
��?��-�R/�� ����@8!sa�A����$C�K�苮�
~��	O�?�/$�#
�"U���|��@�Dš/W,��R
GZ��'� ��la�N\�(����4P\&����B�VI��X�����~ɷ�~�}�k��J�N:z����]#X� H��ªY(K\n=�SkZ�HQo�$�b[��� ��Z������w�DS�u�JG,���jIZ��[���­<B������J����2z�E�w�A�dGP��P?�!E\I�ȥ9�CC��I�eE9QT��%��C�SAE���0�Ȥ��QK��r 4��6���>(G�i��ԕ�ET:ʅ��EV��r�O�믿�9i�Ye-S�1��
�+���B?x�Q��ƌ,�J��+�!K�r�M*a⧊[W^�"����ʏC��(�CM,Ť�e���N�����X���'���F	Ap���\cY~�JK���{� �S�OpN,đ%y_�#�S�� ����$՗=����������ݼ�`��7�>�vz��'��r�F�:,�耏��fo)���h�ۿ�J���s��J}}��:�ף7` ���X��5����f4\�f�/?�p%&�*��T٬�ʦ �A*S�YN�}�J�"���$-�D/_DD��8
��oy�*>y �\l�Oy�p(Yn�٬���U�,��p���g��;�6o� �>�������������C�S1�f��8PCiD����s}�$3�53\FM�緁jv�+��|��Ü�H��b�4��쏢�W�XZ�Y��L�Q���u�n������Ѹ57��)�X��QE%�7VK�+��O��^<�� [�
�-�c��b�G��$AʂGD"�:�R�
������"wG������N���۝���k3��K��1�(X5QT��n�K�l*�S:��<;�T����?u�+��~h���.a<(�m]C��� ��i3�
S�r�؛5��.z��λ��n����_�\M9�)Cn-�6���1#' �{�
^y*�Rr$_N"J8�������d�Ї\2�eX@�H����3�쀠BM�b9�`�c������g?�����lϮ,8��	H	P�a��A*���̟�&�>���V4U��M{�I�9=#���D'׬���3d���!��6}�6YF��п����7o�m��޼���n(�5W]S�TUO%���'k���l�m�JM٢ %�RK�(����	��D�O�%.���I���+���~%W�H4��L�����mo|���nv��o��t{~i���v�0�4�:g IʫK�y]��D��L�=���±�f�i+�	움��e^�R�C�E9��vΞ���u�#L��I��������a��~��?휣g���:��O�/�{�N��&��"�&sbI�[ˈ��S��灌B�q��<Uj����4��^�3�
c����G���7��g�6n�n��/M���cW�9��75"�aM��Ԁv� �1�mQ�P%+<ɷ�պ�20u�-��	\3����e��L"d�@F��\��`�]ZB��N��9|��w]�bj�q�����z�q�Ld��T�'e�I,-i��pյ� Z��<���A8��p�V���	�d���6��g���BM'�w����~�<��B���>h \vM\P��qe�n:$�:��+ɏ�,�e�y%c�%U2�FGԇ-&W��A1���9d�Ip���m_�\��==?��)z������7�烙��u�K=5�M���'��8���"�B&<�I�ON��\�]ᐪ(G���S�UX<HMp5�_��t>fiaQ{����¼����hmv����
�>{��:il���$�w��#��g��/��2(76!�L��#�,����dg=gǱft�m��`�榗sTݲ8Ƕ�̤tZ}K<��o=Ȧws����v��O��7׷R<�Yp̅ff;Ǭ¡6�I%*����H	�� 7���/H�\��%S�Na"�8!Y܊^
M�s�?�����h��Ԟ���ʚ��ƺ��o��@��ƈ�<jB�^�FNy%�@��J����yBD�C��"Vq���<ܣI�F
s,�Z�����~Y�S�{�[�;���N�\�.o:������`v��ъd������F�J�%$k�!!�d�$Y+;\�$h%h"© ���W�!h|g��/�XU@��� ��������W����c���~�>����w���u����g�/��DGZk����	D�A�L{D~:�$G�U��U㬖)t�NkG�u�1.*1v��`WP�G�� ��<��1 $lU2SQ���s�T����vN�^/���.����Y���ܩé�͵ŕ5�r��ݍS6��j�.{b�\ rh"���o"�D����J\�������ε�F�ơ�m<&�2�)���´�o�����x~}�j��0�a����kK����v|�mf3˖;3��Ҵ��'.�i9)HP���"]iNޔ�>:�"�^C�?�qZr$��cl��SI�w������xp�:��7
d��w|4�\^�^���G�Ϯ]YnVui���i4�+��m�x��eQ��ԗ`��KD]�)�V(HI�O~�%=Q8��<	�f�T�0�+�E��ĕ�isB1`?��I�����+q��=3ޔaUuk��L��i��<2I�L�x�\qE�|4��6Gu4Uo�Z�ױܱ�R˪�z��#s��JF)�v�+YIͱH�ߠ߻��r�������~��������ËaҘV���<����=J��f�$����:���8$��o��R�K2BV~�Zs
������֔y��J�E��X��Q��՛Ņ�������w����m�s��?��Y�m�/"�^��[
�5��Ϟ Ǽ�#X���MxIT��Oۈ��",r6
b�n3'�ń�gEk?�N7�@�����R�k��σ�$��eB;�&%�Mf�l3�/���Y�vmH����������p~c}ms��?���_>_YJW<z6J31��I��E���HO�A8D�q�O?a�d�W�XMBA�_��B(d�P+�2!�|©�+̊UA�j���8B�N,p�X�J��Z&nt�ewi�~ey�6���Қ3U���''Z��dAGƢ@�1�z��ȸ����%T�W����I�O�����5� "'
�����}�IL� �Pd�&@��h���}+"�����8Q�~��At��b�E���S|ʅ.@Igx����e��f.�Ğ�}��ۍ�͵��Ź�۩����֖��/���f�F�Ԉ��Z�	U����xÆ<�ɉ^ȓ/��_(�ab��~L&�9�#[������kƖ���f��G]��۞��T3��d��_�Y�0�g�g&���Ps�)�FH�]�F���.�I�+��VNP��O"���G/�~[
\by�r�p�x?����&��`�mØ�ՕA�,���a��sfy�h$�!�:��IkZ�wvxa��99��}�(d���j���e�7a���LaS���I��K�0�D�<�㐪��͐�׊EɊŧ�p �ȃ� �E����'s$������j�,$���|�,�j���X���_�)X�R��D��>��ެw*�Q�9h]���O�:G{g�G�F�l�tIj���g�g�̯� xd���':��]�l�m3��G��?��] Jo��~�	1��L9��S�w)�;Yz��;�Y���O~��Ow��~��\�Ș�n��E���VItr�K!�dc�����I�0彬�_Dh?v�pBɜ�!+""�<���5�e���C.•����*�P�O_�� X8~Je?��+�1�'d	&"Ս���I�B��4��^@t`��6��g�e��)n�/�O��}�nԨ��$�i_~z[�%����/~���t��?���i1"%9	Qr�d���I�np%J5��&�jL�&R�S(.Ƙ9�Y"U�����P@q��".QU�O��'Ϋ:K�$�{��jɊ&����ŕM������%]�~�Yu��ٳgH�6�TFU�r��s*t���M���ɔ�DSBB%�r�B [@�x�� �&����A�'��K4o�m���/諯�R�f���d1&"'E�CƒE~���?*q�D�~�#9A؀(!�Ȁ���5u<�#~r��	%vlS�I�H2a�X�x�o'q�Z�KCH@Z��?L@_Ȕ ~�AN��8���_\e
�2��O/��~꫙�S��I\�Y��][���:����nf]?��YE��L���׃�g�ʕ+�K���-�n=�w�C�n���a7�1e���@��=f!�	�)<��a	K��s��28de4���!~���{E,_� L�J��O�X�q��>����/�
"�f��� Dʦ
@5p��;_�% �2�\SG����(�=�Z�xt�w�}�t�z������)�=X�p_�rhg5�L�%0�"�:+��Xܺ�=Ȟ���T6g��R�S;�i�+Qt�M��>D7f�u*(^FA�)Nj^�gNϏ�:'���ոs�u.�SN��l}����MQ唟
R��'ŷ�Y����?:�SP�m�"�"�v)��cA"V�i����P��P̅��heװ=R�Q����{Qejyzs���u��'�Kf:�
�}���If���δ��_�����eQB1H��Z9ن�eNP�=7��7NZ���f�צb���B��?<xwr���;�zur5\~���̐��x.���'gL�" i(x�6?�����e��؅�Ȼ�e�T�
�+NK�bU��,
�
�UR~V1�X���e0-��p�^�@�^|����{���n
����2����A�Q�ft�A�^5���/c�X��BnMn��QE(c*� �v����N{��8<O�N-���T����E���t���w��oI�Nm=�]\�jM�=��7�    IDAT[Ue%�I�H�GY��i	�)X&�J8A��![��p (A�q<��"V)W� _i	��ʮM̪��4z��?�G�7��K��W^|�>}c�j����3)Ę�1���Ov<��e�ԵH̼F5\�dKބL2�G,��B�/���6�l�+J��ӝ���Û�p�v��9�yqv�z��;25��1�U�:9�mv�~��1�l���nc[B
�Qy/����x�H,2&��!��*.8E ��#J��_B��W��V�x�Kа"�x�����;ӰW���f^���;+3�y��4���^;5�&�"��TcM��'��k���L�;��|�6TS�J�M��Q��uf�hVv�fF3f,R� 5�����^��?9�?�������ۙ�����Fn9�4�$<��'S̱k!��'ݞ�җx+���B2��	ɧ�ip\�s(��G�"6p>�}q�7� 7@ȿ�	4k�f��/E�V���ݛ��=z�bk{��nqzy�z<mVK57�M"&��tv�d�͈2�i�LA��C����d�������o��/�ؙ<0��j�]}��~�͇�{W?��\�ӳ�v�!�z}�jn�(*��.�E�$}'b�ǒ���O��T��T,Q@J� �d~8r*n����)t����	�YSN#�}9�����4{���_�ٳ�9&�r��� ��^v6	�zO�����e2����	����[k�ՊR:���-*So9�bܜ�mwKd��cӖv��ƶ�y���d��n�|�zfo�����^��&�4��Mz��/�+���_��3q�1hٷJ��	�����O�<����0ᗴ#��:�EQ�� �(zt��S��񻻴��wۏ�.՚d5�Lb@�L
QWA�=K�LL�CW:���DN�2���&���@���*3�ź���j��eB_'��\��g���0������:痣S�j���S���N���u��)�`�}�ɚ,ˬ���	��%�'MJM+?ydA���'"~F����M�&L������\0��0����m�ƾ}���u����p4���U�������f��NU�82o�Z0�\���H~4x�̕��g�۹��q��GҪ*�h���l�E���F�M,����%]�l�k���M��#F/��7upqy~z�=�wo=���1fo�i�)]��3S[;Y����m2��K�79�'���N�&:��.�Cb%a%=�����K�b�8��/t8�,�Yh��G�.��GO��~����W�e�H?y�׽���jL=Q��i�D�G��Z�4��^��8�јlg�2�J��Ǫ:ʹ�u��v+&����6�s�>d�==A���2����ƽ�W�$<�V6\��aȽ}����:��<ڒ�AfFEU����ŋ?��?����鞟Ȗ���� �d�uM�J	I^����	����YQ*.Ql�m�kBZE�!*4���N����?R0���)�~��������R���#j'�T�-��L�,��Z�&�$�X:c�[�6F��Ϲϔy�K�J��kk���;L[ʶ�@rD;���Gs��)3����p��}~zt1썏O./��]����:e����µgnnq�ɗO�|��i�^yf��T� 3s�����c!?�1��V~�R
~r�8��@�B��[Q�ڃŌ}�.�6�tO�;KkT۬e�lr7�P{7�4�I��b�Iuu�p%�+�]_{�T;���he,��r�n�����co��\��D�.F"6שͺRtJ�͕k�I38m����U7~
W}�P�6��|l��}w���k.�n{o��W_?z�`s�m����b��Wt@�J�f�_�~M]�}�����X���8����d)yFsZ���D�<��B����
�'�lN%��Yd�>ԣ��(�J��T|�W��zx&�V�<4��g7�V�Ϋ�}�����.����6E�+�.���ֺN�}��l��M��?�j���D �!'
?{�Z|tT����{"��F՟��YA�qJ��<(Pr�)<c��Ǒ}�A��h�NҚd�8GP�8��S�i��1k!�(L6�^�=������={��������^]_��|�vЙ�����[Q�5m{�IK*%
���\N0���������'Q@jn�O�TF��,����nK��	^����������Ϳ�ۿ)Ma�����)
�L¾�I���k���+��s� ��7ߘ�FZ�]�(���GqQ�p��|,
��քcA�
*�tk�0�����l�sd�K�����Q�T$N-sS�o*��v������eh���ZL�zR���vk{�7��L�e�LK�R� �*�E�cŕ������4Ҿ��M�.�a��ȕ��f~&^��T���D�6@F��߼yc�݌?�V ���E�AV���ȟ_9I�p�d��-��H��H=�\�Ir��t�!U�b��[���j)=�urt��7�k��=b?ue1yO��9���Ź���rx=�yqv��8u�;�C;������
�@z��t�a���#�fm�l����5��(����̦y����Ќ��ƳG���1��;Y�^�Z2='�Ձ����|I�Sj��d�M,p?Kc����(%^AU?��\��$
� ���QdKCW�^_�#X�R�J�Tb��$(�o�Pt���I��c��
G�P�}��!�G���8�����3�V�J��|��
H�^)B�T4�/��/��9Eܷ �oA �OU���F�
Q+��$ȳnͦ��߿ǃ���̕��@?Uj���V���G_M�|(���t�Qk{������%E�����E��Ug���B��,(���� �����g�SNe��Udy�0d��d�CC�LH��
qȂЇ�I��׳��pH�%gq��,���ˎ�eY��?��H����������H�O	�,!p2�1��9�/�Ȭ���4��A�%G�����j�?o�BE(�+Q�r~*_���KKy�DP��)����X�~�)�0�yl0�r-Q��`e�b�{2^邃ȯ����LqB1@2p8х������)Z/J�'gӽ_�;��27�{r��{��䈱4�����j:c_k1���*Ǚ4?|8���˭g�pUd#��{F�Y_-v��Y+k�$3�O�Q_�	��x0.Sv|!-�'=a��9K��&Y.|%jȊCaA@�ly��	��)O1XTA�T�(Y��fA�U�*�� T�T��H5�,�����]�L��g���9��wq���ٓ˝͇��Y��tO�;������W��x�e�H&]7S��xRҺ�i�Selc�N3���!�L�5��Qܕ�'s����u������Fg�ǝE�^��9�	ȩX2e���I+.��6ȓdJ�<�L�"�B����d ���4����Y��!�Uq+zA���ӢZ�;)z��j�&LۘlJp袀���V�n>{�3�hQ+�D�A���ڍ�k���8��7�J&�Դ�8����T3�'g,�e�ٜ%Dy�<���;V�:!��ߎϻzA����?�=t��sw{�m{Ŗ��BzE� �*��
��c�G�0qB\	Dޥ[(��	ByD�� ���&��-�臘�7�4��4Q�����}�ᄪ���fDo�����S�a��������_���Շ[��b�b���s̑AݵD�_^XL2��g*��,��9��C1��V�h=�����(���MV~,��ս,0\��t�N{�z�NG���˹E�wj��g,��y!��j�Zsh�-��8���i��\�!/8��7�d0�Se� 
��Ń� y)`Q.�/|�I��_F*�M�������:�tϏ�����wϟ<ޘ�\��NR׌�	2}�v*Bcop3?���(����K�.I���E+��
φ ��<�	I7��N��P��Ic+�K�6N�z�9�;8�ܵaȎ��5GŔ���(�:tsmǯ�����9��q'o�]�1���R��d曃�OD
���+
�D�ED�~��HMf�>C����(.������}��;���/ݬ�3�f
]%��!������ʥ�Յ���G�$F��ݙ%reC�4fMGe�\x�%Ȥ.���3B�,��lGX�Z���c���������I���ջ���M��m�KW֯�=��72�n;@�ݓk�T�Sf�,���s<%~_�B� y�7YhEP2'����x��� �B��?�D
�X!,,-,���N�2�39��|g�=�dã\�3���z~�L��٤��d�}d��g�ܵv&[���]j��r����H7K�٬]vj��U���&�Q9;=?9{�ݻ����xy��V7�[n�NRRM���F(n�I�Ե*>r����-�o���σk�*��Y�'Į�A\E$�|� ��6Ҥ�q�V*� � ���{��hf=̂����D���=��ͫ��<�������E���擵�ӛ+t�9���*u�{�����&s#A���	�)i��I8�L�F�����ȴeV��sD�]F��ۮ�ٱ47�39]8�B|�����y�^������y����!�S9A[2$
�w�\f�����~,@?'N�OyA����&L?�!��''z�Z���v��A*n���U�����͕�dO�Xݴ����U�#ݎ���<����ȹlf��K�&������C��i���M ����H�Ff���f�@�cmb�b�m�N_���f��)A{���ݲ��ۋ�����>�Zc����R��hyeMFng���3XSL�YU��AMBW	�����D	��	?�ih&�K���WJ��Č�Q�ᙬ	���p%q�4N�g�|y�~���׹����$��{���s������ZǍ�yo�-�.�9�d�	t�=�߹p`�]�t<���X"&Fx��S�,u�'=h9��M�hwڴ�
�`������l�2������(�=uOq}�;�.�^��a�`my֟��P�����uM�DQjrMcKWɄ�f�����S�(��[?���|��9����YI���d�����l�=2%ҿ�<s��8��J�s���2�8�t�SW.﷽#i�[��ҍ�G��\�[8i�%�����"�� ]�2�eW.���@�0���>�5�N9K �{Su�\:�-��7fz���٥n�Ʌ76o�.{��W�7TI7I��/����3�;�� ,I7�*�9�1�����n
��o�#��	L�}IPh
�&Si�B%���>9|D�.2�rgw�Y��+Le��cʶ�!��,\:%B���{���֖0�B�Y��\z�+ܑ�R+��I<V����@������@��|��K�*E�x6�޹�7���xK2�&y���%�z6R���S�&��.��,���ڗV�@Ǟf�n7<�ɟ��_���nzv����IS�1y�c5Ãy9��O�'9�����"4�S(i���Eg�t� �-�Q��K��vɎ�+$����Lͺ�������K۫3�ĳ�+^���f�Kb���Ed�I�5q����^d懪g�X��
qֳ3>�광�ݵi���ʈ��Z�"kzG̸r Pe]��4����ݤʤ����^��LQC�*O���A��]��?���M�z=&w��<z��C����5!)���c�ɐ�Z,	���$Lh1���o�ܺ�2�/V}yJ�<
��E�I>qZ��JP�~
R}���W9�R���=j�[��g1�'̊%������zm	���ں#�fP�=����������L̇Gc�jf���I|�+���2@��b�$ފ���b|�4�8���(�ΔF�_6Ɂ�����iLf厹��>�ᬦ�ģ�bi L�49����,�T
�0,����B�A��䌃\��ʁ�Mi1���k�k��i������zck��ʦW�g��<��+��^��8��DU7�';�l�\9�G�M�|I�WN+��!��?6����H��0_�8��R*��8*�5AM\pH��p���iw���B$��̈́�mƜ_i�����ה�۷o5(��_���f�Q�=���Wfb��d0T9)�K���$Ø� .z����幅�v����>�Z��Z��V��2��#KW��)�3���
WZ��}u�SF��ِ>��6$��vz���������^����ۅ�����fy�2���N�����}�k���4�(�Yz2B�zA|��[e����5G��K�"
�%dh���U��5�}t����2L�("�$A�+���#N�!Xс/!%���g%
���s� �j+��]a����]���0���b�ɫ�J)]��6.��.-m��m��ٻ�>q6�0ل���:p7�`/PZ�V`�Zܿg>��Ӧ�����m��((�.%���(+6���?;ۯ�Gf��*����(B�X�T3��g���t�4�,!C�
�@�Bi׷���J'���P �B�i;O	Y*"F�[A�%��Ja|%����!X:���(Ed�T~< �5�	3RG���P�	���/5+��?L�"X�*���Y�c/����r��I�Қ�,R8ԕge�����:�N �����{�]ٔ��鳴J����2[-W�]k��b�8�7N�P��MG��P�Pê��_����1q���%BS�:��կ|��\Jn+:N0 }q���!(��˩�%QU+��sB�*�V��g�{��_Nfq"E��� |p8�WFx�2j4�"�p_q	PN}фØ���{���Z1��_�oA��<s�FG�FŚ"�z��&|@�J������?'O�$E�-�B�)ȝ Q����eQr��fQЗ#�JA�P	�(T�q"�J�\�8��JBBx���GJ}4���d���Ah����px����HR8ǃ%�`���G��s������nf�J�Oύ�����hx���������b�B���e秃8�w�U��;��IG��k�+�K�~ƨ��%���Ns��z�N굄9�\�]~�q��D[xZ�T��Wq��z�|}n�j�"CnG�v�5�YSb�]~kp��۲�%�t�m�7�`�͔H�M��b�q��Ze�"��3���J��'�M\�__앧2Ry���S�Bh�4�8#����9<u+���?sަ��#oEe���\�m��\�	z��ʃ|K[�E��֧�pm.�Ds�^Zmz���0���U.2���N�#ρ���>|8�w���bD���{~��#3K˫+�/���Ц��!i<��۠�r�+�U���?��G�Z&H!��x�a�o�_��)R���V->�WY	� )�}N.F򀊷����}f@���,g$���d�Rn3�o�t`���H�s�����.�dz���ֶm���J��qO9�c��`xyr����������o�9|�E�����������#fvRʆm� ���1)�ȅ�6���yM�-! N�Ɔ�/�V�W,8<$Ya�\�E��P�<���/q��@E��Lt ��RY�kIuSS�l����}9�p�p}7?5�C�+a����5Ub�C&zy�Mփ�c���$i�2��,U�Hڽ׶ߘc�?e�J��t"czmk7C5�|[�l��t���w?|�����ᷝ�c<,�,gղ}S܌XY_e+����(H�de���S��C\�>�JV��r�s�O�I
���E���*N�-��)x
[s���Ș�����eۡ;�����̀��j��4Vd����L&��$� z@E�\L��TR��*��T��Eg:c��q
�w�s�����7ޗv���I��;<�wK#ONXɼ���l>]bf�����]\E�4ǷD���Ȅ�|!�b�*�6ַl�X�N���/��^:(H�!K����#��P���c��zVrf�e�&l���eV�4�s�^>���-јA4M��R�0;��9��� �m��}�M�3��"��&�?�*��OAgi"��?���jGW�������ӽ�O>��p������������S�dQ�.�amF����r4�mI���XhQ>v9H�d�!8�q %R���'�gg���ܴW�x�Bj�4'
�,�X����jaZ��+���^F^9��\��z���hvVà���    IDAT�H��/�gl�ȑ��$�m,�@M� #"E�Ө;Q�0����`�WQ|
��`BG�-p=�����t����y���o��^���7s�[[r'�H0�T�O�"�W�ds"

��*�
3I7A��Z�D�O�'�< "RN�i�[@A
����0SQ�����M�{yp���fO�ݞ�_�!q=�w��T�#BR%�l\�f�+��#t��,8 �j$i�P��< ���m�b���&y)���&jM��0o��vή�.��u�~8�㻽7���1�1t1|�qR�M�"�X6ӷ��6����4ɐkz��L� ��U���@�/�Nc9B���*p�r� ��+�/<t�T�͢��^j�}�Jxt<3M�8+c3W�������٪+-^�9kaZ+��ݽ�-��i��K#�cL�R��e�6w�8���F���3�Q���$���h�s~ux|����οy�����E�Y���d�,�4d��B(I�,�� j�8���K���PB�.}��$)��)&�:9<�
e¯Pȑp�*W��>����N��G|����1]b�h�=�tiy�>�\	�$�]t7�}zzA�:(jDV%��,GZ��B�~��4[u�m�L��a�cJ\ՠ��.߂�����N��-ׁ��ay������i�����o��������E�b�ae���^��"
���Ύe����gF�T�(����$g0kT��3-�a �t������"�/�n�;c���a/�K��F�%���4u{���Ã}O�Zf_Dw7k��tƝS�۫[�n~�?L|�!�;Cw�D+)�#�LH�U�(���l��2��:Ģ����ց\}ђs�&�]br�T :��P��F�Ή%��������v�.~�?��G��su�r�9�E˝3�o��m���L���>iH��:"!�ׯ_���D��vp_�T���(%7<�T���+�T�O֣�TU��¡ϲ)G\h1�F��e��״�j�5��ј���T)[���n�N_���Y�bD��%��@X�m$hRMu�u��Y%��'3�ߖ�4c4OLN���T�d�l�\srr2<?{0voo���r�0�f�7=/j�j̵<7������������y���fR*'�CV�7a�}����w��8	�	��%(2,����D�_�X�>�s�|!ͥ)�^!�h�C�'P�!3rt�2�~�����9f���\�n�M쭻�ԃ4�� �����}�D4$[������
�]]Z�� �lq��BEK�'���� le1:+���i����&�YQ��x�ъi&���7��̕�y����?�뙗i��v����Ɇ�J���q�z�$qT�����y��D(H)6,��$V�ʓ6G�-�Ǜثh��J\� _�*ndԚ��$���p
����"�OZ���"���G۔���GAk��5���P���R��׿���v�gQ� 1��57�n|l���y*��JK�q��2�~b������otFha�� ��6Wi�Yph�gU�E�_�/V����9�gQ�(�FM��7�'���QÌ֓h�R���A,E�*���$M���Sgi���f-]:s��?�7�KV�g]��������l!����Q�%�Xy�-1!�\�ZV˲�1���1��H��K(�&̭�b�2���*w��� ���S���|��*����t�$N����l��۷o5�5l&>�$fr8���7(�"W��^��N�c>��/�@W2J��-~<��u�A`�����V�aߒ��p���խ�|�����F,��6�̑F��l��ͱ!���ɴ�$�DR��2V6W��X�hp밅�	ׇwg���ӫ��CwѤ��IH����S�� ��u�W�b@( ����P9-�-|��#Ъ �"�j��2��=FsR7�?n� >��l�%v
�Sm8�H��L�R�&"�rxP�
KP���.:�jN���\��3\�.�^�s;�Ig�}&���+[��<$E=X�.�9��{7sh�)����;�h}�����zd����/5ʌ{���>�B+hT�q=�0����N�4�f�t������,���h����.�_��g_w\p���ִ�/o׾������L�x����ɁC!4 ����)j�A%H��_}ED
�Ph��l��L� '�f��#z%*
?W���X��҄�5*eT��_� �[��B���/?W4��L* ����l%�A���#��\1,8ʕ+���~��G��F��)ʀU4UU������o�']"'�x$����^����:�E�e����fUU�U�Zn�������p&K��)�\����/��Rr<R�㋠\���2bL��`CZ�� ��� ?�e���(H�P_D?�Z��V�J�0��N���J�X�
,� ��	�p%�W��D/Q��_�U������"�m+����EP�$*��e��V: �zk-"�I�R��8'��/RADIݒ$R~2J�hVl���&K��Y'��^��r8�/4}��˗��^��BQ
�)h ~������� GD�nE@8�G,~��Þ�9p��)���<��
�\A�����'�d�!F�8g-{C���w^~���õ�3��>%iEcG�4^+��e��ȖU�u)�#)�z�:胇�^�Λ$�=��������L��� <L�~�?��s�"��o:��k��N������m�v�_��Z��^$̻��Y�=�<e��;so�#�9�m�Q]�e����<�Ob�g)�H×��8�O�͡�/�B�d�QNi�W4���E+"8��52W�zyu�%�*2ky=4�ru@.��`eddF=�"YW��Sޑ4��!���h�t�u9����@ɑ�{�ͳ�I�4&���..���6;�{�����ONOΌ�3η����͍&��dN�|[���-!�pД��B���[qK& 2S�9@�%����gYA*9D|���\E,���/��ї.q������:�v��㓳ӎ���+�f����j��t�2��x�`L�I#̤<�M�R�t���eF������ی�6�b� v���������w߼�����vO�g�:>�%M��
��G����òP���������9���\f�p�&� ~�
�7I~T���ʰ&�p���}9�̥Xt�#�¡�M��]���6l�eF��m"<�U`��� `�9�SU7��	Rt=��X6��)`I� ۢ]�5-�\ݸI�����ۃ�w�o�?�v��������xni��U^̆��ce�����u}��'Sܲ�?,x\\�%�(<dp��d��Ph���~���,�"���P_N(�}��ȑ�[lGߪ}��z]���Bg��o��Y�͌I� r���[���uX�b�^��m�*�V��c �:c�n�u֞�:�|`G��v�~�R�����!���Լ#u�N9s�$-��X��<Q��X�$>�R�Eʽɭt���@'4!�f�A����'7)_~QJ��%!sH	���		�3B��3���f?�7��1&�����9�f�:����3���L�a��TM.����1��T���l^a�mLQfjR���	��w���v��������7{�ߞ��g�73++[;�����S~�r���yY�
�+�D���2��r�Ph�*��K����+�~��*:�dX��/�/�L+����f�"�Oc�D4�2����:g���ca�o��Y�����^i�2gZD����%��3�r0�2'�qVQg�1Qk�����0/./N�޽z���}���v��_�=�u�^^�y�@I�Y�$y)�K>%�
�Y?�H�����D�
�j��M��A�rb!S���ϼ�W���|�c[Ѡ�#���)��r��^s�C5y3��.�U_26'��\�FzL$u&�� �2ʎ>�<�O��Sa�4���C�)�L�լ��0';ݟ_�O.�}8������pp�sҖ��Х;�\ȯ�p�K��/�*_�|���� 9�p �).L�x?�����˥0Z'����_�}Q��@�O��L�<~bI,hH��|�(v��t���,^��CŷD��ip���'Rz񦮵��/4V�Q4��+�Ƞ��ø>W�	�����R4tG�k�ͧ#4ޟv�{G�?���;$��#:�ђ6�KIБD�<rQR�,r � M(� ��	⧂����+��&"E�7��&IB�� �I/b/ds׃����>ݠ�
OόM#\��h�p�o��GT1�a�a+"��
�P�r�/��AR��ld�)s�2fuSe�ae�V���ņ���
ҟT⼺���v\k���W��^�9y��A�njxk
j=Ϗm9I�Z�V��0����큖q�-ɐ@yJn����N�����J��	2W��'��۴*�&�7��n�D]㯢����̲�*���o`�"d�G+"��'�{�s��rN-Kn9Il�.�j�ҜԴ0cag̠ظ�bb��i���8j��s+笉b��x��NU��gQ�q��#�pw=\t/�;���·n��?����5��W���Ro��8ϟ?���.��'�MȲϑ�����lfZ���ID���y
X~����>���pJ^)�Up�BE)8J��f!��Mg�Ye��S^2��,/�6J26YG;yJ9R��YpW�rKg�-I�e֔�j�|5�\�TȎ9[�5�ƚ���J�2j�奓bދ�w;#�5�?v��W���k�-Z�X���a�ٙ幥͗?�������5w	d��5pJ����}6bF��	\�X�)I�O����B�08W
�a���W�������f-*��X��H�Ў���^�\[�X'�����Q�[�&�{WC��-�*��?M	�����ue��m駊���Q��x��F��Ҋ���B���*f
Zc5�+ ��`�6��ܩS.��_�/��q����=^V`WV=s�������sFY��vji|�����ӯ_~�l{�8���G#��O��Jڿ��oY#	C)�j�����[���9�>���p���|��
&���-􋸟L��U����s���9��qZ�iؓǛ�Cml�>�����������#&9�2��\���FU�OC+P�teel�Wr��h8|�UV�_��1� ��D�4YE�o�)J^�ė�Ɓ�����:��1�J\L��ږӭY!�PԴ0Rf���r�p�a�OA�[[HXBN�N��NBR�Oԕ�S:!6X�gH���݌o��x��Q�]�Z��w�Z�����i,T�DW�FM�$�D�OUO�ۈ7\��ҐBä��,��*i�W(�PqA*!�"�g���@1��鋎�y��SO�� �
���"b�������C��������Q~�%���E��$D#M_�r^_D
�/yp߰nb֌[9Ӌ�K?��v��國��H���;7���kj�/�����TәQz)�����xy��e��%*����./�K�+#�i��T�]��[?�Ø,�r��0!⭂ K��Uh�UA�˒�b�%���Lq�0KP�j����d@��ě7o��B@&J�����x��Ok!jRp\,�]�$.��G�!@�����˿��Z:B_t?)%��7�{=�P�ޫW��6V�6D��<z��T����Uǅ���s�WL���m
$տ81�::�^���KkCw��gf��n��y�m�DA�"y��¥>�P����Gn��f�L�S��g}{}������E���0��?7�V"[�dYI)����>'�#|A��B	-��#Hr�B2~6�S芕+�U��A�Ƿp�%�T��4
r2�R)
~J���Q��� 9h~B�d1,9Ȋ~��0!`�É �B��2���)���BF��,�F��%b1 LԸ�.@��۷o� ��_��_�gG�@f:,��L���$��$����|�6�<RA��DG#��sR��w�}�>�-+�`-�� �����ϕM͌��/!�V2�!�
�"��m�T��T/�G,�
�����*���HE�2�%e�Y2�� �8���#�UF�+	Kw��@V/��(:�2e��#�����W"rT:�Z!�����P�P���9)S?���+"�_t��?�;�
�)БY�ʸ\���dY�_~)H)�������씦�E��"X
Ft
��O�`��EM�����D!�(p�y8��� :�c�&(���'x�9���肪X��X&�Ok�x��e��dI����<�BJ҈�I���7�q�9��g�ڷdp�(z!�HE�5h<����B���Z[]������g����-N���ۿnlG�봁����Y�˦e�i�pjin���`;I�!�Gݳ�~ݿ]�Y�Z��s[��?�3a�����d����؄=|a��b��T�˗m�N7?=?�蹐�Y\͌����ⱻ���Q3��/so������k�-�~��VK���Y�U�[��	�X�)�x�ِ3�[?��8?U6RyĿ��$́p~��T� �W�Cٍ� R���N<�olY9~�h����K1Ks�c3	K.�1�׫��䝬����vNk{l3�h��9t+x:��*@���G=���ONϼT���ء���ڱ���2u���xD�/����%;~Vv�A�� r ���?AqBY�𳂠�P�/a"��2Dp*�����{�:������žbi*l��=8��9z�����O����+ox���W�D���.��V��n�>��d?,<�E�ڌ�\��f ox�17׀�Ҩ���w~r�9b	z{gG�A�j~p�2�`��ې��o���Y�֥aǰ�s�Dt%�
�;��4J\�}@���	����O�@P+:�
�%����JA\�K�0E/j�y�S	!R�����-�	򔛑��ð�}8�^����>y���G�[K[�Y�Y�M彾2�� 1�'����SSt9q�[gKr�$e�z�*3��c�gv���G������Y���i�C�,��;����S�sŹ/j�ӗ�d<BlN'��"��}����''�%1~�����St���Uv��9�&2�bQ�T��
�A\ZŞ���3S���J�m�����?z�d�у����[�%v�����h^K��S�XN$�j��tD�v��J�r��Og� 6���q��l��^�ܩ��Ӌ�K��=j����g= 7��@�dg���&�+��.�_�WI��D���ω6�J�(`����,�\!�[�/�' �PR����pp���B�K���~u�etL�!�����Z/_<��X�쳭���U���Ș�QE�Qk.�:�*�h<���[�ÿ��lH�61�����Iw�[��{����y�޹�l�w]=�s����:�k�����)/G�ܠ`��eV��l˔���Kh�6� ��k�Q�ܷO��o�خUBK�%����Q�Sq�)��|�"[�� ��R.��\!�f{W���~��w��qv>yd����mc�������_^XΪ{n�t�C
N*JY0o|Hy�`��g��B�-�J�.��T����L[�.z��N>ؔ2<0Q>��Y�^Yz��av������4�.	5W"��#iT��K<4N�H�mc�OAHqrQ�.�EA�W,��w�
�At�Ed����7�� }�p��5ӫzw�7��t;�'�<~��pmy}a�`SV��%KO>�!�Qzjmn�ٱX�X�膙B�jf�T�B�z���v�F�v�uSH�'���ڋ�'��GǪ���i��$��+K�+kُ";ż�l�� ����/��b��$�"�~r~��&+h\Ax�q�f�B�E��
x�ε���O�2h� �`u˾;� ´����x�9���Q���m�T�j�EN[�5YMK�&=�\��k)�;�=�)�X�ir�Db� `+�f�XD�R,C��C$Fg����N���c���ǯ�3��Ы��)'EN�!T�d�*ZɤԌD$�?dN,=�B�C��J�P_hL� @C38!v��J��2�xJ��FKˏ_�|�����`���e+(7��clĜ��̵��Nי������E������暋H�\
�(K��lo�y�\�B��O_�ƛ�M#k�9�>|Fɱ`�E.t�~nÊJW��ҝ��u/�O���C<ur����ɻ�
М�����ҚSV�l�P=ba�    IDAT%3kpjV�H��(H��ȧ�؋L[- +#n#z�_M!1����� BEAd'~8�PoC`ń���U��*�����˟�����Y�bS�4���4O��'�s㫕�ۧ/2	`�G���մl�t (��J,�Vَ��]��՗l��3�����jm���dB9��[��
����6����٨;�^�:�����Eގ�rHJ?pm#w9J32�Xʱ'�@����r'���&�Q�:��ծ�k�yp���	��%vqK��j��}�CK*R,N�)��p8�hp��@����((���]��r{��P��r��8�����H�ぎv��!C��&�s�sٌq�:�+-�k2L���3%i�d������85�q0����u
6�; {z�;9�]�}����������"%Ϛ�����������/���^[ʝ�i �3��r�@M�:�e��P�V�(H�+"��,���$�oLA�d(G�W\ #@ܿz5���uʤ�p�����^Go��wu��x{g�wֽ�8�a�D�o��ؓ�����լS��0既Y	�o��$	�R�	�m�J�`���حF�Z��uvƺdW\ZжaK0�7:�un�h�;� �u�7��Uol�u<�9빽f�9�Y�����vϮ�|���/o��:+��������O6l�U��6�4!p�,��=) ]�"��<�[�R
%F�DG\@R�-HT��~&w��(4GC�?�<��_� ����_�� �U�֓*0��9��kiqVK��wo߽w�v��l����Rd�OZ�c�u$b�J4M+�qUЄI
�!������?���a�M� ��XG88l��_\B8'vK2%z�>Lb!�2��Rd�A����<媿'.����L|*;������b���X�l��޺ecn<�}������W�i',YZ��g�5�#���Ѽ�N �Yui�3�����l�B�_�_x ୂ�����/E_p�y��3y���u1��\�9d�42�֌��m�\��D)Q+#F�����a���2��<������t����4w*9�[��9��J��˵�a�p 2U6�l땻s�Z�y)%�ݜ�`��Ilw�J�.��ϱ���v����4��ei��z�,��V�=�_���Ǉ��X���N�ʎ�q�HX��i���O_A�A�P��T���
"+r���u�*#�f�9@~@*R�.j�*9t\]*5��&�u�	)*VT�HXtŉ=_u�hJ?5��o������+{s�����lgvQ��ɑ�!����B$cފ���:�t뫋���w�dd@��֏��A���M-��]/���v4
yǹ9-���4H�St��e����gW��F��n�t���iIo���ˣ�?�_���!-.�=	���0!�h�G�2�� 9~���/��DG��26+"8O�$FB���( ��d�DY���+J�*��8ĉ�1N"~
��DDM� ,!(����Eh�<J2G �*�C�px
���ĭPdѧN�O�~��A������'x)���բ��2���Q{q�&_��/E�H��/H8R���Y�.S�g"
hhB�ӗb��� ����O�9I��S�� �f5?d+��%��(QQǭ�X���+���aF�Ã7��*Lh�����_�2��(�JH*��V��?�Tȁ�K�H��ƣeų�.
d�q���G,	���^?Q���/q�YV�IC�h%N��R��2 >�Pމ�� j~���9�Ib�F����EP�%�U^tD��=�(����?�C��&JҤ
Yޕ/��vqS"� �ҽ�GB�T|�E�'w��(�������m�����-� d�M<��3����R�� y,�	-�K�@ C���R�+K�B�7�X�X�������Wǿ�����K���f��$5��MH�<#v�L0��ѕ�s����ъ�d���=$m���n��Q�LI!�b&�~�U6�,�*~r���� (:�H���x76˻�1����\'�<orњdC��܍��ܛ5��k��nW�V.��Ф��|t&�!'�3ِ;e8�7p��b��\p����s���[���I?�,�a���"w�Y�'%�N��if���{���gݓ}k��>��U63 �I�>�v͕S�dej6W	��,��2��sp��^�l�웺�;\�Q��巛pK��X��I�8<�
�2�4�A�m~����gy@D�q?KVE�mm�/"��ₐ��D}�J���":��'q��'|����?�Pq����)�n��~ �'3���k��F�ֶw6	�imu�QΥyw����i��6w�nd�+C!��G���Av���m����t]_ѵU��l�J����?s5�t������Y��� �n]S�󳄃l�U�ȼ�\Ic"��VJP�~��D������%:��ҁÇP�MVQ�,L��0�/�J��+L�"m�x�y�vvNGþ'/v߯om��l>�Y�y�p��|Y~�%�u���a� 6Yt��z*6�i��4��Q0�퐱k�/�j�Z?�:Juq}f��~��E}��D��hu�Qk�����d"�����H�nJ�8?"�<�o��S!+YNPQ�_�\	�JD*�����IB 8�\?97W1�8�,�cfz�OO�=<��m.>���~��p{�:���,����K-J��m�ӿ����r!�����(���{$�J_�V��q��s~<:!��SWS�������>�IX(s�__�tp�Ϗ���T�y��	N��� ��Z�p�">�s8�_d���b Ώe[�E)j����NE������J�loKl�9}�����N{�L�;ѓ�df2�\��T�TK��n��þ���z?����w<��v��*��-�$�����Ky�
�s��d<�=�-���n��=�yh�ޒۆoh�e_�ɞ�;��Y4�֗��¶�B͚����{3N��&��'�Q����s�ۧ��v}�v�h�p~տ]�p��_�~qY�=�,��YW���H%Ȣ3��>�&����|�j~���Ib@���Ŝ�[�8:Oqp+?��� "����g��[��N��j�Z߾�6�z�i�����/�;�n��$��i8}�٫��w���"�vY�lo��/��'N�B-��A]��	�8_�^�;��廷�����j�/o�NZ-�����2�!1O�ҌR���6����o�Y,�)�(@0&�)ūL[Y|-Y�E:��Gr��$���K˕&N��T�%�}dN�cm���{�l�l?v������l�b�����.�fu�u�����:T��N_O��ZY1�kn]�TW��m�#���?Wg�-��|pw�=�{>�����UFHl�p
��Ҵb��

�<����"���C%�Aq�=�E0�����M"��0��/��M�huN0i�|[��gsbd	�=m���Lܢ�b��o_~��Ӈ��5U�Ǧ��Y�i�t�� �n�p������Z��@��-��������p��L>�]rS��ؖoy���۽�ׇ�7������`4�t��.�>�(���PH�L	��v�s�Lru��ej��Ҩ膏� �R�S_�{��5%�Tqxk.WT�*&�U����bţ�����������7㳉����Y��X`�3>�OT��k�''>��1Z�3ZU=�I��oR�I i-�N��ɥZoP;j_TMP�2LEꒂw�J�+��s�u��o��^��.��=:��;��vAj�
ЃM���!���z��e�%�O��2������V���U�KL�r│�N�/^H(������tP���R�Rc96���H�68>��s5�?��_���5�[�|��Ǘ?�8�9�B�jaaz�sೲ*e��f�������7�צ>lǕ���T��MS1E��[ڞZ����
쥰}@��2�z��Y��.e���ql���������ba|�|�ٸ�Xh{�vg������v_c�q��5�Rs��vY?�%�D�)��r��r�f��Ă\��L8B����(�!L�/��� �H\
G%W��H�>Ǥ l%0LM��4L[��0gbC��z��{�m����;�í;���@��.� �Ț��T���1����*b犕�o~x�+o56�2B���P�����e�\n��fe��˫ׄ�O-��U���������mo���l5mm0`:��)�nq
qqam{��o���_?x����vݗ�5X*��ۉ9���řb&�����?��qQU�VlIW<8�H>���:�b�B�Z�Y~&Y������ꊺ��嫛�};%���_�ۗ�:K��>*{��6���Z��X�qpm���?�=���v�*/���J;��?�YW%��e(#� ��]���SCrW\;�	�����մ�Ϻ���Z��oL{��.O'{N?�X���3-��=6󡽅N�Ƌ�U�D>�����o��o��X58�y���x�o3���O���i���<MB�.]4�T�y�D�8��&¤�h;8HC  ��\B��1ui'��?��uȚP�ͽ��6���޽���|n�A�&p�.��p,��Pc�~���榕�sr�ɱ� ��Đ�KjM�.��f�U��t^��/��Q3ChRQW��3V��g�:��<:h�\�0�0���?��8l��T�OZ��)ǵ���j�1����1��c/�#�&�@O��ˋ����������5�U�q��vݱm�f	U�j�Vgj_���W�ę�GUBl��:	p��F���Y0Y�� HZ�8l��!�:�ׯ_�����8c����w�,:[刜������aW�|������ vb�E'� �G@q����I$^6�_n�I�T��a�����]��.�Z6�ʏbݩd�bc�`�>S�����Y����9�����?��W/��y9=��>Yٛ��Ř�vI�[���v�֛!��*4��/nM� =RC�G�!�Q< ���Q)'��F<\��ͤ�׊��_i�A(?�A�-Ke���W��Z��$�D�X���t��_�~i��}��ճgϞ?�U(Pri����f�� cHLP15�������_mu��ޠ*��!":a49>=������f��n/�:'ǵ����Gߦ:?]�e�*M�/�#k����'3��5���Bu��X+�:(V�6�W�]��ke�P�ݦ�Y���(n�h�@�8�! ��n���:�{T��</P�Y<�	Wj�X>�cMh(աc�b�b�tj/��h�RjB�p �\141xi���3��)>�)̣,�����BTb;�<J��
��x�\�ZD4��!���H��ɽ�ɒ�v����O�@s՞	���q�JmWE�JU�gZ�L�����&�u�ik�����@������B@%Ms!�f���q�Yчz��C(W�ӏʟ���C=��}".�X�Q��[�c5 �����7�_1��
�(I%�8�dIʍc�Ϭ���W��>p@�J���a�M���?�9t��|��,i	n�-*�y$n�k�Q, `���GO�8{$g8D㓞n�]��<bE4&�/�'�O�MߥV��r5 {d8>JP̫
!�~����_�5��G�
��_���Kh�D��lt�r33p��P(��l�Y�`��M
=�!���@Br�0YR���?�j
���������x��^}��/Ю��Ko��)��uo�o�R��W��e4��Z�$���s5>5��*nt=��|���e[SUL%�pKJ<�XԖ` �f�Ǯ�#�2����^o��W;����[��ڧ�:���/n,yk����l����d������7�¬%Ɋ�`,���J�ݵ�(ږ�>����̏��I)�P �d��8�$P�>V�D��X��j&Z��}*����\6Rk=K���>ܗ�e��gxtz���Z�$	[!*���Y�P5vK>��9tf�15ce��t��m\��6�WM��t�$4��L�傴��1hb�b1+$)G<��ပt�@"Z�p�y���ͳ��QVdp7mS�Ȣ����Х٥���W��GǪ�r�z}��s��!��^��ኝ(�m��-��3;��p���Ksd�_�_��<���G�GW7�'�^j K&f��EN�."������]�@O꥓��9����~ZydAPU8\:��N9�#D4ޖ3��)��Ure��أ�S�4Bi|$��mhQ�E6�wkg�͢	CǛnwv?�m�����0��K'V�M76|�aqݧ]IXvZ��A5�Eps�3�x���'G�������y]~r�|�|f?����l�����M�����y�޵@[O	�HL�x	�,��d�~���+��	MT�#B1n�˒�3�?TA����ɕ 7ܐ��
s��	�!�8���I��;R.��;�ÑA��@�_q�|_;r؍8�7f�|]��q�Y7��c;�K�Z֎�����|l$`+��W{G\\�0����s�ڄ�b�ʅ[n(r�dݠ5�c��Mq��eNK�UC�?��ѣ��x8pi&�NH�0Y"��?��
�a.�9	�ґ�r�p �'@���*�����G8`�1l��o�X8\7���={�����������{��m�1�X���#�I�k^��{ͱAB![x0�o��3�g�
m�9:?�;>��}�tz���W.tW�`��^�E}>FzRas%bf����C���.	V�'?0�b~h�!#�g �P�	
<^�M�i�GzD�	(��'����8���d��U�UZ���rr���K��3�^]魍nG樖��;Lyk3�巁�d����Sej!_o�r�a���k�����N���Ã����������D�����:~eg���8V�7�a��T`�`��@mp��Y{�H�QZ5� �MZV�&!H�xr�p �@�#'(���DT�Im@�Ů�K�% �l����fB�~�ˋ������͗�w�Q�1s�����u/�2�[��fnk�03&�!̩`!���f�������S�^,�Z�����r�4ݪ~2G�S��	Xe���4u�c����<����|	Y��(K:@��i7���!D��80��*��!���(�R[�ԍ�Jߡ���#�燧������g��=��\�����A_}�԰���a��\�jS�*v.B%�� AU赟�GL]z�����x���۽�����&�c+�օj*�v��e��?4Tׯ[�[�[�jN����&�� 4���-���i>
g�B� K��J�'!����äs��U���U�H��Q��Ng���~g�������g��?^������jvQw�(�ђ��UɃ����]���ȭ�>j�f��9�Yצ���X��H�w�[��bU�������o�)�i/��*��/��_��~�QMteo;j@���>Yba�^�&�G��?y��2ۦ��M�a�b�����FL:O�3��{g�2�Js)^�/.C��%�{���q�DL����[���[s��x\@�S��lO�G�
���7�߹8����Ҿ��I;�if���ể�~�1v�F�յ�X;���*=�J�G�%����W�>�ڟR��yh����JT��&D!���>�}�tz��}�w8v�hl���ۃ��;��u���:�U=7+[� ����v��t�!(Y�L�C$�:��|�������iJOh�/���t�.&���g��� �҉���f�\ݖW��|�B��(�?��?����^�z���xe�đ)Z��.�9��X�{��{��^r"y��~�ˣ:⪄���&^.^}�1�5���\k��#
]�2��ё��Yk���^-n.N�g'�����3��/OǓc�n�]7����h��[1#�@�c)V�Mܿ��g_?��?�w�Π�q���j"
����u5~^�xa��#��UF�?�R�9�q�ʌD���Q
�ʎ�o}�Q�+a6�;V=�����a6�ټ{ϝ����l����.j���j�羱��r�}ǇY�7�}"�DNt�    IDAT��n*=�������&LT,5d?`�P��n����}XE3���eA-<�-�Pk�^]�lN�<q�zz~j��x����酁έuх�����P�ݹ�w�&�Ս���|�{�������6�i��E�����3:
o�Or\-�L�v������ax��G��Ӹ|��d���(_A !�#�'�BR�*T��u��z�����K�����|����s5��P]Q�,�y#oF.�d>�jH�3<&`���5��	 �K*s��I�?M��%LB"�a��D�6��F��g�[�p���ռP@H�:��8!�Bn�$K'5�__Ad�l!�&0و�t �@U�,l���.�14�z��'>����}zxpsq�����_�����������չ]+��x�i��7ԯ�`	�����#f��!�J��
�4MX�4p��0��e�7@����K�E�@4*$)J����f����jh5��>����}а�;����@����X�%�nҘ�'�����:s��!��-Ռ������Z$jm)Gfg�S��x�?��t����u��ϑe|���G������z���~���V�n-Z꘸���:J?��W�ڀ3뼏��L&:1幘[ �#_k	�H	A��@�����B?�op8�Ҽ
YB�H����k�B����V*ȵF��!4!?�� ���ԐN2�Bs��#h~o��O���@"�Q�C��-�M������y��g��m|��3��V:�������ɑ��/vvN<�U��z�� }��ݎ� #�%�kܧ#4}�-�|�R[������_^��P3�xz~(�P�D�{��ɠ{����_U׌���R����W�J��[2	N��R��"�&�u����h0�$�|�0���+�Rp�b(V^�K��`j�4Z$�b���HG%�DB.ŨM�h��YyD3�Q�Q%4oLp�� ��#oO��)�FuC�DEa�؂{D�9'�Qs�Ns +���4�s�䪐�(�~�ߐ���50�G�($�@"��
�G��1S=����tlT.��v&`Hs@$�=�*<ȕ%�Q`���Ϸ���4�ԓ �+p����h��L� �,�G�e*-�H�H����ǘI���d���r="`Bh�Ne�β���!*q/%���PPE�d��A.|�)���D�B ��<FZ�	<�����ȃL�\*�D���@`>P�H�:��MON� *���[��F+�4�V���]�_}�BF�@
��b��J!���_>	rU6�!>)�c#q��0�G�GV��TI˕���\�&�pN����k���~+X�������am��,���>S��n�u��W��U��������,�7�s�	m��n���)V"�J�{O�ҪR�^©D1u,pVH3�4�XZ�A.*� p�N+O^uzf:.�1�\Z0C�C���x��x|�21G������p�����p}�_�v�s�'S���2������RU�) �t4��>ba�07Fm18͑$sno#��!�	p�%L�8�'aJc%�}��o�~��-{�t��I���MoO�o��}��P����菉9_��~�6F3���,�m����^M��ƅ=i�N�ŀ���cG?�#!$�\<�he%�Y�(H��(q�ŀ�ID"4j�x�<�Be ˕(���� � n�l}�eyea�$�{�:�3\��\�;S��5,������"�cX���U�G����595��L/�NO�e��Q"��if�$��|��<�0���|bWLjq����K��VU� �	qmi�c���|	������$~���r���$�P�8���M���!� � ܄hB��+T͜���b��B^��u�ww�!G��VM�<����{v���t��Yi��`2�$�eo�Ǉ&Q�����E�qws�(m��N�������o7�~c��a9
V�g����&�I[э�,�$��D�!�G�h�{Y
�� ���(-̤��a�!OL"�G�$�,�\�d�\�᱌��[��À��x��p4�N_�1�(xc}�9�/����ھ�Q�ϼj�$����*����/�a�SIN�X������><z�{&h��>�?�m-�}��n�+�[Ũ�	��f�4AV�!heW[��{/���I���'�0�&H�p��y��a'��DoĖ��B@Ҙ�HFЅ*d��lvf���ͻkkNClm�6�F�A�M�i�~ݘ:[_�u�̶3
.M�٫��Y������:9u�����v�&7��I+fl��m77�X��ߛ��Tn�í�Ֆ�~X�&LUV3G���qf|+F�]�*'��C((i���R�I���i	�QE4m�*Ga�Q�E��p5E[UuU�2�jz|t�B�?�4�3�xgk�+�@�����T���s,��4}��,8�\ǹd��D1><:u	ꑝ�Fn�-89a����!f�	t�9&�lm��#n:�6�*�'[�@]Ka?)��KVB���>y0�q\䑻bEJ�8��������0M�4�]="O"A��bA#H.�~�	Y����p���w�W��sw}u8[9��o\�9Z6c�h��|�35�dm�Ĵ�	G&@�v����;G�Ϧ��5}�+��I��N3�������5�ӛ]�Jc�q�-�dC�,+�)�[�@�@Y���
2�,�0�ȕ�O$�LD�`5�'N ��V"8�C��1�@ W_!ͯa�8��n��. ��\�����#!����6r���V�2se��G�~�L��\ƭ�����,�ݛ�ɇ�u���;8�\�\�����w��؍��+�W��e��e�i,�:��DI�5�`Q�u�5��C��c�����pZӘ�3n�{�;�q�O~�"+�RB�xOwa��Z�VSRCdI{3�L��
Q��փ:#����`����������S�^s��MW
����(ӓ����ν����w�a3�[]����溅	G�j#��Yo$d�㵇(KhuId]�^og4�]��y[�\m��+O�zz29:p��S}٠L���"5�yuG'gl�*�����_����<d����ُ6�R�1��TN/����o���q�zH���FYūy$i$ye�9��o�+_����&9qo�
@�~�{�fώN��Nt�n��h���:s�?��9z�f�h�
�ݻ�#_�[�vk��z&XyU�6t���0���c�����v^�5g�uJ��	�*����O���6�����5q�f=���
��f��P���/�^U�oM[?iK�V7e�4���$����?����˿��7�82Pm<�K�K�6u�'�:�
� Y�� � �`�R���[ņ 	�KS\���O�Ik�V4��3�߫}9���X�o��V͟����v�x��jm2�Pa���
��0P��fQ���I�p5��ѫÞ��+s��p�]��>�mI����������pU+�a���	��ͺ{��ov����n�4j�u���Ϩ!�XAM�p>Q�_�;�8�*b���4.���S(����7>�[�To���k][��
> Bζ�ҋ�������_�F�����ׯ~��M�-������F�����ޱ/=Ց;�bl}�u�B#ɾ�p;��ۉ�R���}�[\���/��u�u�5+7fY���OAy�g�_Л����v?���f<;8�?�'�K+C�:�Q�Zm��۝��c�V��ٗw=���G[���ֲm��:����(�Cu�*�Z!+~V{�g���0*nO����� �����^>x ��9p$j�ty��	d��˝˅�T6�"��W��?��D����զ�&{�;?<3!<�b�PM�43%P#�:e�	� i��$�	��"M.����2�� �o���� ��G���/={	ҷ�z���ӧO%��%L�d!�|�b�>q����C#E� @ֹQ����,@5�t%��!��\.4ZR?뱅��
>B�42�U]ؕv}�:\Y��1Z�^�wl,�y��~���GW��UW�VV/͟���u�W�I_�jlu��	M�W��+�� ��y	IJ!.���_,����� 7	���: H��i�� ��	�xI�*AnĪ����lS�|�q�TU���(��AH� P-��!,��*�cD֡����c�H�(���e�Wj[.��I�VB����G�\m�5�:h�!ZU�.3U��W�ϟ�g�Cx?6h9,��T���t۟L�hE:���Xi��[ �8�9Iǭ���3<�t��D<or��*�8�?-�����q���Q�D?0ЄĚ�f`]���L7+~Tp���*w��A��#�o��o��p�h��=
�j���s�k���>mv�ޟ���<SE�~��ŕn������]?�J����t�q�A����s��|�k�N���?�+,��Z�7E�����d��Lm0/>�����j�[8-ܟ���}f3)=�Q��j�m�y�Í�R(�˗���/~��_�9���&� �����}J(��b��M2)��P͝	a.%��cD�y��AH���ꀬp�Hn�H�p�*������\�2 1��F|!��l��:A��.Y�@<&-[�iT'u����}��h�&�������D��
E������ǈ�`>b���A�G+��fH��!Y��t\��§�H����*���6�qҔ� �Z.�ɊW�)I�VII���ҊPj��3�F+>�����:�|���Jj,L��;���=��K\ʔՔ�O�N
�̗��(#�u��şJ�C������Aq˂�9A�pp�����r��A$M%���H��G.��s�X�Dmf*Al�A����;����ϟ={F
#��4d�Ϊ�S�QO~��_���F�Ǌp��	�� sl\�c�
<��y�FYh)Vv.,�!�IY32%�%0��GAZL4Z1� D�Q��|B�X��)I=J�#��V:d顬�V7��VV��ݼ��z�j�5C+0^>��f��G3�ww��a��2�_v��5i3���~}�J���qWШ34��Jk��*KXg�O�J��E����i���� ���A0��S�����lV�#���'�G��w����[[Do:v���'5PZX\���?��=��^�zy���m���/�G���&�$&+�LrBIoJU�V�tt�����%�]6b�\1d�1\��)�-����[�HҚl�^]Y��j^������=y�:�6��_?�m��qE1-)mȑjF��L[��ע���&w	��5P�t�6s�6������(��D"8XID�8v��Vc%�b�mH�Ȋ�ɥ1��!C���sDKÌ\haV��!%eŐ�$��݇�
�*x���F���M�S������Nd��̻'.4v��5���j�*rM{]^�����F����9l�����rT?7���m����we��֘jp�"��/Hs@�0U�/.��;�c�d�tI�4H�44AnT 	<��9� x��9�u�4	�0�_���T.j�Jqԣ�b]E�GB�_�mNP���y{q�ý���������lӲ��+s����;w������%�'j�����I5��3t>kh	���N֋$F��.����{	h�9�<&K���gTS� �0��QLLVD���� ���L��x��y߂�а� �4rb���㧍�O׆��_����Ý�)#��Iك�q�rq}��J׉�?|vx���L~���ٺ�g�&��B�kR�o/n]-;�=_n�!���ʰf	���z��ש	�y�\���Za4o�^���uWb�-A: QB-b��� �Q�`&����ӦG�0|P������e懰9�j��I�pC"� ���(���.ZYh	���$���\�TdYs;�hT�o�uՠ�4��� 7՚6?���[+���w�ۨcg���+=�wXgn/�Y\�,g����H����+W�����!@sX�T��)�F	љ��'a�pM\v��.����4�<����!$����\ �+!�A��q���Ѧ ��d�OzA�CQ�~�������n�c/���7�'\q�7&�k��5d�Ynk�n�I��5������*�C�zW�C��e�ZlګAi�Ej;�,g���{Wq׾菿\1�+HgT�o���斸�Q5`BCH��&�ʹ"�&��p�Xݢ@�z� 8�@�_B ��Z
�����VFr8ƅ���*T٬�c�����ԫ������ꚛ#\��[�&3�6�/{7��=�bJ�mʓ�j�;c;��	/&�}8�x�?޷_��}f��\#n��.K��E�2���I�`�x��y�!TX�"18�?�3�01g2���gP%�\���M	�8��,
��VRb���Q��0<�]�:8�(p�0q9����]
g���E�>�ss����G�d��训�o��[��-�P��vc됵
Ou��^���j�>;�j��۫3w������#\e휱OJ\��|�v|`��+((��Ћ8|��B�=�0�3��S�de���˟s?0�� r��'�8���J�8�UdH�ރ,g���֪��	�Q����(�x�������po��4;x������.m�����d��@'�q�;�����e�Or}k}����{w���kK�����ʰ�q÷�I����]�O���G����t�S���Y̟��'Rwa�!{��R�&���i�4Z�����ɓ'�S��
8	%�SӞ;�ۨ�@G�c��K���J�E�,��߲$R��%�,���w^D��	m��B�CЈ�>����/ Ƚ��/'��k�}�����G��.��3&��L'����|�g�wd�~�]sK�ƚ�b�΀[?��g�F���%N��۪�kr����6��fs�;��G�>��6|�k�'�6�_M{�sn7{��`*���$DM����62�uLK�C�=�U�lpwo��B<� p��FAB��+�%8� I�Ws��b����)�n��m��@(xl���wi��a�Z�}�Զ�^NάĚ��y��F|��õ���h�#�GX����sѯ$�h�N�{��i��?]�9�ǏK.�'��h��&s�՟���C)V꜉[��W��j�yf�Yl0R��=�?��7�~��-^F�&�u����s�Մu�:��	2����k�<ϓ���7�������+��XV��n�y��8�σ�VV�j8������f��Ty[��������k
ݩ�k�f�Y���m:���&�L;���5���d��|ͧj�0���Zq�w(?����;�]�(��޵/��]�8�iV��#D�1z���O���!q4�HcꃲvT�����Ͽ��ν�.i�������R�^�A�b5�T�8�8�JV��4���韥y��(���G��CH�H�b,Z�lV�e�!��i	�4��T� d"昲�U�x$�G鈷�%�{�R�N��/޾{s������>/�*�r���2�:�"�9��Dh�#�P@1�J%M�yf	V�4�V.&�9�#� P��g�g�-��*z<I�k����j��}�U�hp�8Y�Ԃ,Ӥ��շ(kU�*���R�!P�)H����O	‭�Z3�o����;��m�M��t�������������ڊ�Tۊi�y5�w.'���'��;�\m�,�S@"��6��>���2%��dQ\�GhA���"�k����
�\�\�=jp82�99��)qgBD%�}��%�O�>�e �WA�������
#E�P,`!�C�H�N�V�u���6����l�B���D�OhyTo�~��	K��/��xEP{����ӵ9��c)+]����7?��?�ݮM�j��\�冱��W�ԗHU�Ð�dѐ�L�C�3��hb���K�;m%�,��W�����o߂˥6V�1	?�+48���L����?�YM��?��6���@�%�+zRCL%=��'O�X*�ա��{����r��虃�"�������w~��G����o�v&������#    IDAT�9Ǉ����7���^��m�Z�J[6Z�:tڃ�L� 5�m�hH�گ%�/Ej	�6x]���7�&�����IC�i/Sop6�~��nm��k�ݰ*��4R^E����+�J0-�L$pJ����r@�����
��'p�,h=R0�B%�q4��'L�c�WC�(У" O Q�h��B4cAUAԟ i������OS�t��I#�+1>5g���p�t��������������'d�q�:�:&>)����"]�G�O����Ḽ�b�|L�'@����� ��&f�\pʣR�1�4�~�A�������y�@
�ؒGa(a�&�0�YLI���te�Hj�ɷ�~+iΑE
�|�T�T�^_M�̇�4���7��$��	4�K�HU�s�4A}p�X�ǟȢ9L@�) !�
r��"H:Y����금Z�B�,��FQ��x�T:@>��ɤcHa^�PC���ha 3@̿���Imr�SI���,�]�i�4�a��'� ���TE�	�D�3 cA𡕴�3��s�ɢ� 2'�y�@Yh��g =����Q+������3!u�z�i���o�9}���eת/��g�*����R3aڟ]]t�����&��f�AvM�ڠ3rã�Įf�b�`f+~k�ژl!�4gB����B=����2ͣ��K�?���v�L�̿���W�4�y���W/v��on_��ɶҫũ�]OJ��b��z�������&�Wm,ow7�������M��w�n�e ����)�Q -���e�*�6T��I�$�4�!�d�(-~��|@	҃����)�5R7�ڡ>5�����$*�]zV�,#?��UuR�Z��P�� �2�I���$�E�FR��4+Y�P�]�� KZ��L-�p �3q8�����)���!�<��,3B%�'�X��H�%]�F^C����-��u��mb���r�����ح/r)�չ`��]��i����oD�/@����u7}�ꤙ�6EЮzSĕي�c#�Ԓ&�Z.?�,�C(&H,�fK��s��Z"N�/� �J"1����r��*�\�&��!
A�@(!��C�,k�5��CU�����;3�F�:#�L%^�:ݫqmL[\>{�'���px�����U�J����B13�n��?�P��ܘ+��cR���k����YԤ�=��?�h�Q(�>UKi:Ɵ�f�� �(?�`\?H�"  �,�� d1?�᤟	��)�
O�:�*��g*2!�L�TEb�����:�:�n$�&�����bҩ���Ϛnn�����i�|BCuU珡�C��񳥞��0���>_7�S�5�F�:N�Bo����1�_�[ ��N��K�L���>o��D�(	i6ƫ��cW���r��S3�I�����	I�􈛀D�I�����*�y	JC+u����\�_8��r��&p�Cm�.����dϪ9(>��g��k�?_2�]5Օ)��~M7\Y��Kx����_��_pS�zs~���~>��q�9����J�B�U����Ωc�Vʴ N��A�K��ͨz��Q,-�o@��ȃ���a��{�0�! �(�3V��)��\�/��8��r�q5��a��P�08㋉�iUZ��C���L/���L?�zp�07?��1���pί|
�N�����u�Y{v �f�-���:C���'��:�����9�M��"�ZQ2.�uDd�fz�pH���_��	Ɩ8ƃP� �#�z���&PF 7��Pr!��Ljxl�M:k�ͷ�̖�ܙY˺7Vn�N?8N�g�m��0W^,pH��Q]�׶T���}���o�\�\Y���?��gާ^
��Z7uHN�iEZ��̏+��n|�]S����U��ut�'L�aʒ����� �c</��B.5`Fz0�g.�8�6�8q�����U�\��B�A�#�~��f�ꕭQe2�Q�r���f.R��A=u�[�߼96�pBbd?�kT��&0C�T��M���:�s��:HQ�|Q�>S��N 
kz��Ѧ�D_/)�ZQ�-Y:�XM��S���Q:�5�2��v�!?Y,G,a<#a
 �	�L���;�a�JLI���5��
���"F%����P�q������œ_.>x�ȗ�w߼y�f��Vu��&ԑ���0��#;)n�����rs��f���چ��G�U=vI�#��F3��p��:sS�~^����������H�66t���mͦ�mn���K^$���+K�fW�]�L����E�!W���i޸ͼ��?�s�sV�E\� ���H� z�#�=L<�����b��R�֑WN$ʒ�[�i���w����q����/�.--��t�;�ʹ߽vV�|��ژ΢���[P\�RRFCa����:��]vjpvZ�o���ّY����.?�:�f��������b;�[C�aF�k�zX굇�V���Q	V�<m��&�؎5�X��yC�5b"�|�m�:[�)	����,�+i��{��Ǥ|Ln����x$}����%S��Z�>��5S>H�(軽�����z�u,�үik��`���1����wR�kɢNJ�:a鴱='�E�;ޚ/����n���g�v*�?m�2�HqW�`��Qgi�2]�?��A�{��7�<��5?���;><��;O�~�MY*����%N�Tl�3ϟ?7���3MO��s00��+p)x\-�{x-�Q�f��t � B]�8�ܢ��+��R�^,�0�x���h�����O���׆��Ah-���I�	\�O����!��5w&ܗ8e}me�L;�gt�w��T���˧4չ���F�/k�ʴ�������G<}��v���9{vn�O�{��o�lWŸY��k�t����)��׾��o����S��ܯ;���x	��õV�Ƽj�ʴ??0�3Ur1�rr�M� ���b� 0ː6rK� �6 ��B����4�d)�p�*1 d�\1�`F8
Έ��v��~@�c�U=�X�7����s��������Ԡr�q�U�8�YG�<��!Y���i�9�����%T0]�GL�
�B�Yu�ũh@R	��D�Y?~��S��52T�f}%t��	O?��"T��,���S�d�G�O � |E%FAV����h3�Nz�QaB & � B�s�؏=��m���-/�^%�����{�N��,�Y��t�P=�U�N�ءn�o}f{i�ϵ*XH���T����S�UH�j��+qJ�J�UN@p��@� �R��븅�d���c�彌sR^�l�W��R(Xu��_����/�J��v����5�9D��MBZ"V%�4�e-���ǲ�lڲ�����bEM����b�fF���w��˯/��W]��.ۆlӐ/����������~�WZ�:#%�f���0�ϕ@�TY�@�O��AJ����6�Qc8״;���O��� ��+�^J�^���Re��+)H��{��B�ZK��]�� As�,h�\���>9_��I��?��?R�]�+&�hB�dp�� ���n�$���Ã����-?���pb���ǟ����k�����6=xhEߎ�+�N��0<�y?�[�r��I�:C
]ի
~Im�����Oq6�_��C��.��wS���z���6��{��绋>�`��&tqMg��Rʈ	x��:�/^�ݵR��Ì��� �'A�"�+H(M���
��8Y�	��Z&`�'�>�&���`F�'��HC	e�U���B+�(C1A�Ӂ�3�<��C���BW�b�9*�a���g�G%�]r����Fm�Q���e��Y���8	�&J>n��G����n���3�ß���6PC��.��>�y=�����R֧�'K�e��-�0�2?� N�	Wh/� �X�O�?��?3�	rAn��9�0!c)�+M+�
��6�4G�VU%@���`BmMD ��xJ`W�$Z#��8L� � ��!�6K��#K.����\<� ��`��$�?x ��xDE� �u���P'��!�L%��<�9�@(d����B�k@�:67�%\	"d��T�Vȕ�H�v����$��oP�q�'d��B��b��8J�GBD�t�"]��B�G�x[q�i�n���0�}�K>LY�y*���e�
��l��v��a�G�����ߪ���toל]��d�ʬ����vs�K�IY9�=���wW�����K�Mδyp���c�__�0��P5��%:�Sy�g���-��n3�u�����k��+�~q�������_�sO���¢��&��s넨�r�̏�W�n������f�ug�����b��%;ε�8�8��qA̧�Yʷ�DZ�>?��5�m�	�9��VW�Gf��� AB"�?��Ia�z���r�R��r�[)W�j0�
#Q�h8�
�h>�́�QU2�DC8�Ӭ0ħ�U��vANV��ur#��%��-Y�G��!�rX�@� �?4�p�1���I��0�(6��'�d�kEM�<��V�W�TB?ۺFۜ�V9� ���(�x�'RڭV$��v�j�^��B���ś]�;ʲg�d!Q�0�M��� ਒%�L�ѐ����q��1	T�d��xB���gp�4!NZ �4npp�ϣ�ܠE+h��@OB���e~G/�]Y��ixtx�3�~�iW�<F�������/}9�䪍�V��4q�?�6�Kk"�nu�}��oGYMU��T����y�{�LCA�����A���$��HA@ ����G8��Ȩ�PA�V�@z8�{�Ĭ`� 	�f�&
�8�̪٢��/}�	W��,��"�x�.�dF}��첮ﾼ��8|��[)����.�X�.�l'YE�4�ؚ�\SQ5P�<K��������<�+�jӦ��n��0�z �,2(���
���Z!V����P:�@Rd�����8T�s�IN�H���R�E�}����h�X�,�H`R�����{�����<��|����[<P�Z.�$�ͣ��c����i<@8i��%ʥ��� �i���@���<e���֣Vɒ��I[�q��墍D&�0��B�)-�������+���IJ��f:r�X���S����@Vsaf0K�W&��GmC���ڋM���h���
�o9�٪ZWo�Ac�=���mj��fզok�4Y�U~��!΀���I��7�q�&P?�A�#L�aB@a��� hP����
����8���$��bjj\��li�[�Y��j��2Y������mߴ��Է���Ã[#���Y�~u8�;����>o�%�؆PS�4I�`~쒖�h��<�1Ρ��e�c��[��KC�q��p���fl�>�H�b�O����ph�1�|���a��Y��\�V���zfg+�o� <uIO��;�^��%|ho�ɥ���y���q�I�T�&�O���q�!��M���KK�ev��,��x|�,���Z��zc�c�ȣ\�� �OrI��1*����0� �C�:--�����\���:�=Z�G�C�ǣ�DӠVL�m��I����ç�W�����G>J�X�jg�X��T���1���Օ���zo�=�(Yw��}%�bgU'�6M�ވ�՞N��ͫ�>XP�{�6�����V�m6H5"Vh��<��o?��D�Hb�'���H�� �ް���TQڅ7P�\�6�Y-&|η ԣ0�' ��]��,H���`��͂Dq4��Z��l���w�����6�ӓó���j�8�t�`�b��U�g��pms�[#}���r�{rj��k�����%{-�yw�鶉��Z4���ꝍϝ����⢛i�>��}��GHT�1ӣY��:�2K���S���R1
&���.	E&��x������9�ۡ�O.M���i��s�D��\�Zq@%���&��g�'O��v��)I�\�-A11�$�yu�w�l�Y���d�ŏ�%.��%��-o{�;o�+6߯��5�ce���[���o���b�	z����ni?9ϭ׷��C�,����vFk�q����jc��M���wG�}������>��Z���U�][���Q����&�L���+Y��iq���+K�$�C(���8otJ����Z�� ]�z@o�8�ӭ����_㛷�?��n�s����k}�t�{�-�V�;;����!g���.���^o����w�r2Xt!
[ȩ��p�R��O�׬}��7K�Ӥ�*-j>K&s��$Kq��m �`�B�ȷ����o�����?z��\^���.�tˍmŚQZ�"}��ś7ox�����I���Ü&G+ހ��D`˷bh��St�V
�D�1d��FO�qVA@-��!���pF�0��J��C��bn��v��1��5׊9�Աp3><8��Λ�K|}���Ε����㶔h������!�jt�EU<��� s�0�1�'8T�G��� �� V�X���o��|��Z1í5���(�,�Z�|����O%Vg@54�\�!�z��
 �E��~���%��'
c�&�:���dn�(F��`��ai;=����ذs��gG';��~�m/ �,���,�
�S�0۵U6��u��L��S�[
�!���A��QD:qJ�n��d�M����,V3GHh�^����V���ۑ0&*��YG�����?@�Bע����[@��b!e�	
�#���O��`Y4p����f�&Zs%�k;l԰���K}��Xy���u�:m�ܮ��S����aԫ��4���m�PvЮ-.���owa���|��g?���X�d���a9��F��F=�z��eu�P sӐK����ԧ��>Tx ���o�H��4���f�%Tb@��\L�:�r�j�_��_����'�!����+0�C+ʸ�������0�i0�I�����t�� ()dQFLqh�&mL���1#�+�o!|s�.�7W�nn_^���?�}���'��.c��WC�j%{���8�y�`ߡ۳B�B4@U#�D�X�*�������짺Ґ�<������f��d6<և�BV,U��4Z�s�l��
��%��NA�� S!�CF�ihI� +��uI�YB.&A���&KUX�>���K�$K-nH<�T=��`��8LL(#W�ƬXՐt�j���R�[��}�X��X��XM�VP�����'*�v$���r	�@U��ǯ��Z�DO�v�ZG�GH�Q9i�X�I�5��93@bE��ɥ�3�D ��A�W�7�"�o�$�AQ��lo|�[z���SO[�D�$1wiqL0:Ѳ�g��I<	o+cG���VO	�BL~�:	����ܽID[j�şʠ�3*�J�����U��@�4�(�9>^<p�
U�@���m�y$ݯ>'�c(�ਢr�/��a��%���䪽��o�Q��'>�Q�J(�8p��G�B�W�<JLP"b@B��\$�v�Ap�s:C$�d���Ed1T�L� �0i�7���0lw����ͅ�������>B|u����ֹ��J]zڽZ�]�ٲSO."���f�{V8'`Ra���vW�N���Ň��$�bT
<j3JB&d� �\WY���o�r��㓗�O.��Q����ۜPGWZ�Y�|ֹ����O��dKë�v���ˇ��u�#w��-k�*6tkW�IH�'%RFL��	�(�ρ�  �Dba�d�!�'&�U���*��rp�,B% ���T6�)�6�`.&r��u�Z��
NV�����\�O.����8*@\�9d�Q�r�pHdA�J!�(�y��� M���H�&BT������"-<#Օ>T�!�~�S���S���\�O���k�a�ַ�U�ո��yߔPj�"�x|�d���*j@�#M[	&�!�L�Dҡ!��K�C��!7����iJ�p 	h�4���$&n����8@1�'Q*5�2�    IDAT�q�г��+�ź��M��f���lI�i�,�����Q�)��2��iE:n|B"5���.�)!.���N���\O���� ��sGi,�!�e�U�m	��'�C<#� K<GN>VR����,�$>I�@���VB�+�OXab,�P�~�����x���L?�H�jԱ9��9q�fh��+�,-�0I\n"Is�s�P%0p̱U�8@��F7pTI!As}�����#4	1�G�H�F�\�pC�xRa��a��hǈ|1�0���{D%�,��h"�D�@"=�H$�8Gn�T�'��rᄹ4�8B�!O���b�^��ࣥ3��8�H��u��*�(>r=�h$<b�.L���9f�� ���<���+h�"r �@�$�2�cea�*� �[��ʯ$�D83���)�%"B�� 'T�IG�P�iBI�819�g�@�DC	�hw�sa.x�h8x�r��Gb��\O�=�T"*(�@jM�m�W'.|:�zj��v0;�vq�C/WK��h��[ll+G����I��Za�)D���J��!�,�����<4i�GT
%& �a,N�cLF�� �K��q����1UQ:��Ib�0�(#�+��'8��c��&H�U�O�9Hl�K�*LM��U>���0c]���� DC+�XW�J���\�F�u����a�iKU% �k�48>�&]@�#ዡ��h�QB�PB��	|H�sм�5U-�U
LA��R��9z�.nL�)���hfo����d
P�ve���9AeEa�����ñ7�c�h���39�ڟ��&����m������FWV��LY�\Zk~��R��Zap�{���9�8�Y����zk��cf<«<���{*�kR;S
A�hqi�%�3�$��?���y n̏;|R"����$|�K�G�� �: ߣ��t~6��-#md��R�tؾ{�j�OL.��V����w��� a(V|���]�頬/�����b�<�������̽�Q�ʄP�a���V��U�u���ߍ����y��i�N#N�R��tN����ɓ'~�i;w8L��Ŝ���f���۷f!8���0V{�
r�)�#�I��KĽ�E?� 7l@(MC��F\�	�bdܒ`|�9�j�YA�xH�*Ӷr��	�.ۇf�Ys��Ĳ��nNB�-�4����(U����.,Y?�x��:�j*M��3w}��ظ�cd�P�1��x���X��|���Ͽ���w�֖
j+�(�l��l��ٳZE�9�P��)�Tf�9-*��J��6�?�6����3S��d&�?M7���F��?u{z�e�&8&Ө��AK��	MZ��q�����6s+l�'������hM�˖*Z+��/Gt��p{J���+���+�"�c^�g{��j��&I|���l��d6{���?��?����S�Iǐ�b!�c�����W��'Ŷ�>�89�Cf�\�	�8�'ip�'B%P�K�T���
0	� |	�JG���b�@�8��h�ljgcPcl�_>��3ױ¶��8O�p�᪹�h��]@�5�G"V|H�<�t���A:��-azLݐV��%R�O�ڣ�����H�9�J"6�i���ׯ}k7m�2�_F������_d�GdS�8C�
���\�G�R�th��$��@�����ӧ��kZ�?�_5�ݩ��r��u�FX����#�8d�,��g�ط�������*�l����ݣ/m�������g}D��g��|��H!R2%.A11�I�W�f�XZnH$x@���p�m�PZ�	�4|14��4A�\��pō9n��C01�l�Y? GQ*��D�g�"�B�	���W�$b�ǘ!-!H�Y�1���פ\�cW����#F<T��R᷒��Gu�~��.�+,��p'Ɲ��;`��aq��`g�:޽���Eo�*���;8����_P�_�F�h��w?�����C��OT,��� �Һ��Uz�����E=�*8Y+R;�H�S��C�P)%�٨��t�MnZ&��ƀ�J�Gk������?~ldc%-M�(f<aR[֩%��\+�pݸBLp�����������`������黝ݣs�/�p�����������kY�.vW�O\�eӡ���4\�ѽ�qg�S]m'r>��RjQ}MM���,��E6؜;�>\��ϖ���o����O��+�r�r�b �B��Gh�M)���	��%0<	�0eaYZ�<=
��bY	����!�<����	din�,�j��GI�/�ʣ!��2a
��*	�
�k���J(n���6���+U$�r#4VH#�1�\�����XY�pI�Da)LU���^5_?Ns���:=��/�h>�9�&�󿹺�'?����s�3�x��pH�e:$��vx�8b���dG�����lol��	�I� 0�}����[�
YYO>��U}���������"�w�g*C��04.[�{���FȺD��쇭��Q0�b�?lVz'Y0
Bx��5�9��C#N`�h�#Z3�� �'���jMl��&�٬!l"h�ܡuTSD�	`�l��	@,�潐�IV��C��A�1�^��9+�����e�U 8x#w��g��60ƨ?<[�4��Fa-�.D�ĉxMcT���I�
�&0 ��lh�[Y�(��?�2H$���"�	V0�|Q�3Ø�t�nY�\d���M��gg{|�ȁ���r�������Ǐξ�j�����Ž�/�Z�ގ��:��/����p|Bڜ��Xk��?�}���㭕�g��t�J¯ߟ�r�'��#hK�-A�	
�
�`���oL#�מ�_�rE������_����/.O�}E�!ܦ�ʂ�)8�~:G�^�xzu���ª}������։?Yw����.aXv;��}\@A��vђ�S&g������
٠�2��aZѪӣ�MҨ�ƌA�SG�G<4�9G�0TEK�����w�B��4��m{�פ�dh,!�H�x�)�0_��<Xu����
Lo5M)��Z���g<`nf�X�la���K?S����bB���S���;�Pw�ݑ}��79�pn?���T���˚�Oًqڠ�
[S�#��f*zi�9"�RO �Ąhh#�i�E 3_�0D�Rѕ��l���`�� )��j���(r�+=/�9���c����m ���a�a��Dn�����[ⴇS�z��wǕJù<=ߘ� �?��:�	E£���9j�0 �*4`b �/�z��I/��x�Ы�p���v8����1o2�C3����O�0)F�]�Q7�H��m�f`^ o���&r5+<�h*<�yT7M���q���K_��[0���TX�e�P�P����
=���*X,�����+sVd5%����Ս�`��4J]�Cz��;�٩1gN@?��Ā	]0��a��ʉ�2���`��I֛�NH�E�	* ��s�;���B�d� �����l�=���و
��`hdLM.u��RW�$=9ׅ�����u!a�6/��K)Gz���G��@�4�3D����r�W�S%H]��à+M��Ϋ�z�a�S����f&�n!�s�y�Q��Kc'4G�Jr�?<*0�iȘ�3O33kV�)��RX3�P����ՖF��_� 4)qj�`\>����M�~�]�ɽ�ڷ�=]���2ЧӇ���9�1�\���B�N`j�"��,c�2���s��0B�����H�7j.(��g�#z<
�B����Z¬=0&�ɜ���/�^M&��3�����.��J��ң�\0��4#�)1�����\��f%T�c(�ޫ��_�j��'�3'6�3�	 %G� ����Xt)d]jl�-+��i8"4�@E�W�7�B�Vh���FH�$?~Lc�Q��d�:�CU&�/y��0X�����E_��wA������/����o~����Q�[>>��-`�R���7�<Q8�=&kmay�{��:4v��F�/��5����}O3��.����<dU��A��ڗ!���������$C(���f^�?̽\����,q��,��^H#�i�!�!K  f]��H&B����tǯ~�J�Q[0�9BMʦ���3K�G'��|t����r����e�T�sն��˧>�b�.�����
�s��GD�4��f�{�����ЇE�tƝ��t\�g_�D2aD"6C���'������]7T�o£�k��G�\�~��|�^t�k#�,�l�V�LY�axN�u)� -����l����bD��Tb_/BCc�B��?��3]0���d�h�~�ȱ��5R�\����oA���n��ˋ�rN+�V$��xi������[;k~q�A4&�l���5�&��p��n����?B���z����}��z���x��^�_���Si�Dh�\O��k��^��e.`N%jD>-]�D�-9������.zXb�^/�+N��d����KRRY������^M��&,�<�F!�o�=.�X���7G����ٱs�Ƞ��=�3�f�G�֬��7Y{�k�����#y+��O,{�ߝ�x�͸a��Q}t�C9��Z\���8%�b�d��p��YN�ȀZج��A�2*��s���*mjh�dN�@_���x����|aV�#̄/Jrd�3�ËA�,����2ua��t����ڑ�}�۩��}+f(���5��cT]���PL�9���}Y0vq�d�L)o6s��X9�3t2P�^.��.��J��i�&fO����W�K:�#����&W���mאּ�Q#�Q��Xe(���b �LJYQ:$��'��AG<0a�\�qs��[k�n\�u꯿|rt|��o����;�no�j������檏��
����ĄE?֘�0�F��4q�c3H�HW�$�Y���,HH����T/��XUsA�����M`r���m?f��h+hRzj�G9�I���-��D���@XH����hma1�!SV���C�����l��J������X�%�u����c�Y��_��8���[������M�����o<������p�J�σ{#y�@
@<�@`�.�۴'����xC 0|#�k�D��A��ؤ���z[j���r*{+Bs ����n7�;w\�!�|I�ej��5����c�-<$G
/xx�%Q9;�E �W%*������ڎ�n��b�FÑS7T����(N�<���*N�<���oO��aN�N�?|���_9���W���i��Vn\��'R_~���C�}�k��g�c����k㣴K�(�����e�¦2��+�,������7(��l� �8�8���ߘ���X���f�TV�)�&e�m��m��K���Ԇ��:%��s*���~$a:M�UI_$4l�J�&*�ɹ3��LTYq`�Q�ThrM�	IV���Gu��/Hx�`j:�$[r֒��}>l��S�|�fA�i�@�`#�I��`�h��Fq�k2�%7\�����5�qP���j18��adɮ���A	 F0�2�2�"4<�)��(8����m2�ЁM���̤Pm6�Be�B����b��l_�4c������\���pឥ= ��x���;��	Ois&;��!(�!�!�<{;1P�i�s�X(��"�p�*�d\�|� ��v�dBP;9? Bs$Mfˣ��� 0��?�/��*Q!�	=M�������l�-�Ȍi2e9�\�r��,�j�-��N�wL<Ra\d�tA*s�2�9=y���Ȕ!)��(e8�^.����������x������߾qrp���w�|dƧ*�^|��d|d�����_�,�Wo�Og���n��g������{���|�`v8�9N�Ԃ1�qx��γ���fq�iA�<�i ��^jk���K^����u�ϗ�"��85�ꄵU������>lH��8�����F��Ɖ��?�����:1[��8=y�/��}m��_�����N��H����ր���`��@���j����i
A#���d0��w<r��|e�i��睬D��ڈ�2��1ﯯ��+�7%����Shc�NCo�sZTy�ѫ.�D�VrG�I�){j�
062%<�ѩʬ�_�_��c��E� �yW�Y)Q�6}��v��A��.�c�M��K�M�-$�z|S�T�@�
�F�Bl0��<F��F�������R�+���dTHh�`V2��&�^zJ5%M]j���k]�Prڦ]���_So����'F,3$e���UB_����5���:���S�������:.�M�hM\�����CI����f��i�Cc�;��+eX�S���	�-Y�y�
�^$z�3�M�d7��H�ئ�j�HKM��R�$ h��#�� פ��K3�:s`�����Ih�L�Q��rĦ�k��Q�.�� 	��y�a������E��&<MC(Kd/3�a(1ӓըҘn1|]���kr~��Ϊ�C2�A��Hb���	f�l�-�0�2r�L��(��1�5� ��Y���X�d�@�<$%!��d �1�����0�scdO��f��Ɋ��:�`��%4X ^r��T����ԉ�y���H ZN�0`蝩N!Ŧ�
���sv��M�#H]���iJ//��� �`Hx�}	@3�^02=Sc,4J�#Q�ǣV���\���F/YoB��l����_d�2��_�.��D �w)�џ��qv~�/_�
�����X�;"�g�#��oX�	����6NT�����d@*`h� �'�W�
V�	�
�<�ؘ2]�E�&X2*�a2�- GN0����ƤZ3@5f�(Kd#R�<���\$d��U*���K�JZH5�x�D��6Nw)� ���.bE5+�xy�� AS�o�cP�O����Q�ρ��d4&��5�� �U�x4�L���F���hb �>zi�D���%�p�����Jz���CR-�M6��0ߟF!ok�����W�{?��ۻ7�{���?�.>���(�<��99<;��b�+]|��y�;7^!1>���鹗n�H�Y�˓�q�I���^�nA2G ӯ��"TJъ� Z�J~���s`�՜[�$�M���hu���4���(�j^��#{�Z���J�f��.����8Nɧ񻞭�$?�qf�FSm�1�9T�"����;�U��?�޻�������A�Q�Msi����C��޽>���I5w���
��8Y��ۃn23^ĵ�a,�=)KC�QT�Aف�Q�b�<��h�`hԍ1$%C����������Ə��[	��[ld�s�pҏ�'�o6���r�<o2�R$�L��b�X!�
sYe�_[��z�7A0]q�C�����=4��x�:�q�dk�u�q��]S�>&�=p�ȈHb6��뜙�_y%��jo1t�u�b�W[�ە{7��eu��t�hk{�����ow��v������9��ު��XkL��6eɠJ�3!(���F*�բ�$Fm,06�0L�H�G�`��[-���}�.�4�7m�i�9/�D��(��k˲��h^z`B�57���t)c��^�j�a��A�^w�ϻmH�n�ɿ��;��kvL f|����ӏ>�6sƵ8����5X9O)�!�jby[!c=L+�P�-����"$�yB��$�T
)��5��.��
��V/�R/�F��;��1�z�l9�T+u�G�X�+�� �V�E�x��������/�S}��i@7���>�e,����*cR̀�<[�dA�K�nQ9;������v�28�(���ҭ��w�� w�^ؙp��+fl֕�Q�d�� ��2����E�����Q��An�ˑ�v���_Y2���),0^�p���� �x?z��&�"±�W׽���k����?����x�xa�����3��<�����q�u�<�l	{1�����M�iŽZ�h%V=;�dr�#K �8�`�+K�m�z)�)M�j z2r��<[<Y�-�I����R�
҆f��G�`1� �K'J�vQ(ȵ.��c�L�ɺ4�7!��w��t��ݤ    IDAT���$���с?Nq��j|�x���sWq���"(sK�=J۾�̞�NQx�ߧv�]\���]n{>}v��rk����a�����R�`̘�9���aʂ������ �FڦSL�KY��gAK�![�2c��N/?���۷
y�����M/-zu�K�üHl�h)Ŧ�D`D»;=�7�<�P�C~�&_H��&�/~� s����cb��E.���?��?q�euy\{k���������=o_|��兵?�:�ͭ���ō��v�]�v�j������s�:����p�>�ۛ�.�ٔ����vaZ��;�>V����S|��?�X�~��ߌ���ah�R!`���ˌl��0&�
@�Y��y� ���
Y��r.MG��1'�i2T�-ȳ�B-r�:q���2,�`&�mz��Q��\RQ1��'3ǌJd�`�y.̸�E�^)3��jz$j�`�д��O0V&* �9�G ]�J�d�֪�A��ŉG��d{���!��-T��/��� 3@̿��e_Fɖ�v�9�@1�j�
��������Db�t�N�!�#Z���le���Hm�|��De{W�ȶ{ƶn)c�gB��`㨩g.]0�����#�^/ Q�/LD^xȑ�B�D���9fw��J�_����JqZ	��e��xĐ	s��� .��� E�.W2�ӟ����1_����/�qg�Bb8�I��r�!����`t�����|��)�MH�-+J!B�a�$7J�*��Yxj�ls��Kl�r˼�D�����W�.��r�'e<L(Ց��\/�����G��{�ƭ������7��?���鳳��K?SV���V��?��yk���#�85��f��wo^�����Nܲ?�י֛/c��W�����\�������0��^	�¢��?�Y�-�efe�����o���l�Rn}��)��g�rW/�Q�&���<�{7���[^�^4�~���k�X���/��Oka�<6�aQ� �P�.�*�YW٦�D-�rn�5^�𱑹 c ��:�]Hl���fN�E�cKH���#�.�����.N�L�V`p4�8Q�)�C+Jo$�A36��;!�����xP�EHIF�G���,i9eC�J��Q)�X�c���)ɍ1�����+$u��f��x�8������N��>�f�s�/�4yQώ�)4E�V҄W#�a��yT�UR�U{]2�\C2�G�0�;<�f�Lt�c�s��H�J�T[{S#^/���@"��lU@��q*�R�?%C2�)��624p��̌��r����\Q��H�D<�s��ѩS�����AΖ�֌G3ۺ�HÅ�a]NS�����d&�T�q��.~s� �G�[�h�kf�d��a$�x���%J0y�� )B lx�l@S�$ͬJ2�\L��¤'��P�/`��fK��&�B�D�\0�li�)�h��i#�cV4\�1��s���T t���$$��QY�A/��
fǩ�k~:|����:�4s��l� �l;Uǆ�B��NSf�sM��#[Ma����E�W���^` ���b�0����'X�tQ�d[$�# a�p&��I�%-/Ŗy��-��P��A�S$�4"�dUM�W1L<��)�lX�ԩ��%Ϛ�-`���&X��B�f� A��.�m���C��� �/M�5�2	C�a�D8�w
�����5�Uk�i� ��l����8	�����x	�;mr`'n�k3e|��������N=�S��b0}�k:�`nt��&d+_�<��EՆO#H
g�A�j� �z�dE��+z9�:2_3��&�Lr�f<Ysӥ�"溆�ׇ�l�̈�b`�zz�ȸXa��Hr��3t4�%<�.$lÇ;�o�WJ/AϤ#��:�E/e�+�¨9�1m�o�Wf��؊9p5s ���M�*sW3Ȗ2B��4	~�*$j?Ta�Ɇf�e�Y��%���hV������߻��{Ϟ�s����g�Gv�7�������Gn6��
�W�O���oZ����ͱ���CX�� ���^���!�\��_����rq��Fl����c�pI�Kä��F.��M(��n�<x�Gk�j` �o�֬1$�*��dH���%4w՚���&�Aav��BY��3]IkE©�����]�]n��7��3U&v�����8qZ��A�),���o����vB&��et�����
�]�]9����v$�lb�+smA�]%�
��$!�	��ZS���r���JE��T�	yD5�L(����J36]�!+��l�k�1("�:ٕ
 ��,x̮���8ȼD.���𥈕�Iv���w��Q�8���dK��wg��ǻ�ې�-7��=�<�`Az�Y�2�fS����N�7�L`�O�/.
�%���~��;߸����uXZ�^x�EyS�<b����)B������~��Ȉ)Y%�_�@�hȆ c	z�2Q��:0�G�,h��.	r���K�&����֬�#�����*�b��#�\��d�"�T/�.\������x�B�s�GT�S�q��[�q�ń)�+�Ӯ;;{�����]a�3q�K0z�9G%�S�%'�.��8�%\���SxG��0��i����.TVf50@�]*�� ��E�R)����d:l5� �	৴�`�LL�JVׅ�<e۳���z��X����Q��F���w�Ϗ��u�b1{�׸5��U֜K�%'l&�pL(Y�K�h��KJ�E"x� L�m���"d���6�*%[��u�!����!]��!�e��b�J	�#���s��hS��ڰB08O�L�YC	����lř!60N���wmV/���.�S~콥���>wW��|ܘ��l����P���l�Ɵ]������y,-��8�U�1E��+��B3+����(�� �� hk�V[�`�0��T�%H�����s�M�cB�6d{�f0~2}�޽+�_|�N	���8Xj�&[p�6��!bM ����!��P�I0�]/��[�W0y���g����D͎!��xL��u�lzy*�
��	aɷ4ϝ�8<߻����⊷HNN\f=<p�ō��jmucsk��Q�1X�����`ҧ�^��Gu�J+I~�"��r������ˆD!����W��BM��<�QX��S�W�!���	� &�������`���C�-�c.5��o���c���y �/`xە����Kx
Cas����ε�{;;?�{��-Ϧ={~��ѷ{7������-�|�ts��%G������S�e���s_`r+�_�yl�A��Ɏ�|Za�
�+���#����8�܊y�Km/W7��l^���\9]�a��䴾�^[�h�W���f�M�&�<.�Үi�j�k��Ja˰�ð��[�A(�	
�& Y�N�լG�[q�k*\<0L8қ~i:�(x�	0j ��g�Ǭ���b)�jS��/!� ,���)"d��GJ��zɺ`��FTzi�H�X�1�饋F͖`A
�:o�@ECF(���~"a�H�ƋJ���J6�Ap璹.�-G��ۋ� �;M�;l؂xTlmY�~P=0�mk6��~��&�mJ<8��#�m��{��uq�i0ghD6yz��arĊl���Y< s�1��|1g�PYB�0P
I2%֐���ֿ��^�4"�D�W�rD�y�R��#�4���~��F@	�;Za|��gl�9Y�8���D��c,�t˓F��8+��| ��^;I�"s��^5*��AjJ�^$L������WdR/�h��f[�լ�!��(d$��;��/ V!9��O������G��։�'-����K� �w�����~�ci��˗�{�_ZX:]8uV�w���WK'^I{vr�������>��'��������מ������3�૮Y*0�qj�֏HD+H�P��Ŭ�P�ob��==ފ0���Z������������ʂ#���Ζ)�i���£x�H�1?^���Ļ�}V����˧/N/�]�^[:��t}�'CL�ْ�WX陋M0ʛ�̗�3� �4
�X�	4b���f.f%@CNP�
0�La��!B�I�L�^E����
���z�`��4A�d0%!�z�`H�#1.���&�&���� H�*�"�)!�x�,lJ�so#қ_d.�*��HM����"Wj���i)ۦ(��`l� �~��1��s,	cU�`�6�4HJ 2e&�+!�4#�L ��J�[<�b��Z�S<�$C���`��h�z)#��,������`jJ�9�@����t���`�<%�1
�<���a��C���a&��ώK	>� i�Ms�ܦ�E�6/-�a�z��u���� ��ʵ���3Ak
Ԕe��g���D���!(x�BBE S@�h��/lޕ��$(��� =�8i�Dج���(��F�SlF�z$��R3s&��El�it���$c+��i�P�[M�C��dx� jV��!����`�Y��X�A�D��� S:H�U0`L4a&�W�� t5�`�S�0�2�4��\k*��§�Y�i�4ב�^sD��>|T�%�V3��8ç'�P��F���LIM�e`�]M@l���`�h��jz0<QQ�fi�7���FބJ�]I+�`�!)#D%�ST��Ő@�y.
��9d�2A�?��`
��0�=���E��0b+ZJf5R�^���L�� GB����6=�0�D8�MW�3�/<g�P�0���#�ӳ���뫫�����pʳ��F��yv4Q)�z�[�s�W�"Zxz�i�R#d^���>Ms2������ M�y3R�5	jl����\�v^u�0�Nor��2I�Qgܨ���N���8ٚ�A��fꗔ�o�H�aZ�9�#��b�<�H	����(�u��UL0��T�Sa�(�j5� 1[�eX�s���m	���3$6���~x",`VX���g?s1�E��D��ػX�R��v��{qr����7�����'�>��g�n���vuvr�즉�2b������nN8��t.�i�Bp��$�)�_�~���6RpyI#��&�EX*t��^2�Bc���f�o�|�l�ö�K ��Z!�%�$�t��+�4�C(u%�y�m��:��Ȳmi�!߸؂���/�HuE�k��hnm�g9n������[�����n��\ �㦚-z}�i���9���_N �U�+�;J��.������X���!5pa0� ���� ]p��g�xdK9��Q3'4AƮ����8�9Gy�:%��i��R"��J�i0�.��� V�j��Pk����y���L�'��`.���b�{���G�&ڕ�+gA��gSqݫ�u�iI�3r.^��3I�n���]_T}��]z��w��.^��Wƣ����w���#^i NM#Eتv#G��4`4���"By(�N��]	D]�	�#�0F]��5Ũd8�.��� �0�c�頑jۻ���]� �0=���y<zy�G �?O%��lr�>�w]{�s�g�G�,����Ĭl�/�^�L����4�g�_-/ݜn!߽{W��7S����͌�d^��/�������.�ٍȶ���Ic�OIh��EB_�4�M��m8�*"�?��r7�d�����M��&~��hZ�z#�$�5�l�jz ���L;o!(����g���7�K��ozQ����_~���%!	���h���E#���g�q�������q�X<�_|a��j[��)B�Bl,�"1p���h��D�JT��wn��ڢ�]f�X��־��-?�kA��G?�'+��/���.���g�.��ȩ0�
�C��TG�~����?rM�����s��)�ZM�wB�?}���[�g൳v���wa%/�h��{���j����bh��5��`�ƫ��Yi�W���2.��d8���Pʉ���#5C�z)�e���^*�߿��^�)v�M���Ws�	��´�pP���8�;�]����
A�L�����Y��ٍՍ�����3�/}w��s2���]�s�Gf��١/�S����+�[NW>�iO�s���6�����l8��:�<��������/W�/jw~�����Mk]䆩6R�\(�ei�l��2(��ucDƞ���	H����PJ64J'L�
+�6{(9������`�a��?�����lu�@�?���/Mz�ٝ�'N�/���_�5+;k�p-��4)�V����m<��� �\�Ǧ4|�����/#��] ��͑���o�~����6�|�������{�����Z_�����l�\{���C����q�h������ُ��>�:���z�˖��
~Y��E8�;� o�Yp�|C�ڞ屿s���i����������u5�֫3P4eCm�M���2Д�#!蒐z[ҥ��F(3���9J������.�B"K����B���S��&p�HT 2+!�ǔ�>��g�D�k��25C�EȻ��j��R�L ֕9+��4j��
��J j����{����
�J��)0`�=�0�x����������4V,��k[�0����=�^&NьK�	�Æ͖S<<�5���N�tVΤi4�*-	�0�f ��خ��)	L)��&+v>(��|G)�@"�"~B�fS/p$r��S&�4F�^ Nax�kD>�/V��I�`4�'���12d��Qa`,�yԤ+`��m��4�l����,6#��9�oTۡ5"���6*��N�<
I��R�,�@�)�&=~E��$�1k�D ����bH���Aa�(�le�U�yW�#02�4�e�(���e����am�̕����ŋݝ۷?Y��o�^�|y��O�/.�.��ٍ�C����&���[��b�_���߿{s���3{����tv�zv�Dv�Ƹx���x�M_�
�x�Yx�+�r�W�[���=Q��p��ј��#|'s�ʂ�_[Y^��'������~�3f�S�\��;�����d�ɋ��cG����~�r��rma����p�ۨV��٩.����k�����2���)И�0�`��d�01L��y��AK�� ��ڼ`����c�r�*�6����ro��'6<�d0J�d��P� �&}MT
�Х�Z3yB�/[<-`L���R�I3g�0$�$�Y�DWB� a�N�oRx����5[0e�K����]W��g������I��`>�\�QC�߬4�*��0���e`�. !q�V)x�9�/2]遛���53�$���P+�궋�4����F� و�낇T���B����U�ȹS��AkQ9�%�c9�1�ǐ��ټ����Q�S�*��'�[J �L`j`���1΃bBLĚuQ�����)�|JzJ�Ƒ�����zɨ�
r�̈́����)	��_�\R�E�/]�Ou��8Q����KL$l��7�H/��DN9An�54$<�TX1�QSf��PldVx$��@��PN�#K
=;�x�$9s��@H`a�%�ᐣ`.�RD֥4"M` `szP`lŦ��7�8�ڥ�a��d�Z��n��F�Vl -X &0l�e���/-�d��� ׫��`fa0�-� dJ�
0$��)��\0L�	��`��?e�BUGn, �
�|FKCpZ�,�FT����B�=N���&Z+�.$1#ϯ�>0e��<��Ba�\�K_��hb���Z`�z[��jrQ<3<$��RF�IU.�s3$��:��I�뒦 ζe0�/&����y	�[qx��S5}���D��$*��4	e�.2�`4#��S���X�T�5!��c���gl�rH�&WV�|!��L �%��S<�t)V����^�C�����D�$+d��c"<���ۮ�a���B�-�H�/]O�V	b�1��b��Ӷ�D��k�|)��(�E�-B#JƄ9�&=$MH`�b��W] EE����l(�R3~ҏȦ��H
�����:��L}���1��:��ݽ��g���ߦ9=;>�t���>�n�|ؙ�m�p���Kh��و������L!G�~��m���R�_�z['���d��X��B�>A�7�Eb��K�>�{Yߜ��    IDAT*ژ�����1�iaKr2 B�R�#ו�b�et�ʡQ� l���� Mӥ�͍Z$��9�`b�t��D�~�7��]�q�Cc[;��O�rM�oshr��x*�%�]�5H�$���]��@�A$2/*M��X<J�jh�˛��:�k;���ѓ�x ;,����5��Tt�+�!�?�xW ���.%�&eMB'~x�Q˿e1��!�%6�r��^�$�ϸ����C�^lF�Z����<�m4�k��ǳl㾃+�c*=[%\њ5��&k�-������gz���wwm������x!���rDg���w��i���eU˶�ͻ.E�-E2<d����ț���)�e��
!�5V�2r�cӜW�"�7VQ�f-$_x8�Ŗ;9�X	q��	r�����6���d&t�[�����.�ƾb:?Q_>>9�\����N�O˫[;�jۻo���+��o\ڞ��]N�
�ײ���-�̙��N�FĊL	Ɛ\J%3}	g�P*����A�Ո��F-?ܑ�+y��IS�!�h)�5�1�)�`�#��'��͖�6���WJ}���ԕG���'ϖ�}������4$wXfC�����Q�!4"H��Kvή���0���Fl-i)�.��K��x�8FhZ��-Z���>�Bٜ��ɵM�}~�G�!sd��R�	�/K���_÷'���Ǐ�ڭ�4R.,!�䐻ӄ��j�w�Z!q��5R`C���6O$x�����ߏGWY�����/N�7�/��]Z}�3+������3�k>.��q_W���Z��^���m[�,��_c^]��7"�W� �$Ԝ�^-`�	��	�Ф�'6|�4�^I3v[7�L�X��o%���_��<��x���%/V 9eKA�6�� QcWh4�D�\)�ew��e��ڮ=ƺ���Uukޕ�l\?u4�N��Sow9v0z�.l����K����8.s�yf71�<�����I������,;��3�B�W�F���!"t�c��	z��^I��k*�n�iڮ��T�l�<+U@���M�R���/�ǖ������-ez���/�²{�����MT	.��ɟ�	$N0�&����#1�Kq"���
L�yᚆk����j���ð�ˈL�����p7�R}|��0LC~����������e��j<Ytz���w����o�~��X�7��mݸ8��k|�<dݤ��!��0��83�b:y�m���q+ڒ��N�_�tݭ���yG��Vw����
�����2����Z2�Z$Dm�ƞFm�
�ұM �^eO��
/� P'G8b�V�Z��2�KÅ��GaK	0��8���ʖ��
!�]<�z��4ɂ���$
��<�����X�-56��s1��	%H�h 9wh��	����K�Q�1 ���1k)�Hd�
��ht)��S�h�1��8c�2l��gG,$l��z�1�Y��V�H5X
���f�e�w����Q�|7Yq�4 f�Ck��)���C�͹��b����S�a
��[c�˞�ސC2ԔM�70X~�����G攀�^HS`�ْ�
;w�0��c_�vt��]CT�2n��p�VZ�޿�΄����`NՎ����%�Sqʰ�L�S���>j��! �a��_� �@z�B�Bru��[�"�7:V��G2N���E�B�C�B"Sj䥚Nz<4�J]���y��Ɋ���I�M�������zue��љW�D��F_�8q޹���_�z���>z�ճg'~ō�m�Ѝ���坷v���?���~��]�g_|�oI�=?����)�Rad��La��KA�,W�W����?�N�����h��b}}��wּ�}k�g�7��5o������AG��7��G�/�՝{��K~���9.Gy�����W\�}����^����͕�×'�3�N�ݕ��%�ܖ@JKb3͂^��n����&�`\Y�N�ȃ�a��uh,B����USb� Ao��hB�<9� �Cj�g¨���.<H����ħ4�C<j��7�3�20G�M��a��F�$�00$(L��o�S�b���ɋ.`��ՔBf�)<�`ũW�iD��u�r
S`�z�.���Z�@�*�ٰ���3��0q���M=Y$ ��!��7�a���4��MM��'��W���#��/-s�^)f�=�	�8_z�g�qR>���i����ٻƠF��	��5�}����v֐��z�@I6G�d�^2�&�	Mljj ��0�iV��ĆJ�����(1|�s�����R#�Ws�
�:$[^�д ���J�� ��Fz��6
��(kr��� ��C��)`�Pp��0�BN?�9fMC  ]I�7+5L��
��li���SMN������b��P]��ES� �*�jxz���4��1{�,N��(E̙h6X�
+2zHr���п�_L*ɨ*)3��ڬX������f�^�겊�y�ƅM�5Y3km��d�J�f���KSPr]0�4 �91�I�Ӥch�!5+HR*E8�E�r���(9�<� 62/�4�0�H�dJ@N�N3	�J�a�o���+l�+��Z]�b�V4��,^��.z���hBve���>C'T�X.�̍|rv�O�]��@ʉ^�j��cF�^��N�Hi!�4|��Ѩ��z��c.��e٘O�ǛkMe�6MS?R�(b�F����ޔo���( a 2i��I��n����Tx�0_��J?�h"A��G��k�̱ɱd \�zy�ya��1�Hh�AMi�h�$+�^����9�XӺ"G�����ҫ��z7!6�d�d0~Y%��$wf�.+ܥ^.��&˒���q�e�_�z^s�w M�����;�}�t�f\���^�y���yvm��f:np�#�W]ђ�� �T� �y�xtDs��O�~;�^�
��՜�7�r]���_�d�&��s!�`��+-���ë�/I �h?- �b���[�T䜹��-B`�4�W�E�{K��z���/k?�	2�a̝�_g<�EN0�X��^K�ͨw�ߓ���Zc��u�n�O���o��^3R���o^a<��"�l�b�w��ٻ>>7��֬��L�DRY)���5� ��J�K"�����?�%r5�Q ��)�u�(�8�1�:�i2TD��k��j]sNf@���.�̩����9�|]E$4&nv[�����%)`�$^l��/>�O�j��B��/�.���k�0Ͼ{����bie}e{m��6������[�>�swo�7�<�rncQ����5���'�=#/�.�O�X��,�K�n��ܺm� ̣�xKc7
2�RJ�U�^+� �]���͜6٠���=���6��ζ,c�1$�̋�Z/u�ECh���˃/�xl��Z��@�{����Ã�ׯی<<g��z��@2=ZcL�nn�;L�}S���7v��_h�a!�I��_�����.ͩx̦��
���'Wޤ�� �� q�
�S�.�J�Tʀ!�O1�:@`���L2���# r��2M������BL_x�3@��_N��˹�[7N6��7ƫN�l֟�_<�n��E������>Z[�n�y��X�ӈ�L;4�ݬ1�V�˳
�� H{{��%Z*nʭ�c���C���������J����Ǐ�GV5����+����"j�>��3�L�|ҰjM�L3�UIC�㣛bp��2VD�i8�t�em�N䜚8�U3sYU4���A<��k����i��4�����%7&\�]>;������k��+���a�ͯ�v���q��x��d<�6�,��S���,{�*K�z�)]�Q���[��_����
U& ��h��|����QJ�6xE[�7�j��8�Œ�e�\�3^�2K�C�Z�Z/�	0 �4�������lno����*b��Keۻ�۔��y<�nXn�x������t�N���co�dȌ{���������?A��pJ��WV7Wm�~����;�mc�bǐm��-��ehxKSv��_��ZGau�)�$ZR4 �X�4n�K�M� �`Y�R�?�O��En�؊dL��!C�w�d"h��Z�����!M����T<��L'[!�����0������Նj�w��&dtV�0h������������/<��������������W�B�t~��\]�l�m.^_\�Z�ܽ����g�G߿�<?�Z�^_Uu�(`wf�劶��.Mmk��Ys_�4���6�/�NK�����������Gi��>Բ��l�M+�!����(��D�W�6��)�R�CE�&�Ĳ�C����&���H8R`�zu)���w�
�^���	?C�3�)�W\<jV�����3!�#M2$�m�Q��.5��R�LOI.60��R��q�]?�����L�;�U�*z�!L��lYZ�:\�U�8tY�ֹ0���g�V���j�(dּ̐b4~��!J$l!m�64 ��L�@��F��ᑡ �`K���9���dt����m�?���e�;���^�%�	s�g�	[2 �~���1!�a��I���1�.f�zՆc�#Z����P�L���`f�/و_H&`���`.�jzT�
ZͶ���;/��s$fz!�2�4!����^��&�B��Sqbc ]~���{	�|�kf��-�� ��lٴ*��T��,�!i�l!9�]oʆߠ0(d�1��Y��)5��p�m]z5��S��7u�,oo��:0/��<��hwm�l�jao�r��k?|gw�j���_��W�������'��m������o����{ks�������ӣ߽�p�r|~t�xpy�ۃqBP̼�����8E%!��`�/�0�����=:��лm�Ֆ�+����;{���n.�W/7Ϸ.V��V7�WΎ��7n���vU��zl>�=��|��.��^�m������iqjk����҉��� ���?��]$B� �4ɧQ�RK�4�-*���,�ͨX���)'�ɺ2��v�<ڮYeB��q!fz���Hht���[ud	���� �X&li�&5��Sl�Q�W�lN`[��� ɖ�.�lgC�9A  �b@EЫV0D��̐�͜ު�/�x�`!Ր��ƕ	fz �[���`�Ucنü�i�Ɖ	*H z2]\/|CH��C	��&�&�V�f9! �����K�U պC�0/�� �؂�e�􅝕.͐H�K˜���(�̋_����_�-Z0�X�Ħ��4:�*B.���i� 4�)3O�P&=��^�b��\;�̣h��s�4�7�0��"���Mَ����ˋZ`0�EB��*r�d�+���  Q���g�VF� �F�.�F�;A��W����&��
�2Y���ıb�dF���N`KF�W�jR���E~���� L��L	&ȂA8���bfE&��XԚ�1O��mM8�
 �x��bHΰxX)�V�mށg�4
<�x&ӱ8)՚`h�Scz	b�˜8fu�\d�4J�h��cfkT���*�%���z�){4�ׅ�0�:2ץdk17R���>J �Բ-׬ڊ�s����o�4�\cpRG#�z3a�K�0����K��WW��d�V�+�dށ��;]�Q�.6Igك��c��7N��*$%���%w1h&�����``�MMY�@��B�����_zuv��~d`���7�VJ�0�CY��co�
@��^�� lk �N�b`�FH��Ã<��Ҩ[�4H�����VSפk�R��9%��T���]��u�+�����(�a��(�w���nD�a,y<+���r�V�YaS��9�ԕ-}Q�d�����'|]�Q��Hlh��A`���Xi�uQj�4(H�E��������߹L���?�Z���E����@^#3}ە��0\�јv��ǎ��ү~}c��-?�D��C�Nc�$�=(3�[�E� ���U��f�"p�֫�"T��Kָ\�s�L�?!p�j�6 Fa�X_�� s��:sr1(h5#�W�V滦��ӻ�G4����N��� 0�y2%���ֶ'�����w�7��-$�J��5 �+��^�]g��C^�#�h���"��ML�n7b�r=ĥ�G�����j`�e5��S����ޖ1A���fef~���D���+B۔T#W���b�;�6���!�0��^M�B/�"/� �w�}�=-s��'h
�!�h�ŏ�da�`�� �b�k��e3��!ۺ\oQ�r��6,��dc�pW�]kҫ�V�<|Nze��h���k��A6L��D�jJ&�|���,�0ֶ$[ն�FJ��ǐw2+�p��͎
IM�!��ݖmzq�7����*G���NT��sj�
[B��^����V���O�,C�\#��X<�mm��iN�H���C�ʆ`0���HJ%�4M[�旞�Z��w���p!�!�	��mr`V��U��[�;��?|�na����x��5��_�<>���}W���������G�U2i7y3Rͣ�O��SK݊�eU��X-��|i� 3�C$���?$K;�Jד�=�b
�\ȕ"&<Z��=������O]P�(�.۾��v��Sl��A���R��1��~�3A����%��#{z��$|����KÝ��Z�ͅ[K>4L�y��<y���5\Z��FVn���y����k�K/��b�/�Z�v.6l;����s
Cn��4��^�F��[�N3���M��2����A��F]Z�HW�HвJ�kf�R9�.�5qx�߿�֤c�&�ֆ�O��Y}\��!�(Ŋ�K�.5���It�H��R�`���s����\{8�le|��{�������K.�xP�x���1��B�rrf��d����w�ny�vuc���M��]3;�vI��r�����v�������^DQR,�n�YF�����|鵌�6ɢ��9K0�/'0���B-ZI{��1<Zy�9ɤ����'��B���������=0�`(K�۴��-�&E���Lg��z�`�J5F��l��AX��ݳخ��h�ǯX1ŨDn�6H$iKsH�jf]��{�GG��������w������߽qcsoeku��ǽne��%�Y�؇���^��x������x����y��x����a�B���/ɔ��k�{��Iv�����t�p/tld���`g�` M�.a�.�) � &K���r:OmɺX�I2�H��d�X2*�/0��j%�����_$�$�Pօ�	Z�&sET )�j&S�%�`�\(-Wz�R/gK(��,�	y�F�D��sg��6���ݻw-G��p,��Zk۽:�
�Hi}J`�ޘpm�}��'��Ab�����E/N�����b�������n�|��k��Ct��g{F�E�׆@��$�VA�\�0�\8��E�	`�J)~��m�����E��p �GSz˶.&����5L�B8��Ν;��7l�9�)����I�b����C&�k)_0r����]�dcǈ���V��4pޅ��GŤ�����ka������|�ym��#Z]<��K-�C�1�1p��f��Y0 �%�ѡ0@�ыV�j���L��e,j�l���
�"*5�.��4dz����
M䂧iC�+�zEe?�v[d�՛�����Kkt�[��/�wo����{��{{�|�U���ҋ��+�{;���-7
}���g��=?}�s��gW���/�Ǚ�?�Wʤ��Y ��^��b6:�	��>��3��W������xi�#�r)=�����m���6��as{g{kuqɗ�O���>�O�.�^XF}��-����ܺ��7�����q`�N��T����PHb�Ia�X=����;�	ʌ��l�!��Jk��є�7Xy��:a�0#0�!3�/�� L4)�M��b�90B����´E��^�s��R�� �M@/��%�����.�a�~�3�dXz�)�R�	ӅDI 3:�4Q�R�	0��S'�0�f������A*9"��<;5�Yfhy�ma�+6���,�zi4N�.��7m��DKϖRo�i����K�iC�$D�V�bC��hg��R�p�h�5)�`q�E��.���*�    IDAT��4�����vو�aV�Bj��am1�LS��?�OVP�c+�2����B!y$g>_-��x�MN~i����X��0Q!d�6 f��u�	Cê�YL�"Z�<�s6h�0jNz�H2g��2_��&|�4x��*=M��g�A�Qɜ�t�ac�U�q�Rht��9u&@ߌ���
�R��I{�j��=�1O1��73��@JN�́�V��2�dV�J�r��V�B��@�JR�a�9����պ(� �d�!�S�f�7]��!!������wQQƟ��S>	���V�i�WA���h*1 �f���Y���2�0��(dJ�"HY�B���h�&а��$��2@��Q��a���9�B�#�����N�C�|�+�u��p5NJ�;�̙87d�����/Ww�#�q�y<kɪ�d�ZG��n��,� ��e�z'�۶^x��e�`#��nyDR�EJlvmYYY5����Pc�V��9�y�r��̺�3�����r�D�Mh^���[
�<�L`��
�&V.���ϝް�^�,}��F��D��#}&V� .@ѿ$�Bs�B���\�Z��tK�k}�ș;�(��1��|�	��Ж�f.`�i�3�aP�(y�X�4�R%6K�0f��;�Y˰yP/�!i��Y�	3��)�&���ra1G�(�e�P�vQ�쨲������(K��2�5JO�`41$��20�T�	4E�,.0MH;M4�?$,J����̀�I��0[��M8.	�dA2�yɊ<�4������G���Y���"��k��%���B<}�������%_�I��|)e�H�+���i` 
�e&F3!|�7/�j� N��.# �}�튿��x��
L.�%��!�L��f�3C&^�L�(J��)�T,��V�Qe-sUh�m�Ն�ne���!�d�y�cN�?GH�`U�6������H*ܑ��d-gz03���Q����ߠ�m7[�m���*�i�H����-2w3�`E�3��Hb: �P�\p�����R�@c�3��\�����_��M��m�5-�hg��`
/���$�i`��Di.�f��ZWS�}�}*�����
��C���b�J��*����_.�if��l��`.��04F�`\��õKi)O`�tW��ĭ���;71à��E�DB�����@
md� zx{� !<�б�D�p;"�v2_�	63?��dR�R��ɽ���r:�������f������۫�^%N/�������2r�o�������ַ��W�UZ��_:�Ơ�e��$}e��<y"�n�r�'0�s��Q,��/�◿�%�'���艴��hc�}J�x9F���SEm�X��130+dw�%ii���&�G�� ���s�Bv��I��n ���-���5���"���et�*FD����YPU�>�{�q��o.�����J��������������`�^n|��Wv��@<�
ƀV�j�U[�����  l�2��T��;~J͔s�HȆ&�/L/���� s/C����������^?H���l�$H� �b����2+v�Z�6�r$��^9�|a��������\�������R/;�]�=�ҏ��X��uĿ'�Vw�����n|<y<��2�98~������ˣc�tV����z����/�w���.���H���ܴ�,s�÷-���b�0Q�/)u���"�ol���6�#�I'���A����	[�y���7�6b�;�]d!�������2���3I����#���A0�r����kc^V�?��fx��K-%_I�o|���o��`���������G�/w۽�o~�僷�u��w4���Gv|�����w�;�q�ח_���Z`��=:X�Jڈ��y|��?7��IƗ��A�L2��K̝w;���ҧ�����kj��P���, 	�"#��>M{u���Eȑ�	�%٠�Mo�SK�d�c�4d�a,	����H�dB���;��	y��,q� c{t�(;�|yq�%@����D�J63��1"7ș0�^�KC r�e�0����g�g�G����#�����۰'���csG�v2�,J,����e�>����N^NF��
�l�&�/��p������g�81�s1;�zsϗ�.gy�Ǡ�>I,��B�PE�rNQ�+A�(���Ϟ=cE.�>���#�S�b-Y�G�iƠ-U�S�"2��Fłi/�n	�Ss(�����+�Ӝ�1�l ����du��:����d�(: ��c�,��T��Y��]�ڥ�1;@�`5c��'Gmq(��-��+."J�SO0�HKp���
	#7&�u\�M߮��� f8�R� z� ^0���!��K��;�$�]�f K=1��$̖�2`������6�;8�9w��. g��ے�c�����'� ���{�w�_I����������{��͙_^�.�n7׷��S{y7*U���4�� Iz2�gb���u)�5aT�*�Rp��7�Üx^y}o_���ͥ/���w�#��G��o�p��#��}�Z�˫;w���x}q{���޾�·o<8�_me���G���f$���y�k�Vn寷��7�SVl�`�%��0K�_�\�1;����Hɗ�>/������@[������L���d�:`J��'k�X	0K�jؠ7[v�!K��	�����`�aMo.h!0Hx�(0ɔ�����@b�L�C�L�$ǁ^�4�&�P0fJY.f�8��?�p���9�s�!�a�� �!;Lq:F0��`΅�cKs�I�E&S��4(^�I�$pi�Hc�QG���/!ɓ�b� �����7�BDK�����m_�r�A�[}��)�4pҘ-��/(�W��S��	���愧/hsA���X�̹�
g��!T��(IJ9�Pl���	"�#1�Ţ����!i�t�ZF5i�QcTFiO�zR2�L��,	|��-��8	�G#PV����L|�&t ���FD�B��ͬV2Sх�G�ZPBr0xz9��o�/z�s** 2$��"���X&�F�4%�,���bi��TNd&��Y���4<g��i �,:S� J^U׍�4&:�1kGUb0��Lc������uXa3L̐���K�|eN_�&r���Q�עg�7��r����|�eb�DB�$s,D���.� � �1"��p-饧!zu��%�Q�2�V�����Ks�͢��Q�48���x���A�]9�c�B�u�&f�����U�������Q���!@����'��\BF�s�<H,�s����7X�+�	�QWYi�2a�B���K0V���z(4�rl�7�b2`
Qڐ����*�����G��_����y�<���-J�4�8����Ҥ��c��D	`�g�.r�f�Sܐ|��۾�\K�+0��:Z�YU�4��'����Jo�����[�L���z"��C-���,fi��Bϋ�����Ai9M	�R�2��[��/:%d`�*5P��b���@�dVɻ��OH��&�%y&��"Ӑ	���pJ���!~�Yi��y��4�)�-!�T.�j���.��p�A����"���)��\Dr%3�4"�^&)�^!)��+�c��d�EѨ��c�賛n��Z!��$����\���:Stz^L)�+
/��l�dͬ�
�IT�,�h5/�����[nq�o�y��c�
x�^
)ni92�9a�BX�kȼ�Fƌ�,\�����.
���d�[t�����$�F��0C䎐`G��L���a�aF��a`2��D� K�!"G���t�
���[p��ݻ��a�48��.�>+M����rUCҀe5O�4|`x��8��Y0�&K�M{�}���y}nW+��	� "$ǀ�f6��V�������� �G29K>�\Xg�dxK<d3pJ`ǔ�d��"�f��٤���8L~�t|��/n���O�u~vy1l�;�g�q��7�h�A8=UAe�H^�D�j� �!
��_�\P�f�u���b�$_�t7~�_Xz�Ժ?��K������3���
����u���O��O*����u�Fn�9��Hh��p%h���n����=���I�p�rT26�DV�nʄ;6^�*2�˕��.z����e� o?��E
L�.G6���������g��8���;�>��潫���;�W����f���×�׾U��^KE��r�C/�YO�0�9 L/H��o{�p¨�#�n�E6��L9��rvb���E�̬��&�	��]�^8�M�h6��ȧ%��kw��Hk.�Q�@���#ܸȍ���z�'6��<�O2�K�_��+K���#�������j�����ګ����{�/�ݿ\�|Pw�·�m�?ߜ~q���ޱ��(�3��USζ�'3��ΰV�Ŵ�������)y�q� `#��㡛���ۿu.i��݅LM����-����'� �;�Ѩ�ΣC��ؠ�����2����/��l�[:v�8
��u��!(������{���{�a���~�m�#[��?��<�ܜ����ï�'w����o���ww���w7o�|��������^���+Ǵ���er� ���x|����;�|$�Q�u��?�Q������8���76w~�����h|U�j���>m��ũoR�4�A�KIV2�1��I	6�,��-�Dv9��h{s�1�/����qp�e���1,��S>1�L��Ր ^0�9��SW��!}0�%$%6{� �Bi�eTZ���oN�� �!.L��s����.�Fr�b9��0�����c�W��<1�"4��x�q-������u�xlKV�!4����)l�F�\Ei(�$H�F��`:�4d`[]��4{�����&w��7/�{��eF�Kpʀ���w�H!v�뤪ES���B��d��Y�RU }m��#Pg=Z���\$,=�08�`Nj��i��~`G��r$ &�G��H�!=�c���f���ĝ̅oi����@H/Ol�D`V	pq���!���l?��K\m����B:dR�����
�$�m	�D�e�PC���/%���뛋$0�!7Q�+�ȢǉI��p�� 7A�[�R�9�Y\z<Q!o�Z	xd�P��/��Y�|+�x���v�+l�G�����f�hu�<��}�>}p�+�ֺ��\3���_y���B�.�.�0�ry�wqu}�{��܄�|,����,�!t�W!���U]�j$/U��������W�7��B�_���>��O��nO�֛����s��e{���9y󭷹j��lwy����qiܻs{��ڬ�u�[�|��~�e|�_��3"���N}�F��i�d�UNɓ�$_�k� ���C������ki.P��>�Y�é���<	�!�NyJ#X���r�K� ^U::�4�l�m�I>����X&8a�֕	 ��f�/sx?� 03&i4�[�
��@��L*B�BN�P5~�r�C5RZ��G[Vf�C�1��L��z2���O�'Y)�O'�����w���:@/:�%I��(CZ�sA��b"�@��7d�1yQh�ȳײ	|��������j��j �� #�8�@(19�O@Vl�n��� �z�@Y�J`���'�-Y�d�%$����.����a�U�`�`fC�B�s<fV.|�p�����Tg&Cc;k&?y�ف% *2~K2x�Ē'�U��I�2B�N��J>�2��$=p�0wY��+G ���Ai BP<4�I[��Rj��DIh���+����e�0�-O���Di��[�Y�!Dsx9Xs�aʚ�S	���;��/�"�if2��,����f�2h��`�4���y��vrŚcC��#����L�N_JVKx��Ec��ʐJ�Z#��!&[i�p)"�/sxV���G��đ�>P��-0<�(�:�Ơ73�Y� =6zۦ��(�1��@��/��l�lPV�t����(͖�ɐܽ7�F�Ϸ|h�/�C�f��3��B�Q�4�ze�5��>7Ӏaf���ˡ̫T� ��[�b�L\hX!�4~�j�'P��W%��FKd%��L_D�Q�0�W�3h�L\���һ�!�l�Ag�2�\D&KHi��d���v�'F+��f��@S�4�	3#@	�<Q86�O����ȷ%�ѕ�!7��_8�ƒ�;�//KB3&�?�	pl�a�$)�(LH$��A�O��~��^p#<I&6�����h*j���C:+g9��#}��װ������_�nY����%_���p�дDȋLp-�>,˒1˿L�	�(��>�D�c^L\X#�\͚,����3:�^�\�|9�%w�Xe��!�#��5��1�`f]�82!L`
)ɘE�=Co���1�>��b��U�f�Nv�����N"'d��ƌm� s9�L��4s��H��f�X�u��!�m睜�,�B����4Ə
m���E��4�S�$�H#�Y���
�հ�i�+�k6�:s��3=�T��Ss��s�����.q���L �K�L����\�2�L �aE�����$��b�UMvJ�Ϭf)�d��G�МZDCna��i����e��i0Q0�D˰�߬�ܝ(�v��8K ��3%C�R����D�Y]p�/���K��L���� @,~;��� L�	H:@���);L�b�yl��p�c�a�Q�8���L��x��Р��������&��s�׏*����0�`s�=�r��[���	�۹�WJ����+�.,./ ~�RI�  �1T�����#%���QO�<�裏 E��L>��[������&ӯ~�+�-�W f&�Ș��>{�̣7q;���&.n���Y�)�g��KÅ�g@x\۝jy�����,�����uz��ԭoL�;�������Սn{|�F�K�g��`�^�6�r��f��b] Eo,�qM0�0���>/��gY�1H��Ru�=K����i����[�Z�FO�:����:�3�����c���M�˶�A���z��!F��Y)�Ө�����r��������o~��/�(̗�o}���8!���)׸���+_G��x�~��-�k���¯��y����z��W_���Y|���Ɵ�o~{���}������?Wd�"�⶷�p���dnG�K�m��q��>v>�!mu�B����w؂�������9%�@�o�6:_�6��@�r�";R =�� r;�/��/]�x��!�[+�Q�"-�l1;��4w�8��D� ���|�9���D�Y�I��c�.�bǵ�����ד;��.��<I�n���׿y{���������	�G�~eӣ�/7>g��|!y5�!ѧ�|6sy��2�K��w�����'y}l���dw�Z�����q��]��I7�>U�9�q����B;����d�k;���P%���cH^v�KZz.�y�2 �LY!�.U �����4��'�j� ��F��V��SN�@h��l���z����@X-�dC�4�0�"��x��E6�6���R+�.蹸�{ �G2��D�%�v>�R�It�4��s�V�������!y9)�rA��_���L�g�Q���5�%Y8:�Ki�������z��7���X�3�1𕶥(=�?=�@z
t�I�|玹�%�_DW�ٲ̀�3�*U�Ҹ>@��+���XeUh3=BWY)���Ǧ^`�-������z�U��e�D�/g�\+0�[�w��X�	��x�(t&����Q�]K ��4���<��#&L�£Lx ��ܾJ)(w�n�b,7�=GS[��78�+���#,�#��`2�fVB����	2�l��X�,	Ҩ�r���5�|h��L�!����g���wx]����98!7���ַ{o�~���ܞ��8X��?��z�л�?�7.��[��<��R��B�}{EKL��o�-�ebI)�T��1y�Cց|G�^l�'.o����Ó�ћ�wξ���_�>?���%�{k�,}X���J��y�ǲ���_m��m^�J��k4���|��}��w/��z�����C�\_�n����    IDATVcG�GD��lVB3Y�����3�c��:�_��L��a(��E�0�0R�i6b�B��%�l���%ad��X�-L�)E)��j�l�ٟE��XU0a΅f�H�sj�u�L��L.�1i	jaBR��)'>��/+3e����E���b��P�N_D3V䬍�	�K����K^�$S�k�&�G�/%N�
dih%2S$�\A�$�i���D�Wò|bc�H��I����� ��^�����Dȅ���e���r%0Zs�dbF(O�V��e����)�Ĝ�F�= k��0\�L��N�Lh*'�4���ҔF�Z���'3M/X�)]]*��Y%_`�%�,�q��)��`s�'d*I��y$�-%����i3+���ʳ�aʜ�,�rJ��;6J�y
���=� rT��9ڒ�M�R�����\��Fg���i�` �f]䒤70� 7PYR����\�r�\��y���gJTd��l�N	`Y]E��++Xz�F����lƖ<�п^+N�PJSY8���$JKYYrY��	E`%��$#6J���s���48b��\���-���U]h�7��!x9.� �Ҕg���@��R�θ�Y�-��˄����r�	@c `����@��L���f��Ho{�8��F�a�ђ#=٠/ts9�A���I�g2W��dTh����,��YK؜�����]��s���FT��S��U ����4#�W�����d�o䅐I\#M&���E�:K ����EBO`�$�!yj �M��K;G�FBi�5�$���;�m	Ƒr�x��#P!Ж6$6�><�3���R����q$H�2}s�c0K��ܪ���}d����f}�5���i�La��4Az��<4K��s�ۨ��Ty[��+T剙LY�r�I�F��Ʉ�1��x��4K������2�t���F�����Q�RSU����4� $63L��,1����
i)4��c��#Y V�%Q��YW���c����I�D�3OBJ�����L
W��d�F��@0��� E�9����ӧO	:����t�RΖ�	��g3�ЋE�7�$Ą�,�ZDH��of�����А�/��s�R8C	i�Mb���p#�=V���@0�Hh���Z3�PVd2e��қ[�k�� ����^���z����7�`�mtf�G����t/�Ʌ�R����%���*�F�x�f�o�h�y�Y�`|��x�7G�~�\����6|�1ã�66/��!y���Y2�K����M���"��� s^�ܢ�䉆���5�*x�!A���27�%�p\f�|��n��෌�\J��z93
G�#��K���~K�|Y	�O�eQ ��UV6���כ�l{}�`5�1���������r��ރ{�=���+{�K;��=30N���2f��e�H��H��JE|��[��nx��?���mi���UV�!���>�$0r��ӧh�ˢ�ة&O�V5�H)	����?V�Ĥ���z+C7'��9�.qn��&@���KUtr�Y�fQ�gF.%�A&Ґ�M�d���{O,��Z�&��;U��������;Z�g>���N}���j����ة��k��~��3r(��^-B��kDH�l��`�Krsǋ�`*a��q�+���G�Qf�^M�3(��x��@M�Dqd�88�t���V��
� Qs&| ����H���P0�82��x�40��{���W4��v����W�����O����O���7��!%mn\x����7�B��z�`���o�tw�Mӣ���{7~�k�+�.^^Lcu�=$��Ay*���n��H�-��UꁥB^=ip������ѣ��L���8l_�����.�읟G��%�?�O�$,��$z��._��cs���M�4���^P�Y���N�Eg);^2�-�Y'Y��1e�|Q������b��YY����,}w����翹}��������5��立/n\K��;�/�'�V�b�G�����ϙ�#;��Z�����ӝC�����o����N3���K^���ِ�<�v2aj�,;myU%M���1V&��I�̐"���!f`T�h��diF�|hP.��Sb�)�%#�4�1s�$�rg��+=C�f��=,����C�X09�c®�)���a�����Io�u]�]�GyK�v5��v�u�{�qe3�iB�'��\�8�eeK���v�JU,y�s�rqe[�x�GzH���v9p��j�B	`�2����,�T�H���Ȫ�C�x�+L����hC\�>��R����E����w��U����$c �$6�{�;_'>}-�F8W��K[nɮJsR�(����J%7�eN/4�+�Ш��G2.)�([2	�J�q�tĵ��]	�� (
�vh\-qrT�#�@8�`H4F&�o ~�!%���n�(��0[�.��|%��T'=^��������5�q��/�@rNOi��iV��,5�mf�n! +��mIF���8�����W��ț������������x�����Ѿ'vM����lw����K��|��SFW��Qv���n�>�9�p�����L��P���$C	$=Mz<bx��c\ |���������;�7����_?�|��n.�����W�z���/�O��]����շ�^^_�ߜ;_��7{�I���w�z��s�^���xl�[��ǟ#�W7ɒ���d�l6�̞�XB&�4S��Q �!�x��vJ�f&��	1���f-"�X, O����9wBǋ`��=��̅�`C&[�C�A����^>%6�q���H_EfrK3 6Tf����ĳ�g2��).@�0q����?��� ��K%0]b@�9p9�E+��4eK.�d� %_�	U*�r�l�l�{8��6Z�c0cKF�2��L�Aht��cCe`��3�er����L7T��� V=/(�f�3�%*V��\'a�ip�刜��(:$�ހ̅���Nr�9�+*}r	��P�6p��yy�Y2��h1��*Cٵ��͆�ˊ�p����^ɔfɗ9 NV��J&�ns�4,a�5��JxH��gd�]7 
���D����TP�s�ŭ`�`H�J�9��|��8�R�t,��3[�1�#�����1/sA�B	��ȅ.s�%�ߟ��IU4�!@���)=Kz����In0���</z�`L%VД4)��3c�저Y����r���@ s���~�m�'�Q&Lu�@#f��VufC	��Y�N.J� ��g�2�2 B�� ��0����f/"᳚���/0d���9���*I�Xc!%ϫ������i"`0st��ï%#V�`L �WXJq���L����� �jH��4Aɽ;��h�(o����5��%���چ�Co��3M�0I;zֺ�r�ଢ69<��	U���+s`���Q�3)p:Z:�lL!J	d3�(����`	�!Tl!���%_q	�#�����������7����ďs^$��*�;���(+�A��!x���W��5s��X0���,�(��b��X8Q�2��d�x�	�e	�'��	8�(��% ��}�L4��7�����ǩ�(e��7<:�jfy�g�I�b R�U�2! ��`�E�}���@$�t_���{��9�.����L��6��HB���=�v��x���iiJ��yyݶ��\*<NK^���h��.n2���ѫ�d�����(��aMcLh��L3+"�bf*��lL�`��F$2�å'm����f������dN�� ��.!K���,Y�����TĪ�H�I(���S$�� �	 =���L�O4Y��2�d��BYu��c�! /��f�&k	Є�L#O��-����Q3[�ް�mu��qG�����<MQ�b���J � \ �jwR���&�$��M3rH��1/���K�Y-��%���UEý����,�V����Z$�͊�?ͬ�Bf,qg�	|b�lI���p3y��}'O���rw��.�F��g�S#�-YU���h$��&��&��e��vʼhJ	G���_�V��� �)���N73Yn��=�qr�ӵw�6�Sw}�K��'��|��|�!�/����+�FVnx0�"j�<~/rh���Q�Rr�m'����s��;Ҟ��Yr1�4t�=�iv�3?�O�T2N�� f2��������G���i�6�Y��g�8!��q"رbiQ���Y���
�ꜛdɨŲ���1�"��;�n�Z>}������O�<�@�����g|�`{u�BO�uv��񍤾Q�ʭO���f\Z����=�r�'5��]Qf�����#�F�6^ �(*<�!U#%���`Fn	���g� �*�4	�d�z� �@U&ܵ�G�h5E��s]v��B�9�������3��Q�0�KŖ��ҕ���g��{W��d�����!쏿������ԭ[��Q��`�L�-���>�y�~�b���Ϳ��l}x�h��7�o\�l��|u������p���%v��h��!�J�#饭�c��}pz�Ks�*v�n���k�|��3������n�ٲ�+:f�~;�{c�l*����K�ܿ��:39:�=z�JZ�$y	4�"�%gV��Ϟ=s
!�E���� N��|��r��ͼ�!p�Q/�~	u�l����H�|js�Kgo�n�u����o�w�g�u��s��������~���d���K��?X�P�����z�l���T�e�Ǡ�����+����S�[O}��n��R}���o�x��a�2�'1�s��42�4��� ���}[]��X���R��%��!+=���Vt&z$fS����̐B��K^�PxJ�����I�$�4�f�3�`
���*rAΫT	2���!�fV�	(���o��h�-?~썅��R�� �ܰDU�-K������3;����������UP�r��Ȣc����dcW��a�I/�/{�!���m*/2q&
$U2/BX&HUVg��]X�W&Ni+M7Ȓ�R��J�8O���4tt(e��u?�<�$"����	��!ħ�~�k��*��/6�9�E�
�����a)�M .sl\P�w�J���������R���T�j鵓�<{Y��7��@�R������Ri��Џk]=a���*��hPv5���F���/�U����_�>�"���*E��(Y��C��=��E��և��HV<Y�:4ͬ�d،�?r��Ң�f�;���������������ju�����n����đ�x8��8�W�q��b��xu����Ԣ�0	a�b����@I6��O��[E�\�¾[a��sM� ��V���bu�����'o��?}q��½��l�z��؞n�l__z���m7���✧�^��~�{���|��7�7��\�+�(����P��䯤�F9[�p�$C�ː`.�yt#��Ϛ���No	&+*�K��	���{�?X���1p��LI�P �Pί��8vY3*�/��Y!�Lf0K�	ӿ��:l�۱�;�"d��]���P�iJ��4ʐ��$C���8���;l� iIOCf��Z���7�U
�E��Q�&z��' I*Ҁ,%�T�Wd^�H8�\��D�Ɍ*�\Xi�T$�Y��LeEI6��E�!8:b�RH��c�
P&	d���ʅ��B3��i�'=�E7&[�.�Ԋ��ji�g0�Ұ,BiȊ��d�5S�>�E	�$�:Fc��	lɄ�<�Sf.�X�f��N�zN^8F#�!�ZЖЮ�&9/���!�h�Qѧ�$H dq�8�!�5��!-�y+l�˖���ʗ�#Yn`3�Jl8���q�B���#�1��(�+��\�h̢�s�:J�QV~3 }̂� �g�
�A��X0��4 )�$��`&�X9ʿ��p�W�42�XEf�a�#@��DRnChz� ��X	$��*6<_�|�T�%2�䧜H�: g�L����e�Ȭ7~J2*JKJK�����w�[0y�MV�񧁴̝���?��^� �L���G����nl��Z�s9@�7`�UGV��2�%��$�
�,UVz�K	��$wJ ��^�܋Ȥ��s�_�4�J�L�1���@�},roG�+�������!�_ V&I"���/�i�!��H�/3Z02�A��L(���S3e��XG'kl���	y�g\H2���%���#4C��e�m���}-�AJL�3GH.H:�`�n�*�R-�Q�EA��[��K���F��4S�
$	���֒/���Y�F�h&��,=|���$��-a,�w��^D���Y�?O�_������P'��۟l��:健�=3�yig&S�Uh�E$ДR�L@U�?pBZr0��yS��_-w��&IJ9k2$��/�檣P�Lu	/r�C%�xˠ���JOV%?L	�%0S4\&'�pfJ�B3���`ʐ�E����;f��� ��/�P,T�6��LfV3˥��S Q���&;��GM��O>���{���e3�]K<hc�a(;37�P����`-1i�po�k�%LV���]���!p�DzwZ4��Q��J�s	����k�(�V&�B`(gKrc�3J���4��sѱ
�Fii H�l?["��'m�&Im	��ϊ�O���<fR+�#���p��.��Q8Cn�W������JF��/*�`2�J���T��f���v��nk�&s'k�Q]qr�\r����U�dX�Ӳ���Q��+�k��O"<ԔZ���
3�%�s�������h��C�/�`��^�dJ0��ӳR����rq�<�dS3<���ד� 6K�(�L9��<�����~�~�|�ѱq�b|o������ǧ�W�7�x�.�R!+�>�'{�D8��3�7h?�</�a���K�t����`�����)�"wb�qz	�(_Q+��%�.W!A��\�A=׌P�>]&.������xi�eEz΅�Bn��]*�X�y���������̧ڔ#($N���G�h��s��&�O����ĝj5bh��z�������.��Ϟ�Q(�����k���Ϟ]\��8���y{~�_G�-V���;܊�	e��R�U�Ȅx`���^��\2$Xr0��kQ HA����u�i�8ic�#nʻq������ F GJC�^�1�L�����Ǚk���6�a1��;�ucW������W��c��s��q�����}��g��n�wN�]�� �o��������:�:|~���������s����+v�f���(��"%��� �٥P��	��m�6�ay��(��&@��K�F�	:������~�왶g[:���uJ���0�˿��WwG �w{�)$G��Q�����S�sJ}����{M5st��}���I���`�cp��(Y�ba��@�<�����V�g���\m}�jo��{����͇�t�M�xs��o�?]ݞ�����
��]�t����ӗ9{�ve�[߬�
���^�}��Ϥ/��<�ex(��M���嵒<�����x3�
{^:����lB��,1�h�1 ��^�qdR/+��N����L�&klf� ���L
��Ұtf�dVq9�����."r4Ģa���)�˓l�\l�^̐K"�
`0;�#% ��I&g -��\FZ뵍퇗�6��X0���mcϘ��"
0�7y�b)=����l�� ���^���[^{��d���
�XNx�t2R�� �N
ѝ�r������lm-V^�X�Z��5����IQ�%��	��-�郶�	��4"
A6냺�0�Qt�st���w�B���L\/�02�.�FY�5$ZW/�\�u�� ��'�Egh4�������_PG-��Uh����>��(��ar���N`��R4���
!.���x6��ɓ'�U�
!J��K����.�ͅ�@�G���EP&oz8�HUK�"�(1�ȳz� �p�����L٠�Po	�0S�6<%+~��$404��ty�FJV�ſ[�E	�    IDAT����ˤ�����9��u�`s����/N�����x�
�u�wx�y����O=�h+�%j��-��K��P���c��0������F����t2��؆T����js|����o~����/��f�K���%b�]����W>g�Y�u���r�Y>|��+�}������~���?T�������}E�6;����d{���`I����嬟-KXz��f�jI��`s��ږ0r������@���Z��� ��$g�JU2�q��	���'��(�P�P����L����+G#�ir#�pĉ��l�f(t�\B�*3����a��Ҡc�k�$�ܦ2dI������d�X�[��Ȑ�E4��� u!�  ���1S� �$���僜�\E!g�+ �|�^;����W3�9�p)O�
i�v&xT�z�5��@���H�ѓy%TLQ����
�%�~vu%���d�pL`"�h&�,Q�	�� ��82�K~��k��$�J �3G�4 f�)�f0-E�(D�d��{��.Ʋ(�;��#�R& ? �4B��F�+��� �	C�� ,@ӿҡ$0q�ofU �A�'p�9$�] #7<�ʐ�LO(��!)�U'˚�� ���W�0F�2��_��Ku!�2��fS����Vf�a��JQ��X�|`��AE�i)n��Bs�l&Odl4r�)&b唉��" �-B�r'�jYPK#�R��{=�	c5���A�T\.�50�9ưlV_z�1*�Lc�+0�8���2�䓒#Y
G����m�x ��a��
]�31��H�Ho�3k�r

F΅�l��� �� ���$��'}�;+w=�n��{f�1pD_ڕ<�F��nX�ީzC��K}[��Nh@0)p�&��bˋ<��u��-�Um)Uq+ME�3kM�Q�4�kT&�Qϲ��`�2��ɬ��e���e�W�C�?p���")[K!�b2(����ъˤ|����ɲ!z���A^P�eHlN �|͔A��:~یL��2�<�%�YY��� �i&�,�@r��6I���a/iB0�1�dz&<�#t����`���+��v�����"g��77g�X.Hʳd���%_3MQ�Bee	�#=�ٲ=�.ɸ��jC�LfH�;�dꆸ�	��LZBQ���'$	�0�FCHY�h�G*p��V��Ȝ\ $0�f>ظx#J�"_sy��qm!�����Ҹ�I��*�L�����-_B�Ҙ ��S���n�%=/Ki��쮈!�v��d�3q)�%6V�Д��8� ƒ¸�,K�P�x�LYu`��1�hP%wD(ӘY1����$��WuwT����mr�v��o�Ϭ��*�%_nfQ 2j�eY�3���,x	���z�ȍ��ݖ6�N��C^�沂I�i�l�FU5����^2�"bS��u��tʃ�%��BZ�h�	e�Li2ǯ@��ԥ�L�qG�m"�vۍ��Ռ>��2�P�� Ȑ�)kT���3�h4]O�f��/~�QJp��[�tɀT��a$o� $�B�T��ȥ�|T\B $�)g0���ki�zB Cf�
J�6�XR���g�[�&1	�L�� ��ūS{|�������*��狝�;����<�7��T����?�C;����I�Τ�Ew�����YR����л�]���N�ly"�ų���2�(>��4{��C��@���f����pv/W/U��!H[2�,��=����Ox�"�@!N|�����]eA9j�����0w��HF�p��D��;���ʥv����O��g�&��h��k��lڋ/�E��z����\��h������rtn�%ڃ��s}4�~���)�*K��r�1��,�� �7s4 ;@�mX�B��W!�y᧴T�>��̪����� �X�y�ӽ^�5y��e�&�S
�wl�r$������a+��i�A��F��$��������m}�7ɺ!�x��~��g�Ǘ�ғ/]֍Õo��YϘW�k���?������	��9�\�d����_��;��y^z�G�Oƿ����Fi�K�2qfj�fJi������?���{�= ]�u�0xp�f���˅Ɇ��k����'
���9	A{t_>�(֏>��a����Ĥ
$�d,��b���S)9F��~�'�����젺�r����r�=�Wt�8F�������%ó
�H��:?��g����]�;<���rr筽��z}u{�}�˓�[��o������p��7�Ǉ�V;_:�I�;خ	v�#��=����;r^���8���ww����������m�M���ZԿ�'�s{L󫝠(�������D��l_�}x�������̬x���o.�e�������C�$`�:oGh5d. �����E ��"�.�dHs��y��,ܢ@�1 ���{/]��rP�6ҳs�<At�l�I���m&���M�۲B��N��+.�%�%06	 ������o(Y\��9߫$�w0x�_��S�(9��.�iEI�]�3���x��Y8'Z�� ������r���;�P�4j������2���_��vb:U�*[�0��}P/s{C�L.Y^5y"~�|50]�L/i�U&w!�)]u�I>�X�{����I)+0w	Ã��戢(/��d�^�59�KFg����@8�Yc�f2��/l���L�����4?��S�J��b����LR�̕�XK�^�r�+�(�Sʳ����c#А	��N���L��|)i0s���R&|	��Z`���`B���{q���r��N]B���!�r��wv�y:>� �����k:�-Hȥ�KQ�u��Uh�s��l˼mV&��0�\��r���=oaƻ��M�k��n{�_����.���}��?�����yzy~��=/.�?�Y/_#��R���܎w�������[?������������w_��'���\s{{������^y��Y8����KO�a��$O��X��S�(���z�#I��dVHT|s�C��� 9N`��XN&J�l�t\������5/&�#ɷ@投����;�XH���F3eBI2���x�IoXV`< �M�b�
��q6v���,+=_KV�)	-�i,	�5�H&�`�hD1R-��LYV�d��2}<N�I #��)�"И�gCh���n$�a�V��dO ��,c ��(kNC(l���y==��f�853$����ه. �.�����.V�a�5r�հ�B,3��Kن�^�9.c�\��/�����i�d5"�wJz�<�%�4�,����lν���`��2�lE�E�B ͼ�L�ӛ!�£��?�D4�lX�3d&3ߺ�_>0�`B II_tx�,e2�eY1�6f�[�T����1^�V���^O��e�r��Ɯ�l�?u�-6.�K]�ؒl�ON^L���nY�[�F &�����Jޠă�RPKʂ�[�g���u]�޻36����>NT�p1�fJ�d�r+�@�P)% �l@��
J9#�ULx����]�����-%�f[ƈ�UI��EF(7���ɤ(JKcv�-SJ���!L$f<4���3��;S;�IJG����3	7��˲�ӥ���!�ǀ'A�}��.A�PE������S!�^�r�֟�|ˊX��Dhـ0ㄗ�C�ɒޜ��1�L�����/���T�԰�K���O�RJ59^%VE��>���Bx�UQ1s!�! �=�%�NYP�./L�f�X�k/xr��5�=w&rz$i,)e;�,=%�	�Ez9�*�ت�$Ȑ^ ̬5�����o�h��H/�4�.z2|�Ж��d��� 8ve��IJ�������h ��r�$�W���'&�t���7������b��z�� �P�"�i��2i�B�@�C���O���̊<H���\��@C& �a&Vn��4����c�(=^��'ē5/3���fQ�	�s9�Sᘢ�j�+ܟ���ni�~�4z�R�AD.1��r���Wb�-G�jt뙯��^"�?���Z�fzJC� ��,�Vz����p[�Y7�K����  ��zJz��!���`	����lP)���m�L��m��>�8f<4�a
F@��^tK��,!�ӻ�S痛6���U�7~w��eX�)�\�K�Qݒ�ȜF-�2'(��D	bIưd�!�qr���Y,^�����I��R�j�3��̬^����r����99;X\�c�F�f2G2�%���R�L����J������X6�ۛ0��204b�2�p �3�Z\��0�\��|2V9���tX�e���[cB�Ys�t �[D��)�-g�49�i����AJw��^��|��k��Y?6���������w��z�|�]��O�y��n���Jixh�z"���<r�PD�w�nC�6���Z�Y�>*G���sw1��ͳUx&�a������w���
�:UoϞ-�V+�_!��}H.�:/sK��,Jw�E����9�NT6�r��.%�].�N��d�Yz	3�vfB��i���g>3��ŗ�߼wr�dϛ�վs÷�-��h��ק�����v}4>G(����g��2TBH�<ȺT�
L�t��O	�lv ,́3���Tr�1P��pw������Y�'\�=[:^Z1~�4.M�#��.���m�!���
Y���%Le����G���GP�'�V뛋���ɑ�_�sy����Kie�c߷�������������t�4��e>��z���]�ܜm�/�o�w7^6�;_���o���~����	-9[�p]�-��N�i`l;�ҳI�q��� 	< z0�����u��?�)Y��a=5du���������9R2<J�#�����d���}���`����;���瘍.Il��:�����8\��)��Gn�-=�0{�������{+_F;�����/��u���������ѱ_E���z�=:<�r?����#���e� ������g�]�޴I�k;��m�@�G�kS��>���Q<8�o�K�	L�}P��|u�8"0 f]U����n�A!X�;(f�y!Ξ�U�L�q�^�1�D�8 *[�^ ��T�j�	 �$g���[BY��3����5X'xs�2!X�Yb!��+wT��1����c.��	��)+��i�C��9��R��J�*gz[����io�h饅��]Vܵ��h��\�."�= �����<u^28�5bI^h�y�6��A-��{�^iKǜ8���c���y物ˋ�^��V�J��Ź/s�j=w��mL|5!�z�\:��� �3�Ft�r����Y,[W��w��䎦�]&�~LE�q]"��S��p�V�jG�Ip�aQ�ƊX!��4\.\� tX3Y		W�(�R����(y��`������GH��EZ��iQ�Q��[	3�V&L^��G�Fm��w?*u��fC&j�{�p�ze60�hrzx��4�JH��4f��aR���>���ug?�ם�k�Z�I69�d����&EZF������W��7=�I� ۰-yу<B�bs�����KUfU�|�~�Å����s~�w��f潝Y ��Ax��h�r��Oʮ4�`ݫ�ܑ(�P2f3��XQ&�|h�\D'`iRBƆ!wz}���
����`��w��N�۱���o���On�����/��z������$��cJ�t�x�{�z�rw�ko��?��7��}��W8϶��~\l=��Z퍔}�S.	��"Z�49��-�1�($��u �� ��g��@�X�90вi(��3���k��n�a�i�:�d)e���h�HK,�d�� ��	��p��E(0Q8���#匕������1��-�c�C�r�7f�6a`֔	梴$3�Ѡ)=G*ߢsI�@��0���N_�9�E��9��LFu�ˍF&0h�rK `r�[ �U�A�$�Ңqa���#�r����0��cD�4���_C�K#%�k��Y�0��^M0��4�X`��]� ���-LV�z+
X��b1����9C"1c+2kz�-i�����f�� ��f�2�f�2�� ���Q&L4���2�'fJc�.�܈L6 䪘2=k�9G[���9��W�0�RDe���X �]�*�ƒ/*��ϋ�9�� �Kw.���C��S�BD>��&Hy�͝���1���
�k��Q�b�I6r#���z�BO�>*�#NC 3��K0�1���!����+�7*-�%	×K�fz�%��'/��J��l@���NF�E	_�ӗ�K"��d�L��O0�1�U3��A�h�����@�)�L�S.Ŋ��ɤ.<RB�(��L�:^3�ɒ;2�B,�c���6��D/1� ��4�sE!�0J��B��뭥l 8��4Q�Q����h)=x��[�>�KR������z���gd�l��)VK�CZzY�Qi��%):�|i
Z&b 㜻�����Koƃ�lI�Ӡq��6��$���� K�2�d�K�r �D�!9<6z{���e�l�Zz�4�e�iPa��-��*��;%���F��1q�xu.C&�D1h 0P��6�!(k�.�ӝ� �	�D���=&����X��0=+�rrr�1��I�d��KIM��J�ձv��ۭ[��|H�QT�:c�1��4�B^�fJ	�tӄ�h��!�l�F�Ϗ�pY��o�VՑ�e��d�a���s.��VK	�-�a�Zd�ՉF���g2p�Kc�@hɷ|���i�n}��!���P�"Ж�}}���~�H��aǎ\,�b�mϝS>�7���?�$�*�^���I��pf��%���@l4���cLs=[�:c���p�!7c6�>���_n�C ��Z*�� �*�-玊�mϗ<}�����EwıI��꘸�����^,���fǷ#ҍ$�3a%tiE˗I,�o�k��a"H����z��|t�6�(�@W{�
�X��-'%��Բ�� �G	%<��3��L:I�����-_0J�Z�d�;@�X̖��m�|zݶie��:��fA�����i���	��U�gi i�\��FGs]�O���2$��`݀De�o�\*~�o�2���J@K2a���]4 _�E,3�QJf{GI������`�W;�^|y�߻xz�>��ͣ�q�����s;����j'{�Ɏ��
w�T'��;"��Ҩ��ݻn�:.n\t�Np	�Vao�lW�%�5P���h2�6������L�B,0�r.�E̒1s��dx�i���%L�r���zB0���U��\��O���Y䢼��{R�����^��ݻ�#���l�Nv�\8qݐ~�Xq>~�ů��7�����˫��G��\�������9�8|���������"�Vm�3�Ȝ�UR*�`t,a,g�'���l�I)�(�+~9(�R7���4��F�z��h�����XY{0`h�&BhSG#gyCWUK��bGm)��B&zr3���Hl.^��wzt�	���s飪��\~�y�+u�X��dmg�[�W��x�I-�y㧃������|�s����G���|����*��E2겙d+��Jz�-�T��ΰ�8R���h�&0a���w=ۀw�م4�hO �Q:����)��b�:Ndg��KåD������y�ak��:O�\�o}�[8e%y����W%%����T#dGMP��#
G���
��~�R4ңT�(~Җ�ѯ&���ol���
��X��NOvn�������K�{��v����/�����3��$���A���2�XCJc�_���r�9_���t��:�ܚ���y�+;m��\�=Mx���8�0��+��%b���	�H0ڬd�8�rd��x�6����'����c.��!�P:Y �M��o���,�E዁�Ti��N���b6;d�1�q:v%,����q���_x ��"<_0�a��W�ٱ� fo�'?_`[�*xu�$Bx�����q
�p���x#"%^�����މ �q�:�4��>�XB�T!����W皓ι,��Vg+GJ�C�D��k�*t���7z9�����̪Xz`����{�,m�EH�p�}�wD��~    IDAT�t��L�(�:/��i�M�z+�������Pi��n߾�Fh`Q��=�6r^ �a��HS������j�$.rC���zu��4� �v)M���^\Ae�LlG?@,+M+OH��ex�Q
Gk�Et̊� A&�é}��&�,���ɹ���"�X'���K�(U�m�$0d%x���JiI�桴4��/��Ɇ� �B��0s��J��j' N%3��Q�ɨ4\�u�3w^ �R�4��T>x`�1�"n���/Ox�/���#�{�1���c������������޸���������ǎa�i/�z��[��z�_������_{��O��Ӽ����"������/���>��I3ՒZ!�$Ӑ;�'s��Gf�1���(�4\���<�,{@j����|�X�pb3g"�@��а��̴Dx�z��2@��6�!�2A;K_��LE)�%SUӣ�i� B�b�V��a̖%Fn �)��#����Y-��R"ϸ�%�,�bY�NS��\8��f��"DU�����C����aD)z�`)[�W���b!!ó�;��X�l�l�N��Xf�>��*�I�,3$%0%pKJV�g��&�mY1q)4��f3&���F�� idjY\����T8�)�����e	[�h���o-���A�K������_hKS!枇���daqYgE�X���2Q�T"1&30���+M��`�!t�a%�
J˶SG�>6�樤��R&	����"���x0z^H6}��������ZV����|�9�!e�՘,1&J��jx�Y,s0]ǫ�+gs��M�b̈4ʜ�DaEEO�]�����h�u�<�{�!�H/�Fq��I�7��H�ml͢�g"����^�[���㇡���i�Oz3S9ă�;Y�� 󜢇4&g��h^χJx�MrAˊ�@xf�8�Qt���Y�.�����M^�0L5�'B�${[�1�`���"BV=*!�T�%/H����(��	L���p9#�mT��j�D�4י� ��4fː\J[�2��Jn��
S�fV���F��QFK������$^4��0y���K/��V#ZB36���,V�Xr�� >5�k�>J��i E����D,sϊ��X!S�0���%#J��"�F�$�1��	�"�[
�Z,<}D�^�\�Lf&�� QQ>,P�4�P2�ɼX	͂�pGNƩ4���9��
�� %�Fh��H,���Gr�d|d�ٰf�Sj�Ϙ�$u>��f���Oyhi�k����'����l�^9~r�2�?gJ;��#ZsV 2�j�,(AP��� ��ex)�F�������)"Bi8��
QN ���e�x�1k)%LV&��S3BJ��u�@��n@q5��}�zOS�#��_<�XHTᶀ;�Na��x�`*�B�s$	�/Y	�1�� �&%�U��B5�8Y��FF̐3���/!X��W	�U�d��u��lCZ�׍�#�r�̈���r�����A�	f�vg�}U�QfiT��,muM��R��F��߷��!%����3�[�6~��� h�����@K�㎐r��4 꼠�Hr��>&�%옸`��X���ʧ�� V� ��f<���p$x�
�J	1p��!uۥI��)�g"�ț���pH��cV��"6$O6�� ��;Sѥ$7��\�0q2qQ��xv#|i���L 3L�fK&��𫚋���Ge�̨�xG�������C��[h�o���^��گ���&��jsz|�'R�&�"��z��o��GP��+_��Y9qt��7��($�a��"��}H�q?�5��Ⱥ��˄�J��z���裏����!����Y�Y���~�hȞ�ꖣ�����۷m<8k����i.O�m*��>T&YJ�)y�f�(1J<�d������H�xph��LM0S"!�����f�x������q�m}pt���������7���߁�:��}�@!��2B5Z���ؒ)XȁP���"W; ��#���v&�i�!�6�j~���(te� %ٕ��K�֭i�,�4:��@w(L,b�W;F�Lf��TKU���5��կ�+��ˣ�L���\g�� ���������c����3�������}yf�)�8Sv�On��9�Ҿs��Ó��
���r���u�^��lM9�yv���S
T�����=r���D�B�w���L����&x�@O/�� {�����*ֳF��mGWD;UsP��0�<��j�0ؼ�뽝�ʱ@(��+��u�dH�������?�餵���*Lt�V���V_!�(X��HX�H����Z������g��=��n��\�ǳ�����S�[~á�x��s��zs���?7닶;�r�� ��76����l�/�Δ��%6_�M�Ձ���&n�x���7in������o���/���Ԭ�21;5��qh�X:
��/K0�0�vr<�>�|$9:�K��@ªլ8�t�4���K�ͬ憴aJ�:mTe~j�EǩRI�*%�r�3\�d�)	0��2�-e��*m�$G�x	$[��α?1��d;��	���K�G9���N~��Ah/.��ҹ	fg��K���:Fpն��V�f3���e(�9~-B���}N=z �8��ɹ�$���b�6T*�L�Z����]��կ ���-�w&V��J�ꕞ�p��r3Hf�	
��NX�[��(��b���w��HA�V��'���uZu4�7wF�V�_��BvXQN��O>Ѵ^�\|$êR �\ %��*��T��7�� ]L�s�+09H�k�����7ne����c�C"���ڥ�Ν;�ʚ��f��������mQ�@���1!����u 2M�I��$$C�W`��`\� ��FDǮ�S�M�^%�$A�Ϋb��W9����%�1̬��A��\\&$`��23QM� 8��!ӓG�W�s��٣�� ��ʟ���w������o��#�5����O�z۳:8����͗5�[�G�z��h}�t�_lƋ��F#��8�,)-?B�|˧��Ī�l���(͠��j}nii&c3+Ͱm����L�J@�Ũ��`FK ��*��a������	�C̋)�4��LOȗ`d*�%B3�`��Ҷ��30/�,m } ��@I�hʍL c�40�=��`X��fr�)�qr'(��1��HOh�h�O��ʲ*"}ǝ/���U&F砜g�d�	�b�NR�^ߜ4\�)!fThG�e���X��W%K�E�Th�\`pF)
MVsMXB�͟@ɤ-ɒ4s���:I�^�j�F`��lH����	}�UJ�DeI�����!8�)�,�p�⧏�\�%I�'����3a3�On	� kXV������K��!�XNK��A"�����RZ�,c�lo̸����b�=!߂���W�i�J8�i��3p�CN�4X�Js��]��� LP ���>$�ʷ`�L)hɗ!0����*�`d�fT�0$f��̝>�fIf2��ɘuq��f%���X�HK���u�d�8ӌ�-_xc��\T�̧2a.% 0�~��� ��j&AfV�H�4�d=% ��a�icp���*	Td���^���J��zcɓ�\�僁�W����״�
u�������{W��Q>Lip&#�`��0' �#U1���`�H�Ä�<0�Ac)a3�>K�;wYŦ-4�4�0dz�/e3a��ei�1��8=;(59&0�Y2��Yg��5�Fmi�xK F�%����z1D���c�,� �҈�ƒF���
)g�F�a�u�TK���FV6<�!���˖S�i�}	8�<�Z�%^,���g3���i��Y\sV�˓�p��F.7¬��[Fn�fM6+�,<�%rz3YD.���l��K��R\s��f��f�̠��s�>��1��d�!y�` K�R	��8��
�'�J}n����
ԇY��tY �rAi�(:S��S�BX�)�yA�8R_��<!�\$Cr�3S��3<$�Ai���g�Dn�$�R����6-=-�H(��ml��.�fVC��x��E�ㆉ�@�[pP�HX��˱$�d!00� `3��2�@C0�*4$Ab)�HϪ���,[0�̄��
A�&//�L> 43�a4�(y�heI����0�Ui���LÏM91�N�vG���1L)�Z�Ё`���Q�U=3�L�u�M˻&z92��;?m-.8�8͝�'XVsl͐�\ȕ\�%�� v&9+�p�e2A��]P]�T,*H�dQ`�B;(=��-%I�aU&��pn:9q��J#�籑9?��1Yfh�TQa  *?M�T)�ƈ\Ʉ43
��b����X͐3z�G��I�����s/��(s�������{A�ߡ?�	C)NU����|�ӟ�r�uI�W��c��{��خ��b�߾}ۣg�C�J{��w��->�E������<eXg�LR"��	r�:���W
�]�<x���܀�-t���<g�qw��!<6B7�=;�6�)w���u_�FrPxI��j�:����c�;g�U�h����<ۍ�N��޽�Dnxj2Z�����(��%�W��7/���n���O��s�OקǇ���=_�<<:�O,v����3�.����=�d�J ���0�$!k����d�_K،aj���hf$�ғ�p�`�TH� �d�%�N�'HV�G�;��H�q�W;x�F:� �bDg�"�A����D�1KW�������g��}���١�"u��u���r�mő�����/6�Ƚ���ߡ'������"����h��٭?�����۽�ǧ��u�����G�+B�✫����C¶��F�R��dh7�@�Uw�\��6�����C.�'�������۲��)�+:G[��6%_;�sOPV[ӓ)�������w�q�`�"E�{���$�fK9���9N�8?A�N[!BQ��y�ۜ�
Y}��_�e:�r�﵅��ۢ��f.�:ߺ�������zc���m�;���>��sG?%k�l��v�_�ӟSd������Ο�][eG���<�?�����-��
��@��%��2_��:�C?8�l����	���2��[�x:C6kN�W��@C����aiXR��{�mc�>K�����#C$�L�i�1K&0�0�p�y#w$Lh�ɐv��DF��2u�Є̱BX%@ϗ��/ɒ<�y連oK�wR@R���v��a���(`�-m9 !�+Td��q`dYڐ�,�ڒ�c3rC�/$�+4N�I����Η�q]� %��܅����"_���5�w�ȝ��44ِ��L`(��4q^Dn���{���ӊ��Sz����a�T83 *�`z�/*%P�٥FJ��HIɬ�$�
��G�3G�DCOV��J!�O�J�|5�`z����#�.�Qhx �&̐�	�
QX�w�ܑ	f^�i����3p��ȝ�Y�u���f]2`�̷��I�ƿ��*����5Y�MWZ��ĥXs���Z�e�**
��?��<X!v����L���b��!�S�J����6���+&=!*�De	F^\�Q�qfD���$�l�B��/�,�-�E4s��"m�Z�	�%CO0Ɗ�^��7�pP s�1`�<>��7G[?+�|����7�is~᯾��嗏��A���rg�_����3t}yu~v����n����
����p�r����g��*�@�J� а�%i)1�r��i�|Ȅ�Ќ������`�p]������r�	XG�FtV3���l�K�eT�#���}�2������Ԉ���l,L#�`����^JA��<ܞ�.HrU��eI�C=+Y���sC�1	Z��iK��d �������\�:�
o8A�4f��"�L�k*J�{.���+Xۏ��(��%�#=e�|���+w��U��4s��p2��pFN�L�FCh��0q�+YJL���%Y��T�e�D��KT^� s%#����g*r�81�V�L���Z�Ov�]s��J���Q�
y���b4]���+!�d�� Fyb.�9�@��j04h���*2!7 �z"4p�|!	8e"�B[���\4� C.�p�ZV.�0ӳ#�	X2-�u~�1]"��oNt��̥���ګ%Ӕ3)G"���G�AV�4d��Ņ/.%a&��ɑ�(K B���9�����%9*xK`��$���YǸ3���b3:���H�~�EIF Yڔ���J%�>	3��2��@���Rܩ��^qt,�5��gH���+sz����q�A�[�*I.La�0�y
L Jȅ�J,-�L��a'&�0N�V$S��@Y,TFق�L�ϝ��,1� �j�����OH���kJim���
��N@��X>%y=Vl����R&L��N0��F�8%�T4yhxu�.h�d<��U�B�� �,�\��.%@��	�0E5i%����ĕ�X�b�U[2���1�\���7��Z����rxK�,�$�J��ܑ؊\(X�K���%?���1K("wʢ�iNi6��6漚������l �� ��`DRnҘ!�"P�e�1J���L�M7GKY��s��u�J�OӐ�| �.��|�uP���ŕB03�\4�� C��P�Q���23����ǘ�d@v@�䢈+�z3��� �@���2}T��x 	j!ȇ�d2���_[��u��o�+ ٺ`V��=/l��s�t���{	 �`  ��9M�p�����	L��j�bPV!%@�Ѹ��ili�@^�4Qk�$�$#��aXz�F�|��E�lT�� �[tVK <1/cаV�X`�)��M^�31��<n�D���^����S@2R�9dlA.��Ē�r��1�O �iN�":K.�b���'���96zJ	X*ܲ�-��_ޜӔg��������Xsa����|�뇃^C�	�K�����v�>�8:�n��6Y� J@8���\pR2H!�	� �Fձ�VSI�L �����8��f��#`	Z�Ҷ�F�?�6�%�n+r^�d��?0�)*HKcx]�ht/��OK�N��?���>��������S��|��_K@膡L����G��p]rڶQ�乕��~����9R�L 8�r���$�\�|�A��n sȭBx�]�	��޻wO^_��(��>po�I <�{��׹K̽VA1��sP{�������;���~�m;�E����(���4	HU	�y	D"�T�g����o�FDHA뒓@���h����͝����^������x'�J㱋?��OU\4x���o;^n�=�v�r��l�WV����5� �� 0)-�4��̈<��^��5�ml)�E�v �05,�X7�Dw}W��ك1 �4E0���ݹ\:����`b���GcICB�$����f������{��7����z���ۮv5x��xM~~��(F�ŵ�_5�X팯�/�쎂��$<�����.=<8|��:>�ܽrY���RJ���#{�l�8N4�N��	��̿p����޲�=��>	pI�	/��-~�"�)?��#��a����o�;'i�c.~��9�3 '�T��Z�N*�s���YH��+䘝<���������Ug��~���g�}�\B��~������"O%�����h<�wٟ�ۜm��_�oo�_�s�^L�|W�~����zϿ���驥�XZ즵����l�{zi?���\�cl�9g���6���x��f�b��b�b��m�4y\X�g�fQ=�e G�Aq�m��<���#23/-M�d���(s�i����N&���̍;�%�Q�]�
]�L0e����j�D�Ԉ�J	�0�ebГ�4x� �g%�O`���)m<0�uL,..����c��l-����J��mx�ڙ�������c�뎹�D��4�X6�--4���Z����
W��0"ʶJ�`4��p2�m0��Y�)@v.;G�V2W��C8�R2#�3f�NdT�=n�9�R�3* i�h' 0*Vi�������d����LP�k�|D���c�4��������    IDATs���+��?�oh<�B�%"�@rh��@� h�(D�0�(q� _x&���K����h8y��UJI�6��8XB�p��a`��H����Lj�TY�:�
���p����
��U���$Iq%F�����`T�DB�w8jB;�9��+s�`C,�� �LfV%�Af0�c�_�wʁ�1$#gV<a`v f3�a�)� �6�\O�f��V#TiJL�	��ǳ�����������l��+}�dG����������
��_~2agsq����SK�3	��ۧ���Zo7�������xc��,��U��%zɠ�j%�S��p�#Խ6C$�͝�ѐ?��O��L�!g0�Y�` ��y�!�a&�H2X����8�;�^����l/�p d�r&8�.��$��qU��_e�3g��f ʙ�$�}�L-�9G^b��`����LAD3̴��Q���L�rS������!���[n0��m���s	0݁�i��%@p�w&��ȥ4&Ғ��A��7��X4�c	l��K�L	�b���7$���� ��2�r��mq9b���iE���H�,޵�1�
�ytf��0Z A@��09�l3_�%$�� '���@�//��v2��U����4,�Ś�<3�P������	���Ws�@b��(d�4�[���Rd$%�l�a-O�/�Sڥ��
xj�i�`6�M�_��)��n�3U +�Y����ϝƁN�KL�Ųl�9���l �U�ͽ�L��QxA"�!t���rO��^����3+.�r��9=/yb���\,��jK��c��H���@I�f�s��r��R�R��J�Qa��L��`��R��,1sA���Yh�ځd#/VCĢ�a S�r���,-�������=w�.��͆��:�`�Ʒ% k�,�C��	BK�pa��K0u�(���r:����Ybc��'CC2f^��i�%f�02[⏉lP��W�d&�й}2g2�`J�*K����Z�
=Sjif���̗���*.SJ0K�4�:��9��'p�)73_�	���iЋ`��٩JO0cN?�GŅ�M�/��f^>��g0���)%��-��CZ�hJ!����&$NH�kY	��H�9��Kn��4����(�&�ǔ�[�|(9bNS�%板%�eh(e�Q�%c�f�	�#-e���hX�dAk2ߒ��dH��d ��#��[b�J��$ Øi�b�:{�	&r�s4|��\V����+�B$ `6��D�-e��+=k�w�^Y��\2�>}ë�	6��K&�K3%��%4,	L�2���g��D�)ϊ
 <�&z���(�x�h0���z��oi+@&v`!��`0f�Z�� ��	G3=w�J��{u���\�i�̒1�	�W��h� l�7��@���҃1�f^�ƅ�([J`��X�a�!�S,�2Z5&{Ń�ΐy�a�*rK}ssL,�`�	���K sK3J�d����1���cKVZy�e劑ceb�X��!��Zh0��#M}�\ 3~�Jh	C�`�����MŲ��CV;YV匧T�``S`�E4s��!d	��{5��`�X!� |��	@�x��� �'��񛜬�Ұ�/��x����_m%p�79w����%�nvI�Kwh����r��z=�p����z�-����[��7h�.��͠37�-���p���{�r��B����w���g�)��'=vauXV���j�B�(}[ �Ç��tv`w�ޕ�|��}��)��R�u�W�ܪ�^w/��}<�r�6�[��.���o>qY���+�/��C�'��t�z<[[�`�1;�o܏�Ĭ��Ǹ��|]p���q���fC&r��n)�<[pY���r 4`�Ĥ!d��N�kI��f��[J%����;�U� ��f�B�.7�����6���p�퀹i�K�	����x"2���H0X^��P����%�����6��8��/�7|�c|��ס��x��g�גQ������;~�ԏ��d��:����v.�{�"�ou>���jo�7�IH����W��dkHRL�(��Q���Gv��a�`�ɞ󬑋LF˖�`���X�L�Q35�QDhߋH&���_��'˗՜�~������'N`&��=�q H�Oh���3'����*$�L���,={�I�pq8����GJ�����(��N�w����������֋'����V>W�����9Mפ������;!�}7��\n7$��B���K�N�+��q����m6��q^�GJ�;��{���9{z��un�`s���ZW����.���v ̲m��<��/��H�A��` �`J��,);Ўe��8�}�^��es��(�?�6	!$N���4�<�q�%Q�0���ׅ���h�C�*m�H ��0A�%��.!1<M��{p(
��k��o��^`Dt���lN&��!�.�2�{�A�������$��Ȇ.yh�b�<<�v�a)�EWC0��\Q��d ^N�d����^$��;^��
��������RRE��[��Xxqun�ko9H ?%wH�����zZ)(��a�{�{��w0�;�$#+� �E�[��������U)7�<Ŭ:V��O����X!E����W�js�cꊤ����{��q�<̔:��찺��������H�D�X"
��UP��t�`rd����U�#Z	��d�E��)U�t������y�@z����!��AV�����M�ڷ�dѹ�D[��K����`�\n	�	�c�RB�@JH �� FK�>�܁��r��Fz��$0��a��<R�~[Ŧ�����a�я6O�!�<Y]���;ۃ'7�s����}�����*�]���{~d��+�:������g���^�����u[�3C�ʑe�P��2$@e�3dy�a(a̖�f#��A�pt�f-4�ف�p��#�2��BR�BC��rzQ�l�>�I������&�Y��4&���-[W,��9 z^Q�[Fb����di�(����8�rD]�����af��,h��+ɒ���DA�D�Q2�c�SlY-���8r��� lF�6�F;C]&sI��3"*9����(!�)ǔc�W�9b˽���G�*��l0�Y�x� �ɚ	^9�ǖr�A	 1�"D����������@�`L�f�o�����S\��v%��(!Ȕf0sT�ДX�*�&<d.`��!��i�BXkM#GTLQ�K�,�-rْ�!��9��IFR3�1��PH�d`K�B;�B҇7#)b�� 2�P�GDɔF�L	��I�p�i b�Υ%0��{�J�X� J��4�\��,(d��1�RS�mz2���-!�đP��R�B�7;pL�df��cX�יh�s�����L/JH�2ǘ�h�0f䔹O�#�D���%�Hw��Z	j�!s1�pZ&��g[Eܐ�]�q"�×I��E�i��0�,���0Q"1p��� c6 Vr��ʅ&<N�B��.+�0�d̄|��1Gf"{�����(x�R+h �I� �>J�7����?a6+*��͢�E�@C$� #<*C\�jp�Lj� �4�X8����;_J��ЎH�/�4LFA�s;�̑��K,^K.�=-��fVH�dB�0����}+��։\�8y���|��SZÓ�ڒc..L�P��[n�0��Z�,kTV��T�`�d���' =�2�K �j	YE% �B�FʂNG��c����J`��+�%���謔�X����(D�2�m	��)��$��iE�Gii�`��6R���P��8̅�͆.��DO�C�|H�%��0Q 'CI���1�2��i��90�l�#SN��0��ϊx��a�+B#~ xK�e���)O�% o���J�~�2Z`����M�dC�(�R"/"B���a,9�p!����`�z��1
�*IrTh
D���@��	Y$���L ?/��3����� �T�@#s.FQP�G���V�0#�%�z�L�J8=Q� ��L�զLJU��� �h)E' �f�(a�%SBJ0gk�-�hK`�����/�%��)NzJ!��R �W(Vzs.f&��� -��d�8��h0G^\�&tP�)+$*�Rxz$L�a�f�uÒ;kgA����@RV�?���	
$ �.,�X��fq˼Ta�˗��al{Km�ɔ;1/9���{�u�8Ρ��\�e���l�c��
g ���9���{�c���qW�������O}n�� ��z1ޥ��ȓ��dl�����
�%�!�V�}+�P;���p��;�n	Z��`��m��z(���HZ�P��Abx �٤����|��*����݉�սY�j������(o������e��<����`V��aV
 ��Ex�𡪗ۥ7��ӟ�Tg�y��0y�W!bi&B^n2�U�{���1���ǟ��g��G/������w�����|r�i��֗�G��6�o����w:�P�Hc9�϶+%~ѕ�$+�J`��P�AOi��-=�~��%�w�h�������5-w��C䚠����Y:T��7�w�������.�co.c�0
9�[6�#Z6V�
 �4KF��V	��j_�.�ї�����-gؾM�Y^&bǃLO2�]s�W�}�	��k����G�����������K���s�9[~>���l�5Hin���Bb�������I�;!U�H8��)5H����0z���`E�w^6���,�?��?���yK��L�$�ّ����?�s'��~�3[���ޓ�c���
�=��ۿ�[Jǉ��k�:X�B�!?w�^_�JFn<��N���N̪FE��߾}��G���%m�$�+�'qO�<����=������w�կ�y���W^���ۃW�ǎ��r�F���b;��x����5͋�*0��r�$��l��q��ӀqZ�=bB�g��?l�UŃ����qG �'>�ڨ�j$�sZL����.2dm'$s�,/EcI�L`������f|G��[q��� �]U	\R:!ɲr6��%/�b9p�aǫ��@[.�m ��~�1`�8�'��@߀�(H��*�l���g%`�!3w ɸn�<x�@�����';م��4��F�.N��=�T��f��[.8��Y �$�K6�F�OC3QIҖ� +�~�t��������ё �A���Lw�����7 �r� O������;�d�3 ��޽K����^3rzq��4�tL�
s��<���
C�Y�Ҹw�$)�X�.yI��	f�C�V@, ���i16���~�C��0Z��]ʄ';���#%�j�/��U�WkG�pHt�%�:&C,�8�'Y��p��_���x� �n{�p'�=��î��h�YD��_�򗶨�+DJ�c�6�TR�7a$��Γ	�`f��DD�d�S��DWB<L�G��U���\� ��#J��[zKV2r�R��?w��i 
Q9f��1g���[���C>X{�u��l\-�z�~�k�c�|s��5'������ýs�ɿ����ٮ-W�Y�"���xԺ�(�yX�����U��63Sb�	��`d��6HC�hX�
��8/��u�  �sKs���`#H,k�y�C�X-�%O����1b�ҜoU�ˡ4h�hr/=�F�0�R�)ӗ3Z c	2N�|����(yɁ,(kJB��	��@bf*9NK̅�1�P��"�X����d�r���:�F�b������>�|��J�,$����ff*�(��f���9���i�+�J���X�cK�PHX	��H���`Η���+dy�^13��iĢ���XH3Z� 3�0ds���)��i�K�@_�� 6��r}I3b/C�\f�UG�,�9�p�酆�{�R�ixu�d1q�7+��15��JI�Ž3X܎8�Q�	3�\�R�#�c��3ӎ�4��*0|l��L"�E�������2X�LUM�֠��k.�g-�\&C�%��U������p7�/$��y9��d��MH(Cs�2�%zC�U,K��J[R9$pdf�
cY��&P�cQ����AE�\�0�L4J��4$L����K@JF^9Z��3�������>9G�eDޞ�b�$�	9��Y*�Cn�hxI�<�)�����M]�l�.��$��|ȲU��-o�1�VL��'x��������(i ȑ�~6�9�l��U�ɑGK�ΡDU��@	�T#��#%�19��`����L�ٽ$��$�d`��^��6>�%GrV.�B���l͖���g]3+)-�S��V��R!B� ������/!6����L=*�f'&_&0`��̅� \A�e2�p��%�^�t�K!����,�� �-����F8<�`(�l�����%_V��㡯�\�4\�%$S\�᳚�s��=W�+�O��ee��(&�2��6S&[�h$��|#�c��Д_¬=��0��!�eT�GC/�����ޘ 2�e0s�vB9�ғr #�����e���&"���d��Il0�C O0C���0��U&L���>6T)�7s�'�@��d�4��S��[�K	���QP�
a��s<�ބdB���I 0�M	�C`5pr6�1Ј�ތ���#Y���h�� ��a�=O!NsTd���"Iʤ@Ƚ���]J	40��{z_9@"O�D(1Z�
�Kظ(L& n���%�p�AH!/�,��@!�2���ph,��jT�#���!7�dJHBQ���Rڑ��c(
����i�@K.ӱ�*dvO�0��o�#D�dYnf2ZJY�g�`�&�iȔ���8�TTM�+d�#�h��$=dK6$�2��T�%F�^,V<�&\��KS ��"�S�������ge˭|[͡<.���o��<_�a����y�į�9�����,�ɽpxf�L7��kϰ���XܹsG!0�)��%�M�R�w����g�F������s�L���C����pw���\>(���G1�s'���_��g+LЏ?��Q����[�e�	���G�j��G([�Qr}x����=r����O��@�,=��%����'g�{�٣��ΎOV�|�eao�2���'�7��9��*�5�����q�,J��*��!��L�/3̄�a�v,�$P826Á�"�q4��'���a�FK-	4���#fq|�U��b�ѕ��*��Ϋу岎�J,IX�#$��,�7W'�{������O.{�������&�_��ӋK?g:���mY>���y��z�n��3���or�;�8�����ۥ/�~��Ƒ����7~E�/���l.�u��6���<���Bu��<�:���|���霤�<@v6��y��|���c��4}�Oo�/	�ϣ~M�0�_����������I����7��C�܏p�:�q���x��7����q�X�X��i0�q'���-���&���?L�Q~�d0AzN�{�{�ͻ��v��W6�ӛ��y��o}�[��������"�\�k�v�/]���\n�|���w/q�����0���������v����l��x�=_��~��x�3��Y]����_�o5�k��-U:b-/�fʎ���?jYNQ-%�Br�v;��������?����U�%�����BXR�rP����E,�ꄦ�!c��aCR
��De ��p����m��	�l<z��N^<�sW &`KţdJ�0�����b��Nb�^(���y!��#NA%�̢�<�	�#=��]y����V���{�GV��Y,{�\Jha�$��F�A"(~�R&�GÝICd����<�,�!"� ���#��B lJ�cx��!��Sb�d��@@��"8�\0x l�g>��.�L�%&U�|��W?��H���
�!�@��狟 =䅙,Yq�b�ƵB2ȑ`�<ZV-��)��$H���`f�4#�q�]V��^�e�4�x�v��J�<�
)O/��
/IƱ.I��FԜR�Ì��9s�DV��gg��'?y����7QP��
��%�}C�$f����    IDAT0ӰN�%*�F0e��M� ��`�ђ��(K��:P�q�)�/��0�,è(Y&Q̆���d�<{����`��P�A�|Z�qY�����Y�����͙G���2�h٘ǿF�٬��]O7�GPh�Z]d.�����f�K���h���^�dJr� ��p$�<�7!sI�����&G�h���k$�w� d��d�����m�lN�Y��Y���3O�=wJ�8���i !�J��lP��2��|"i��;�W���CO6X���`5
D��wQG�J���f�|y�V29��Tq� ������\\�:CS�X�s���-7���`��Ji�`#���/7�QP ^�gb�i�L8�ц�3G<�X`h��0�N%p$�+���H��m)"��)B��i=�	��C6y*�r&��!
62��"q�����V��
�KYh���R��Ec�I/a!4TҀ	\tr!�2Y�1�#1Kɒ�A�l�%l�.��
���g.�b�0	�/J��R���Պ���$�8�ES����Wf��A�JcI6�`�4"��,�|�`���:d�`f����8��� ���	��rC��Q>�`��p�4`$l�TQ����-aBH�eT�`eR����K���*���-� ��,���󂜉��2$���7�cK �򱄑�X�hX����ǋ̫X�b�1�掓ol�gJ�</�#B&�S×�-9}��co��޲ZB6,�k�Ʉ�)N�%φ�ONrQ��!��fPFh��O	C@;C��g-P<�4`޴$�KC���-�4h���IhG!S��uq6�'Г[��'L3=NT����s�!����ޟ���+}�xJ�R�d������R-�@6���0��D��V�`F	��d&�v�Y Ch�8,�{􆟻��0���� X�kfEKI��b�4b�'��l�!3�% 1�ާ��J��D6X�Dڥ�DI�A^��e�y��"��` ��6��Р7(�N��	�-�қ����� f�Ӝ���: 93'�K�2��̖��pi���+�	Mʼ$&�Fl4�.a��3
8/Jp�! /d��d�6�ds�g+���1��!���1�,bH�NC.��H*�Ln���1��#/�����0}��Qr�a�pr2�9HzB����J�F�j,1V�L%�T��$��d5�XNd�f�]�d��`�2D�f�!�-�eB@H�ӘMc�W���R�NFld.f���� �4�#D�˒56�lNɊ�/yzK�����;��d�,�#�����ZB��(a��(g�4���KiI�6��
�L�ƒ�� P��DG����ǀ��*���o3����Ni��'`#@�N�1!G��B`�<̈́ɪ>㡌9dyRQ�QW�:C�,J�d&!���]�	 ����ŪR���z����/�cm����)J���ђ^D�-�c�`���d�CS���WB�,&���^�q��=�����Z��h/6���N��{7^�ϒ�����n���oW}���_:=>:�=~E�~�ytbv?��E7�F�����峻�{΂At�ap����n6J��O7K<x�Q�����[�"rD"����� �-�~�#�J	�!+�	�댛�fw,-)ݟD☊��oۃF�cq
�K���;%#!���A���}�Y�n+\D���3���p�����xg�_��.��e���э�|��o�������r=~�t����S����	�W��+��f�hGDW>h�U��ZA`u�CZ�p1�#|�4�B��5�1��D!�s��I5je�©�����w�Ա^��?������;�:荣�*��q�(!��쒮D�Ĳm�Fs�,����n��`��Ҹd���釕�� ��v�z��{G���Wg]ɐ���fz`��˟h�z��h׷}�p{�޵�w���q��q�/�\�mw7���[���� �I�P��@	a�*��1��<�e�k�]�?�Q-�1��N!;ɒ�^4�"�����|��0�7i�!f��gڣ=u����Ou�	�^�7#�(%����1���rv�E�BIf�?�9 m�d��E�	,I&���ۺw޽{����oy��p��b}��_:_��݌ù�^�C;.͚6~v��6���]]��ƃfO6ɞL_��ꮫ�7C�����|�����������?��|}z��	�͹�*z�nL���[���e�.�$�_���G��������w]�D�Ë��l	'���<A�=$r�@p��DI��)R$�>��w�2PZ�U��_ժ���ݎc�.`U�H!��iH���1 0³�.0�4 $�2�pvʤ���A��W���>� �QTv�2�F
J�D[0򖋗B���L,$qi���q�#W�H���OF�K12�"���"�li��eq��	�Ğ셤j�w*t*Q�xY����E¥ٳ@xg���y��rVz���"P.g��kKK�#��٭xmT�@\,N:������0*L`��Nw�Ts�����R<]t�0��Q15����3���Nj�*@�ѝ�IM�awҍJ�j�����4$�/���{�=5<*W�WAe߿��b�]�( 	�\R`� <Eg�C*�u�tlu+r�j)<����.n�(5N<�rqy�/����US�Y$�
*
�E],�F.�^��*�Օ��!0���%�\�B��N` ;��(@,;<p� l�@	�a$�],���@��"K0�Qi)#B�Y,0rFF��2沜81�+��,��Jx�
�:c�T!�ۻ�L��\�$:��I�͵/�W���B��p�R9~b�͡1U����^)�j*�l#�%{U!a,����9�YC�(�B�Had�v0��b�jbL;
ZWUa#��`0:v\t<��G�n��B�[�zL�r4�b�P�(enr��&��˒)����4L�6�뢗�	XF�#Kl�fF�Q��6kE�Y�=�S8c0�bY�"��%э�m�'�fAn
�e���"�$c�q��� ��>�\zE���V�"��c`!,�P�^%\������1�x��,�r ���t"���:{�2�)/~��YҜU0�X:�P��)�F�ú��F�B`����22��Z%ͨj��	(j0�"��t�l*0���s��|I�,I�9ĕԺf.��mN�bd4�T�im��T�a�	/;��	a_B���H�FH/P�
+J��3��`&�H�:2N .:����e����8���4�Xz�,�盼V�����1d<�)WS��H��qR���"W��ّeG[����2ҥ�f���h�Z�YHQ��QUsQt+b4����N"d�30�2Vd� �g4�^2B}�-�����"ѫ�m��9�)vxṄ3�3+'#/K�`5ir��`!�*�,>���U�Ѵ%PL�K���d$���K��N^=d� ]Ǘ-¢0���`��)F�2"�m�1�Q+ ��r�E���!q@��`F�3���,{lU��b�W��{��_��5jZ�aA E�0���?%��65�Xv����5V	�W�qv�[Z!�pvHvQhM��B���}�� 1Ћ��������Q���1�u�w�񰛦�T
x#�J4�5Y�XJĒה����O)��^�V'��2�\� ����eE��q2
��B8a!+�CQ�u�1L��3���[ e2�K�H)V�(;��� ]:J.T��[Ne 	PH��������]�I`#*.Fg���
7�e�͔ȅ3�iI�a.Uub�����$]�
i�F�j ��00�U��H�^lcI��!DU^_DA�W��%�Rv�,n#�{X���{�[�Y^T@GV,�*Q)�)�$م0�-�i`&,Z#����*BVm��Oi�VZI���,�FIYji$V�h�yK��_�-��T%su-?*ޖ@�"�\%�pڥ`�0ŉ�e�!HvT���X v�P XdDB!v���r��%�e0*�iQ,�e�()B�- ���QIxHx��W�_!��쳪��X=
pXが_%0�a�������a�k&W$,�<�e�//%�& ������ݦ��qTF0F�,�Tjc5�b,�}�J��޸ {����==9������O�Wv����O�z���ut��	�9�T'��>p��sJ7-��p�������+ϳ�۷o��ꎱ;��y��6n�������۳:���><������N�H�jv�ڽ�K!������M
<�����=*w��<OA�����x�z�t�螹��������m�1��T����逺�+������[~�px}Ü�J��:�x��{���~Pݶ"����(ɥ������歿�����o�q�K�O���Ӄ���Ke�ؘv���9�4�X��с�f�k��÷�����z�f9�ō��b�`
/#�]X�J�k�G,�`�;F�������-;��@����X�����)����@`%�f���̫���~�t���d\^]�����nɻ�����y��v����G_�\Z���{�M���OU���~���kW��^�Wk��ٽ�u������v���J/�Xy��)�R��l�Z�g�}��Z��ڔEX�ۈ�Ɏ�n�=�Y��Ee�礕�ۻ�,��ľ��;�FU��E.���ˇ~�|pb��6�:}�SR��Ht網����|vrΕ:C��4É�����TI�vZab���81�?x9~������g��_��8��ھt������/�6^��zyz2�ND�?z����S�q-s����r���Л���#k_�=��P��K��$�~�����_>�:��O>G�	v~��r�o�#��Ų��q4e�R��T�t B!Eq����g�'�b3���Y�2�$\x���76Q	���q*CH�`��8�v�,����ݤ�M��"�5����);�#�p�,VT=G"5�X.0��@������ń��z����6������irٓ5�+Y[L���E���9����w�����֭[N���9\�F�BQ�����M�b�D1�j�s ��Y	�a��t�2���5x94�:�aP���B���:vM3rY�Z�@y�,Z�p<�Jg�"M��'"��i&�k�ނ��{]�Q^�:��m�FUY��:|����*�qs�S�,b�j�����=��H^�c7b�&��Hai�2y�޽k*Jm�U���D�tR���X`�D�<FH"DU`M�ȨvI����� E�H�X@a��Lt �.]�ً女�=Sz!rY��S���+x.*/*c��+��
�R�0��(Ƽ�!��=��-�O+��ؖ�G�i`�h��x�v���SK��խ��f�)��[#�qi�-���4Dͤr��E"R�H*�v��
0�z^#L�ƺ�?�L~:��������_ �i{�KT��4�0��}$X0�H
F!�j.uI-*W�b�˾�z��[Ub����di�8�M�*�B�^1��(�YU�EW!,��0�ㄑ�HL��]�Ѯ��^�h+&B��7��Sj��~�,�ZQ���,B\�d����0�tvQ1`�-�, F+�q�A�O �P�Έ��F,�[�J�& ��\���s9�2��-
Xo3Jj����?V��ୁ�3�x:Z� 2!��HT;p�H T���FQ����N#��ſ���ÔB8��.1�&;��B��IGҔ�k��@�y�I�,�i%S*�	�k2�Έ�7�,������0/"Ec�1��f�F�>��]x�y��T�tt�*�����a�	cQtƄqq�_9��0
,�N2�B 6�X�V@��,��3N�z"*K�� Q'i�)��5Sv�p#@Hb��-c^}���c	@`=G�U��i��_^ǅ"�T��,2:�A�FQ �xMIǔ�̢Ɍ��(T��I!Ĳ��Hmd4��R8|�4��)���X�Ŋ�SRsM;��=�0H�Zc�g$�0���]8g�yc���"a$�D�Ѵ����l/��"�l���[Mx��a_(G�R
�+�[Rv��RS
�^�zFi:a��f/Wb�@Q��F�����*�&$���a�hK.J+*6��ʱ�	|V@���[�"Ll�j�` c�S���b����3�@<���
[^T,�����'Ȯf����y�߀�~)�8�K'zKWf��A��'E0:ᥳ�i�3f@E�b��m�М_�E�H1����^�E'%Bc:{�FQ��̂PvSಔB�+���K��F�z�)�
��٨� �S��J@/��\��A�Lw� �q��%K%�rѳ��+�.��(#�!�״���%Q�by���5`�R.r�S�U�v��c,c�pBg��ؙB�T^QtyG�W��c�=�k#W+� ϣ`^v��XSF 5�Br���J���1BHx��<�20j�6�D���~X��\�)��Ơ6}�); W��� ��T|T��
��C����/9ZB����.Q}k������D�3\�~��#�P0��bຈ�-���(�I^�x�_.��i��&�)�FK%����U��5-0`�2fs
7�GX�1O�\0�¥��2�P���V��˒= ��_HT��(����Kg�.Z��[�x(1�J�LRJ��M�yV�Q�P� y����� #�@���B ),�L�a4�!�4EU�MQ���~��5~��lD�]^��a/_<���ӗ�[g�O�/<>�x���on^�u��}O:��b�"�����[�c��3�^+����h����Y�)�[�j�#�XF:�`���4���4čǺ�E��3��Y�;w���	GN�ь����j��r��l��?F�:���S���B�d��s����J.&��ݍ_�`���|������{�Q�	��{��R��/�m�囯VWNn_�Ɠ���9�}p�d���3�m����ϯ
�X�!�X�Qٌ�@=,���`!,�D�3 $�e
�FS��bՎc�4 �O�g��Z���E�=�6>J%�@'��q��w�R�Ƒsy#>��>���v0�u�E-�5�qv��g=�<9���ӯ.7ㇵzJi���x�����Ħ.�N�\��N|���͕������`�����K_�v��W���y��w�	�?�Co��[�#�Ã��/�R<�W�R���&0.e�.�s}R����)���x�b�
�F�5-OG?X������ ���mM�N�O>�D��o�V�S�(!���o��i��� �ˣP�`=p"�D����J�,6�L��'�*�U�d�=1==>���c�_?����X^��������ަ�B=?z������>q�>?���w�p��u2���N��S�	������ۛ��V�f'�j�l{���ͳ+��g/��WmW]�]Eꛩ��\F�t5����0v���1���z7`*�0FXgX��*��1�+L.BAC�?7	*b*P��������X�\��Q޹(�Q7(I.��1S�E�3�iDX^^�p �3�檒0N �z�^�Yڷw��U�Ç]�[/ Z�ەJ���x��y�JUF��іs.F�6��y�n�۞}�A:5T�(x�P
��>/ ��MNx)Z#aqv;�p�e�N1+B%��Q	���t]���H\�j��(HO�fu*��M���+�(ͷ"�)h�.��8	�p<Y��-�E��8�$ e�B\"�.�y�!�n��o���f��*�h4q��W p�LT.�S����Ű;�`���b�s�j�Z
���`.��K�
зzn�E`؈p]^��U�:�e�&��� �M��f$����)L`�Du����B'3���Xv:���!�ƨ<��1��ҁفM�)@#;���n���2�3��(D���ZǕ�����rS.v#�1����q/�^FK���_�B�'�)�C2j���xm�0�(��!�P�1��2R竫4@.ᲃ�7�¨���Y��t�H.:pl��Ug��U�zfSIFH.$$0A��ݴ�S������%��ށ�4s���8������xf� �#O�L;���52����0RTFY`:b��V�LW�pJI�Y�.zF>��    IDATK�8^��!r��) ��1N���Ll����.�H����45�h���[)�	{���S&�b(�x	=ڢ0�r��S�T`�um;�"���x��e<B  ��AX+���°O0|�k8@.���EIQ` 'g��(��MPT�\��-$�,�R�3R���E�nS��@S`�\5/ad�z�S���o
 �b�9���eQ��f�����׸N����r d`1��J�³T�
�R� ei���"\��a�J�(�0��b4��]x�u~.�T$���c� g� 䍖%L� M!y)F����X�2�1�n,�,��x1Ԩ!g^���FE�~�S��S����G��E*:o��4@�Q],RIHZ<�,ȍ��$`�r�%l��	o# rk�^ �R�^d�C��ꡔB,@!vT�l��{��r���Ar
6#�@Q�`FSbJ�'@�Q����C�!�Q�
%m	 \�!J�Q�3���.�Vm��𢅟�(��e,�)i��!�]�޺��AU�H
�./e�zQ�)��sI���Xtt`L1t|y�/W�k�!�'�5J, ��B��S:T�\�0�K�ڹ��M��9F`z��ӄ��R[�4�eX���G
)�  ����H��MZb��1�	Q�M�ѩ�t�H)��萒�n%D�������>�u��8��|�s�������^r�eARq����棐�C�M%�!c^R�䷥X��I�'iy��{Hn�1��v�U'�dTݳ������6�+���E45[��rɄ|�A�G"�Vt�/��nG��w��cEY��l�):0��[��6���̫��4Œ�tV��4�J-�^�Ύ��>�8-p���ڜvj����	��� �~3 �����j:�����[KK$eY�D�`���Q}�����z݁�i�P�8w+a��M�����ak5�ˇj}W� >:5P.\!�i����i!**h���Ճ�>7�269&��i\sی��8��gH�0��l*%��Xc�X���-蚟��L��V�
�����X��l\ui�N���lb9�धĈ�&p�\wA8"xa�j#�U��!��74�M��Y{[p�������2�(X�6U%�/��FF�ݡdRԙh�����BnxY�Q�� �����cHh�s�o���Q��)A�w:��)�0���Q�|�[�C��ړ�z�kA2�%	���m�(E�D���A�\J[P���Z�bO|�g���km�{�<Y3��\�����YД��x�`��ZUk�Ә;���P/T7���ġ�6�x�<RA<�sp�+ul}6�Ϳ?_�����r�����7͖'���v����,��S��>�c-]�yީP�(H�/p������+��Hs)E�nBB��a�N���Psv�aǟ��݊�w۪�9�I$<y���z�k�/�f������N�̊E~}���כaߞ�H����Ϝ8��/ff�m���t�؛�W^77A��+y��K�՞���,�׻��Gg	I|� �h�N��a^����b�,L3,Fp����k���<��V����V��H�f��',ʰX 
����w�����4fOf{���m��i�yp�����a	K��;C�o����d��oQ~3�G����tt��zն=�X���Q�j����7���<�<e���PM�l��_���^�����G?��W/�کi��}���̲����hS���\�"�z[[���B�i5Ym���)��e�C��n|5���D���鏑��%�>�{���������G.*t����0��dL�L�F/vK�qy�l���NX�C��Ÿ�n�07Q��K5���
aw�1
?�/v�d���o�f?�{0V![�'w�z�������.��ٲ�B���>~���������)Z�?H̼�Jp(�lѵ�����a��n�Mu����a+_�>�
hhi��XY����]E����G]�F)���D�T�߆���K�E��*����mՊT]u�U��/�����ir8��鹎����p�\�D����V^����&h����Œ�|u���Wk�ƪ�+}�x^�)_�C�����x�ڂX�J"�ITM�䚚�R�_���IG*�1��${�a͒���k�A���M(&�t�9�l���.w%$N03�~��4e�G����^����P��vL�����ن`��ΰ��]�{����t�K����	"���2���}\��~>���#��5���=���фɸS�/��i4�|^+�*�j��f��f�\�?`Ψ��v'O_���~�5��5+�~��&D�Dp%W�^�oܓ;��^�1�F������:���i
�n:���D��Ym ���k�
�!��k��)�����7���*o�هe2T���F|��� �֪�{�Vޒx���f!^�~�x!��������ZS���] ��b��]�~1�"�?���=x�o���E{X���!�a����y�hZ�B���beX�0eX=Ӧ���]D	���N!Gp����~̊em�a�^p�m����Y��Ŭ.k��^첓�jg%P�\)U��K�5*&޲(S�p�2d	����;fYo3�z��Y(Lh���6���k���t�2�Bdو0\��'�W��6�	��}�DQ��B�U�b�2��n
�`���
	7�_��!.h�s�R�O:^i#Т�B�Fl�)�����h5����o&�sWB�'�@���%��g�4�R�C�2�S��������.U�˙\wŤ�'h=7b~d�TA⮾5��	���0�FYb�1�Xw������p3�6Y��>L^�ʟ��$"\�~��EF�����@� ��еG8��D��mz�`��a"n��f��R=-2�oVz�Zs�$Is\�9��ƍrxN4���CX
�����e$�ã�^:_AD�2%�Q��F���3�K{x�0n�{'�a|��$�f��)z�jV���.�2�-�3byH!&��]F�l�R�&U~����K�O�R�2!� �'��������7ܜ��j!A1o�
bh�,x����i,
�P"����敮��8��%"�Vc,9D��7:��ߋ_�\E<�p��kؔ�S��r�jħ�S��獍�u���}~���$�wU�)y�\�{�	k%�@�"6�<ޙ4��<{5��D����2�������ϒ�:n}��B������m�̭Ѻ�)bi�E~�!��)`��x縗	�ƙdS"�F�4)����J�:Y������}��(ک2I4��x�^ͷ��@S�p�|zm��Z���BB�,X)6���AB��a'�a����Zޣ��5B�*f�����a�� }Q(�@AiK�26��8SW5�X �&�Ӗ�=�u��$bE�6��˦5W�1ܵ������@�D;�l�[��� ���87#�����H�f�(��樞�U4��z)��L$/�{\�f6�����y�#_Y�O�]XVb�V�H�(�L!x���dU{y&���U�B/2��gA �!�C�%�(���RU ��Z�h�'X�O��t�HS����:��+�kJ[\���е���C�����,&,�R�v/���;ni������5!�� ���C�!���1oʄ�<��H�l2���w�w-JN��H�ԗb-�Pne%��'��}�c'ŧ�(T�v/�	�llHN��&L�Y���5��ϧ�h�[��8I���e����e�/3H7W��]���{{����uj��������SS�e+NF_M�
3dP����? �>�R���樧ֽp�� l��o�?�HȋO�d����ϓc�o~����|�9�\{���R#��W�8�n�	:3Y
�'��kNw��H�}����y�D��{݁BAsh7���������#&A/�����9����!�)�N=��:��&�ҍ��~6Oi���)ٛN����zx�V~5���������,�0��r�Ǯ� �z"�9��:�������ּ�#�W�e߽�/}|�'Q�����ႊl��������w:n�D��?�|{�Zq{�r���-��ؠ�ɻo����/��YŢ��g�����+�ð
�{}�����)i@�x����ǝs|T�n�-�8�/H)*��g+��O����d���.���oÖj�N[�s��ڕ����8Z����Bii,?�?~zҧ5��s��6��x����_;�K�T�)}e�
���o/���?��x�sS�H��GC��Q5�$K�0u�y�c���C��e�&�o:}��ƿ�Ew���CJw8(�������M��+�,�N^�ky�+��7PH�L�Ytd�:�<��P�����N�Kxq�(���rt����͎����-�?=�Z{���S�j�ZRk^�����Z�l3������Qw�����{������A��{���|b���`I[�cgw�ïv7o2uw|A�IՋ�8�5�����6z'T�'$Ih
��Lew��x�P�5�lD�Q���ԩȲ�Y׃/�����=Vn���=����QI̊;�l"�Ꙙ��&�w���u�"��7���4���,{����R�R�G%���qk�Ɉ�piX1��C��C@7H��q4!�h_�6��Z�[�i�-c��_��faD�;WX=�	���D�\G���=ż!���h+�֢�p�^�1�x�&�u���R2W�Ā�����[P&���f�g��̌ZxNS�6�𴪻�s����� ���Ղ�%����;��ʻ�ٓa�{�i��pYd�0�T�Dr��[l��n"T�b��q�M6[���2���At��/�&
��6��:d^�i����	�����J~�w�b��|4w�o4��H9����h�m�$5�U�:}�Tk��N1�ض˲FH���`� ��
���H�����Q�ʢN��8`�^?4�) �*�e�4Q��mz�}Q�����	���#�4ںf���	S���99#���(H��o�����/]��a�q�44Uע����P�%�ZI<��{&J���ϸ�7:�/{GΨ�7ј4���n��=G�O�24�I)�N�u���$\��k���@Mx���P¡ �j\k�iovK�?Rj��s�ȣ������
;D�w(#U��h�&������h��	k�k�[J�g�[H����{/��jЙ�6�( ��o�'Ŝ�Z���'lc�(�,�ċ籗�]VR������R^�)8e��$1�\�k��L�Qߜ	�4|�̛��1�ɡ�MTx�����`Om$yJ`O��l9�_�8d��<-��P<?�m���y�Sg$x��j�ª�~׮A��L�#���<��X�hM��A�pl����մ�c�ŴPے98���g�,!@4D	'���hV�X�^etf(��ɤ����MWDq��Y�>H�y����iͭy\�'�ާ�A�g��{�Z�P���$���U�椢�\v�)�,�i
��1�7X뛇{��~�!���D��/-�H-�M@�yJ�x�[�_��4�@��Qf�6���iI&��-<iI�0bc�wv�驟�s�7���.U�xHd�=`P�S��]��W��"������� ��t�1��09���<F>�6���+�)g�����5#�lS{$�Qؠ#��R]�GY9b�c!�W�g����˂�C�i1�]���d�8M�b~���KF����I����W3t�G}l�vu��x�(�} �/�7���Rʌ�����f��\mHH(���4�%��N"!��b�~8����;�v��p6G����{«� WQ|������L2�`b��Kս�0%��+~���o@&c'i�(3�1V��W>U$?k�to�����v�o�!�Q��H����c�2���U��3Tט�I�O�]�p�	�@������r_3���V����b+%�4o��OHh<�T<�K�0����C���Ѵu6�HV��n�%���%z�g/(�l*���h��%��h
^ʚW�;�8�%N`^U�&�o�fV�O��?q�b�tˡ�A���	L�ޢI͵��1���=��}�9Ph���UI!�U�pQ�tD�[��n��֚��V�
 w.0�@��,�^���z�2(���w�CD���d��(�����>�6�D���FO�u�� �-��-aT�� ��l����aV������B4*u8I����q�x�7� ������Jv+��;���E����4Hr���,����9M)��׋v9&6b�~�6$zAn@��bퟯ歹�;2��P�L�b�b�񛒎`�,�b2�kz[�L�����v�y���ۢ{����S��uQ�W���~6��??�R���ȹ������.��ϛ�?��}�{���]W�o_f���v�M����T��[�FD�ɇ�/�����t������<��W�w�$�i���G�n��:�T�Rc��Y<7%�ݕ��ȹm'�d&������o�+�Zt���U�}9Tl۔�j�QX����J�����0e)�� �G�c��J�r� I��R������Kv���c���1��['KS��W�mV��������*���������.¯g��M�S������6��?��M&$ILTAW�S�
��V���5�E}��^ �A�����6n�m��%���\:��5(y�{��|ח���Wu�YF :�G�2D.�)�`Ҕ��E`��z��"����ؓ�7�y�m�c�
�����J��k��V�vZg�]<\���L�]n�k�|~h�7��6�rmm��QWbp����'xk[�����v�:��g��տ�wZ{�W��<�9�#p���������I��}��K,>���:�;���jzX��#����2��[���_�Z��K����)f�Slb�eN�:�G���~��=�)F�ј�s��R��n��K7��;�{���}%w5����ZF�����wOK5"���ww?v����r��1��k�Pם	���;����_?�^*��{ytA?�7��!����.�H���g�F�� ��$�����ɜ��Y^�����V~O����?�>��}��|=xe>�H0��{Az�Z�#x���o�'���Sh>k�6t%��l�����:��T��M�:&4�P���vxqi<��"Y��v/��2R)��Y�D�E]�f��λ�٣�r}�ߍZ��kth����B�J�,�3.���6r�Ml��m�]DY*���3���w�v���o%5K��b���]�K7�Ar�������v��	/C5p0n���PHt�D�w?풯m	�i���M��͞��֑��f@��[����])8�sD#^��I��l)I0��N�_?4~,�% �4%!�|kn;;���ψ�ܰ% �'E�܂�2�y�O�{�I�P���ߓ������mɷp#���?��LZi���W�:�@��8@�����2�"J5�Q���@�gj��:�4O5���o��9<An�LB�̲Ѯ*e9�,�]�]|���4�`���[����p�74�Qd��I�*��wt����f�������L�R����k�#F�`xi�یK�2���P9","�/�^kRF�@6k�����W?Ήv��0�@��Y���v��*�Euh9���ʡܔP&�7y�I����yd�c�Ww娠 ;���C�4�+#�8}�g� ��!w�����H���w�9�Je��,� �ynz�R� �h>tHn�w��{Y�O��ROM��)ho1���Ƥl�R��Qe���E�[�
M��b΄=k?�ó�f��0F]��{��(�BN����e�I�B�!�Y}ԍg�l�Z^����H�����]S1���@v^�_N�W�M	�;38���Wx�U[�����(E���@�#��!f��,6���^��X��Mya��8EiN1�t�������lX�A�6_؞t����\���7ɮӷM��di���^9l-Mm�3�`Ѩc��!Ω RMO�,Uȋ,:��$i}�t躀�z�@s{��tM])����#y� u��}��Y%���_����Jj8u��aY��hOѳ�/	�����d=&Ժ�F*	���
��F��,�����녁&�-M/�Ɉ���Ūt�]�i�� �������Aj��c3���oixtSۃl�<?%^�be�@ZF�{�7Ÿ��7�b�/6,��mY���fV��y��I=��>��2@ e!�op������������oj;�7��Ҋ�A2x�$L��[����8�]K�'NY���z��9n��L�-�!�s�[2+�l�Jw�b�EfL#;���Rm a��|�z<���i��u���*��P��g��Ae�[S�Y2e�m���f�<%�H����CjM�'�pE���&����H�i�QQ�M`�L�(	�V���7�	�"��>�h�F�����I�oi�@�I)Q�6õ�XTU��T��oZ��n0�IC�x�3dD����B�����f'ȡ:�e,���j�Q�G�	ݐ�k��m&�-��n,�Dwoc(��X�	�>�Ik�G�J��Q�Y|������Vܲ�#a�{!Jꢒ��z��A�Ne�c���?�5��A�+e�/�d%$���ٍV�����{�ܮfzXN�M�a�V��hwV����X3�=X&�<��!l� ���3,������)Ō6����L��k�$xy�O�+��6�O��ƴ�>ˀ�~�q����^?��Yjƪ�lZu��'��J`;6tPώ���O�M���c��,��l�j*N[04XR�RZ/D�N�8�&��HNc��:[�!)e���i�@0]i%xX�4o��9�6Y�������׺�Z�W�W�aO��~��tq���/e����!H��Q3�gP��?a��>F\���V%
��r���0 �x��=#I�44տ9M�<��s0�'��ʲ+����I_B�����~򿦙����e��E�l�F�;c:ཋW�g�����	��$�`[^���Yw�_�{��	񙪱�Y���m���i�;�����v�I�_^VQ��'aBӻX�K�Z�XyD�o+C������{�y?�I���6���I-w�>y�o'pf/5Nb/U|��<��x�bp�,�+ v������橇�oo�}y����] ��S� _@�g���f����}��#��>>������I�dh[fͰ\x�km%��k%.ӡ�	h:����zYh�)oBo������ (RNZ���_{r���{��kT�A0h:��s8��t�+CX��;� ̞V94��p/��Ԯ��w�v	��}~}TXKC	��ۋ`�C�K��C*C�/|^��|������D���J�~����gn�Ͱ����+7;�-�d�E�՜0df�3{'���k����-}	�vM�|�gV�j����SA����~�9Ea��Bx������;�����bP�z�T��u2_�5Ӣ��ɐЯW9�ƛԑ�V&��U���]��g̿��w#}���x������|����<y3�ԍ/�qg�&�&���+����Z϶�k��Լ~R��c�ۇs�?G�����|�}�������P^�)��Ȑ��i�Z��®�º�G����=���g}ǒ��뙮�w/L�n���mu������Ʉ?WZV�_+.��	��,�<)Nxބy��^gG[��w��5B�Ao/QEH���V�̜0=�4Q��Ф0H����9@&���x���'z�?p�&*��8i���=��Nҵ5�Cf���2j��/g8��;#Ε��5%gia�aa�j�t�9�0[�;����� 意�%�k��I:���Q�cY�}����WI�aGa��䡈��X	�J5�����S���;N����w���,�D��~c�,n8d�N�1����l+Ψ�1�ҮR��5��n,���G��J�K���q�-��/M��	�h�/2'��R��JZP",l1@n�v�d
&�Jς�D�E��U%�l��IR�G�CB�5��'9 t��c>�[]T���f圀�7q����b.#�lZ��Nգ� gc+���L/՗��Wl�����vK���_�
��E`�A�Ӿ)	}��Y�����;�������(�7E����9�=ʈ�C�ӛ���>�|�cbU��yb ���Zv �-���9EU�er�a@�]�Y��.?���Ѕ�V�*�v���e)�M*��,�G�p��H(�O_��&p:�#���%/��>�Ӌ�Ir��" SA��@5���#��H�eA��������u\+AV�[�Ɋ�/X������������C�cx�t�r
0'  ��#mcR
�����z1EU���S�cz)+ �l����=���R	��f@�.t(����e*R�֯B.&[(U@�׏�M]���N��)$Z�h��&k"'?���P�LBJp�h�#, :�NU�AŒ[�g>��b{]�RU�N�j��ֽ@ �U�x=�z�f�/ș�|a�A�28�OCP3�l�V��rũ��-�	K��9�B��kT���x6þ�s}�=����of�zy�?�َ��t�fU���&����(mJ�a�[E�55�Z�9��6)T���.�F�m��L��W �Y�.-Q����ü��Tt�2<@g�^�����t�mY�H����"�u�Pn���8�:�~uuPo ��;Q�����|�7�q1��0�v���p1�"����⌲�P�<\hJ��_�Q�N]�:ĝ�:E+zO]�â����O��c�b����B���yD��Z���y�?UW��#f#��F�P�J�Y����E��G����Y��H�޸/f)���52�<0�`'�����HA"�Ir�&.��)f�]}V�q*�T�(�mt%�Yּ���D"���NR&��H�#*x�A�)ӨJJ��b���@�������,�� �LHϙ�s�ת���o0�V`PwTj��.���DYJ�CU��iqw�<���1'�%L9=]հ��LT��;NF~��v����&���A�Y�PV�&�����+)'�GG�N������2h�
�c�|CC%��ݷ�+�r�YE�ߤ����yb\�hu��-.�. %�~c��_�$�bJ8,�F �%�n_���&?ȭ�c@`y�Y��i��|��#�P���`�?���;� !�f�~�4J�uw[�&iO�e���mܟ)�< ���C�-�Aw֍�X�fo,�Ӽ,D3�U\zi�* 3��wf2������#�¨�dh�M�H<�bYı�R@�\�9=߁ޗ�)�9���꽐ꔱ�j�(���/&����F�GkX�xnG����e��{(�I��2k:�*C��89��G��ű�qq(��"6ᅘ��'�B�D�����3�.���,�~��!-Z@��ò1��V�j_�
D��*�31����l ��lZ�DW�Bvu��Z�t���Sr�RW��¢뤐��*������#����/�����U�4N����U��-���ud�g�J����0��j�ׁK�&���
W_%�H?`�F��{��i�����G'~��o�"W.m=�
�:<�{����hfΖ��b;"�?5��縀ǋi��-�"u��W������os?�c��I[@��G�����3�~c����7_w����d��j�fF�MA����߸kH�gtAK�.�}��w�c���&{j����N�׋?�xD��p�jPeʧ�+|3l�o9|eg�]�g.:�N�Bɜ�fq��-Ĭtu���u�zyrd�^���}+J�EǴsB�t9�B���<b����O��<�p�#`؆Y���$��v��u���[��-�= ���cb�w�U��o��_>��l;y7�_w�޿4r�?�_u�0�־6���w�OrcoT\U���;�MmY��7\6���>�Kx�����ă��̊;�2����P�ב���ޚ�m����ݱQ��vjSS��YjI��L��+����|.v%�J|_��}�*���P̜�e��֦��vi�V������&@�T�uH�c+[���aE =�Wҟky�`Jj��[ ��N~��Y�k�g�k��&�ɕ��[���o����h��B�!Q���]�亮��[b�����,O�Y��
蕩{�����F~�ǿ#�3g+�^/�G~�X�W�x2�4y9���di�^\T�ǻ C���>[r���u�<O>Vx�$O&&����]�x��D�ԛ��a��'�Yy��߷vWƣ&�
�Z�&5Ly�}��Hr�����E7�B�夠L�48��l �S6�"VHХYUY3�ԡ�"��LT��Jý��j�F�m��R,Q~P�6�@�v�S�g�.B���s��'޴�^��E��Y�%�V��@�^m��9U�� 3��;�1��Q�>�&�F\���Rx��ء�'��g=b��`�ۊ)3j����j��\1�s�_w�j�J�)A}KS;W�S?~�s�e�ii��;��JK�NI���l�k@tխ?�JuF�$^�~�����Ci�b&g��R��!�$o�ZgK�[�ZS������3׳ą� {�t�'Ԙ�ב+�ت���ZS�R�(�"��<��r�^x���'<�h��,ƒ&�.!b0Q��z�~Rg�|Z~�o��H^P�猙 i��Zg�G��[�'$J�-:�&%�q�>��'�uU>��	�;Φ�����i��0cù~�5
o&�� {��+�5R�x2������/�^�N,�a:ZY��H��rNvj��2]'[���!�M��$�� Z�R�Q��lY�hм.���Ҁe�����Ҍi&;�z�����m[9����)��Q�ے�sLwq�}?�nS9�D+P�:����'��n͗3���M�jސ��Ay��y,�D�VZ�t�ž�`�;��f"�hG �*��zj�\J8��5�``�z���21/!j1��P���N)s����׀J�������i�;$Rd�W�/��-_�����9�mL�V���/?�ĕ��1���JXC.��o��(R��19���ݤ��C`.�8����t�9xF
�0m¤�2�!q��ѰàxP���iq�1�$[�g\��hB
��_���3ֈ��rW_�S�$zKOk��K2X�/t	�9�_ ��T�m^r�ߪ�qUq�or�#-�lH�Pj�����3�=�E���~]�\�d�h��0xx���qD*=�%N��~0sE[5b��Q�['�P�f�l�U�ubyo�� ��0�����Р��Ⱥ��_�b�]�e�'���D��E�3<�����W�%�Hi�v"9ݙ/l>9�<�L��E�h6���=�a9ZMrA�{�7��XV]����!��D�Qm�p,��(�mN���I���ɫW��#���$	��>�W{\��zaS����h����bFSj���ZFX��Τ�����)cIT��O�ф�Xg���Lm{3ho�]ֈ=�!�w�����}��驾_3ЉS��u=�ofl�@>[+�R�K��P��$���,��cf�	@0� .~T:>�P-SW�8�	B���u��3o˧�Ɓ�v�D��VrRZ�x���x��K�C5Nѽ��=��ȷ����$�}�8��E8�!-��@�Z�'F\a�Oe��;�Qvl��QHCf֢��YÒ�V�[x�?��^m�_�S1�C����W&c`B�m���a%�(��+5v"� �3[��]�t2�D��:�3�=v�+�4""eD: 1�����Qqz��eJN�����U��R��\��s!�T%��1.vFf�f[Pb��d�`����'���k�X���|h4��w���9�>2�nT�"�?z�� zt,��
[M\����ilqy�iD<H�AbÁ��]i�tZ�ɝ���	GhL_���q��g0#]C�I�H�-C&��\3Ļ�Yj%;�x���KA9�_=���x���B�~�u�j7��r��pE�6�?M5��bh�Q�E=��3�!jfB?C3:�/-F"s�1�� ��f���K��ZY'����3?+�A1VR]�$V��{�ퟢe�\�u��pY�͍��W�?8����T��yѬ~�)nѱ��LC�����w|���d��~	��90��?��â}O������k#'</�~�����-�Zh�̍H�o����Q�A_��jߪi�X��ù�q~�>_�Ꮥ��9�B&,�ش�E>��h+s��rK�����`K�Q�W�X/d}�ס3��$���B�ͦe��b<}u�'Ns��d�ȿ?v�MIf6��>=a�Y�^L��ak�y��*�Jx� �ڛ��޲������}L�ю#.��A��ʍ�v~T��w���Md�H�Ī�Ku[��������vtR~F�W��O�4��2/�VV5�_1�t�D�֋&�4l���Bֽ2";z�6?�[րZ�c���7��5nq������m:;�;ְ���&�*���ω�.`���Q|M�i5�ji�b�p��OW�O	>��{ib��o���;����'+�Vy�B�_qg��*[Vz�}�8vY�?"c��j�/�Zn��|W���o>��J�"(t�*6�����w5�5�4^��9�������˥�ͽ�����[)ٽ���x�n7���r����l�3&{�.���<�y��M;USU��� �: a��i�)a����ww2�n�|_���c��Ŏ.�g��d���ѹ;���+��M(�taE��H�(��cm���]�?r�-���ɥ�o~�%|Q�^�w��?���kŨ^rVt?��t���6���ך-���.ۿ��CI���-�S%d�َ?g�����]��}~�/0��f��P����saXZ�u�.�]O!.��f�`��-v�/�>�-�6S�b�ڹO�b�B�@,�^���D��H�T�;VNm���O����g��5���_/�^��`��4p_	Y�I�:�v��:�m��?�d@��i����E����	,(D��i�K��f`O�~����tJ^�B�f��~Âċ��	9��l�Il��������z���=f��au�уiMNA����F�r�d�y���F���b0ӡ��l��w�y^ō7��S�>	��8���F�ՍN�
q-�|��Ӻ��JQ�F����}�L
o�p~Xg7����
Ύ��)f~�!l�"
[�N��4�h����._}]�5�t
"��M�xl�n�H���+7��0$v]�̬/(^~�(�*V]���7�2��/�q7n.���G!!BR���!㣷w��_�2��r��'oZ�w ����j8�7TH�M�t�+'����ã_�a磗��e"C�x�_�ݏڊ��o*8���wI�=\5\r���N*xN�D6����d�;�V�gJ�����k�kN�����2Zn�iQ��ٛC뚊"���$YY�	UݽH&G0 g.�P%6<>�`rm5��;��u�|!B�X+���^���B$�ƒ_�QXɪ{A`2����&��=���>kO,G4��Zf�<K[������(E�&�,30N�f�0@�`1���C-
e���F%Q�쾠ھ��ʚ<W6S�	�i��{!��N�����8�f��b.>�Q��h�0�7��X(�r(`͉�Ȭ�ΉN��^�uV�ac ��;v��j�\���W�"���w��bg�t<��^q>q�(?O,�"���y��TإWNVtc%a�p9:s�!�#����I�c!K�c>�*�A��r9umV���Cy�[��d�{T��0��W�E���X���,J�o��C�MAY߈"c�;�^W\>��DJ�n�pu�giH'�(�5o�sQ)]T��S2=�C�+�`Jpƍ �w{�y�k1�����jހߦ<���I���=|
�6��> ��6(W�sĭ�%�їC�Ǚl��a�1�^k�w�[�`	Bc�ٵDy��J��RF�{fcn<m��R* +�%C�9œ�ʚ����c�F��]�7��-3�Ԅdbt�!{�̬.��Tl��i��u��aI[%���E�|)!@z��AvY8$���W8��?��d0��9�M��nƬɏ&e�w��۰h�!p���*����P\�;)I�o'�B��6h���=2��+���wkF+�B�ұa�� 3�3q12ip��q��<���Ӫҭ�_9�]��r%�3E��&[e���P�o�8b�H����JmI
��bu��v�nZ���, '�)*%!5��R2�ԕ$QLp"��X<$J\'����;��Sc�-xs��vx�"ށ?�'�@�=��Q8�EԲ�+�Pg̈���m3{hC/�q4k-{yٕ��k�aj��(kW̪�nܾ��R���k�	�)GgQ�-�~��7���H�\yP�4f��m	.�]���+x�oDwD��X������V��lIV�gKHe�Br��gf9"��8!���tH��I�R�{���s\�"H����U�"�Ѽ�iş�+Zf���f�4����N􀬅�I�����Qx�W����d�-���L��4����k	T�竅 ;U��HL�*eIa^gQ�����>BM:�g��s4�SjR=��h��D�8O����ol9��7�-�!�)�S�J<j=t�!��2���a "4�������kNU4{�a�jlz!JӬ%i��k��rm ���rD�(&�"V��	2:���'���^L�dv2�� �B��ʚD��M�,:-a���,z
fw~�Ȩ|�`4�� w��P/Nt"MR��T粲qH��6=�CR�N>��Bt���4�B����6���]��䴀 B��z�Ϛ0E5���9K�jO������u�㫐��y�Z+���3�G��|�c�͟�>�.��������J@��~���/��χbU"�򕫦��\R�O1��)��Em0;����o߾��ZF_����W0�}���\� �,�ҚK��?�1�?���Z��&f���$����_��_{��	⑬�|���;��
/,�������ɥ'㿅���=N=��|��U�"��t�{��y�鑯(OȽ��]8{��q��{����Q�.�E�^�=��w�G_n�^��ͽ��K^�����vԃ��ڥ���co�|���,s�o�\�����@{M1+��a�,�:I k&L�޹��&�	?����E�V���$�X�e5Vym���r|:j�'�|Z遯Gո �K��� _,%]��� ��2m��D�����Ή/����&߮�m�E���k[�������
Og�w�ּ�R�����F��A��4u��=8_�����ث��ݯm_{�������ӣK�;�!�:;9�J��x�n�SWԉnX�G�N�����cnmr��ܹ�l����;F������i-�Z�+�vL;�N���u���s^a��"q�0bp�u���)b�'�8Ď�W8��Kj��B�{���J1�띁
�E�z����h��C��ݻw�ՠ�Ȩ^+��~�m �y�^���X{��o�������K_>������7֬vwsuɿ��Ke��9�9?;�����Quf:g���g��Ʃ/nYܺ�X�˶�t�|ˋk/�OWg�[������֋�I��L���⛼��'[GY�Τ���3@�V��X,h�03*�&����)<�`��C�p��n�h�]V��I4��l�h�=�T"�Y��(��=�~��K���y`fac�zY]������⢋���!��iA.Qa.�Q խ[�?7n�X5������ޞc&\T�ށ�8~Ϊ�N�[3���$��"�|������"��0����1���$�����"��2�{��ՓB+�L�j���u��W���2UuCp�iZ.ף%(^R`��	�5X���󫽦��]�5D+0�����L,O�{+�@sԠl�l>�!�N�7oޔ��H�aW��Ѫ�]�(!��b��5���HL�C���������/����'���bD.��4���rY��$��Qae(	#�:eQ���Qg)T�`S"J
����� $��	�;���R��������B���UB'��2��,avF�PXx-�b��r�rYQ��3���*֨$T�g�OQ�,�52��Rv����eA�Z���J2�[��D�@V7x����Sv�
�.^`�0�������Ka��J`:H�j(�o�&0 ���Ȃ���4���첳��Q�,]`��ȺJ�%*�H�����b��`�()�6b�Q�Y���4�#ES.#ZHc:�(�X�Q�,�Z���`S�+�tFx�n�\f#1-�Se��\ ���l"�D�/;���,ȋ��^�YF��8M)Հ�a!t����ou�	@0)`�"y�9��}���"SFxH��:�8)0\a�0��&W�Z����j�Y`
Ab,�bu
./p����+�k��͔�l����<U�	\��U6/�Q1��E��JQ�+�l!x��t}���zE�� ^��0#oI;	���@* ����Q2��*B����*0V��Z 	�LS�QRcwB
 c;�BJDi��D�$2f��R��B;C�ʹ& �D�p�RO{�֢��� �� �)���Eo��%5V*�\,F�F��T'c&#��;R0c�N'��a����+�a�%S�(��+ʈ2�ǱR�'o����^�-�
V[
L�ʋ
�\E8#��u�,1BY���g$t$��"7%�\R=��Yj{b�e�'K��-�Xv.`� �͒ؕa�H0gf��B�ɒ��RH� ��k�x2����`*�Ox#<;	��S����t�bL��n
�O2�+i���E��E^�����*Fb�҅d�YZQY�R�ȅ��[�ʋ��p�XK��Ei	�����p�Pf�*�+���Ei��Q��|�`�.�)$|^���sU;f�v
���kF!�b��	 �@#��\����%$Y���R ��%t��{�,��BX*�
��VǋD���3j/#%�(��%��*�J2��	��F`�t##�`�w5�� 0���BK!��e7e��즥kd	OzT�!U�U�)��d�,���X�FF0vb��K"!E��%rFR����Y� �]`
@L�@2����+f"�!}�lJH�'�S$b�����,�8�� 6v����Q��j�ބWv:o�����V�� j�%�٫�{:��R5P�+��l�nh2�T[��@E����@
G��VWl�\hJ�%ę�HT�Ќ��K���W�(�#P8
<��t��W��s�%���֘�-G�Hj~F� 
�'�H,�@�@.В8U.��0�"�\`v�ȍ��X�X�)$�)iZv�ó`�-��di��t�)?�1�30F��#��!�K1�
f**~���F+�+�UT@���C�yIIQ�mF��Q#%;ET��1`F��\�$�g�#��H?h�<������`���-#NG����-�H�r�% ����)N�E�E�-)Z��ؒ!G���<�4�p-�B�8��V�����O7��<[ml�6��љ���K/��o]�_�]�����/{q��#��s�btIz���o�'�{�(�7[�#�g���������ݻ�z�����֐�����ID	��0=+�'1��%�樓癖ߓLT�+V����&��'�J�
��%%���Q��碼�Q~��r��I ���w�~�*������'�nP�˂�����ѓOx�b=P��x��m���~����������N?��Z��g����X�:�?:<�?o�6�<<������~tj�v� ��>���Mǟn�Z��M������Z�����q0���.��ܚ��k�av�����%ŋM��縩*K��i"^7e�����L	
9�B����h�px�`� �����������������͝�u;���~���ln�C����:�a�:�;����G�����{�雜7.=��ʭ���?9��h������*�Z?�?�?ՙ\_��ܓz'R�t�z�F����^*�î��p�t�7B�p������w�R����ť�3�@8�N��`v%��p��N��η���J��6�;L��`�dwa#�D��*�.	��ӟ��?"`�(�/�W �^v����܇~dsl�崏*/���e͗��vx����m�\[��o~핯>ig��ӵs?�l�_6{v��^�~�>v���P�o�w�������D?��뷾K;��˳����v������mmk�tl��z�1n�>���?}��D�҇��5�?�x�#o��������¥T:����B7ВH�� J�赋��L{�G���`J�r�XK��Հ�a/�THK���fSQx��-��+?�,$#��j��z'F=D��]���ҕ⟊8���S��2�Uo���?{�4,�i��"5Z'M�����*HgUmF���R�3�`<�{7���r	�!.+0�.
�
��b�;ܼy��!�,nz..���*XKƉ��Ad��os�u����.Z�(�⭅RC��d���L�X���ȹ(H�!��J
<���ا�pe[������Bj 6���mG��Xr�2�����H�{���o�m#$�n!>�yY,�?�P��X�\8-��.�����V*��SQ ��*��s�
eqGU�v
�|`w�u�׏�ŉ��I�ITz�N+R�ضXCD9���-]�8�[>E��i/�X���9�p�"4�X.!��Sp��\	$<�PL�)H,�H��:c���G�N!�22Vj�e*P���EB)�z L���K��V$�����og��F��i�h���%Jm�J�y�?r��#��ExH#f�ƖIAU�FƘ��F#ZӋ��.5Zy�b��1�%hy�p1��,�F&�\�����4E N�
�Wx 'E�`&{Kl��ed�Bc$��	@��v� ��m��C���nʮ��D F ��J��Y<;� d?S9���,t`����s	���8y�ꏃ7���qÄT*}�-^T.� ���?i�14u�XH��1Z`z�m���
���N#����,0,�^�ҹ(�T���aK`�F�OL�LfQ!����*�v0c��t�i�u�b
<�,!�$�R���{'
0 <�����,�E�"�3;$/N#�	��u6�X�
[$ ��P����| �L���m��³�.#u�g䭼��b! �����Yj����*����+^"i�9���t.�p��Ś�b�����e��[;�)�-�����c��XU��xL�FEgo���b���,�=�jnC��P���R �@���T�0��L/���I�`�y��%p�K�\�.����i������ϭ�VH�U��R���2c�^ce���F.�80~ ��N`�dt~�����k,%�bQ��5��C����DF���
T�(c?�C�P�DOfMc,#*�v�����+�OF�����EPA6"�0S������z�h�%�F1V���	!c���2��e1��eOn � �/\`Q���Y[: ��-�����&�>g7�֐,��2J-�V��j��Y��`t�����`,�XbO�y�MƟ��j�;��%�*����F�����P�) 	������U��,��
�����+����DB)�)]T+��+���@^x� qh�-=����(
�Xӱ����6�0cI�H�|5u
Z͉rȲ3�kVU�0� Q��^RS"5Ia35
��H*̘�Ȉ\Tƪ�̎$ �%��J�% _Ƣ ��D,/]j#�TI�E5��#��b�J�^��p�C���@ټ#`�:/K۔��(���N��
1DRR!>ь�0FIM�2XY�p�m���X�����uGu��2�@<�h=@�D.0F�n���R0FR��<c͑q.��.  �F�� �E�s�);�n_��B�M�gk祗[Q�)���9XS ^R�F �`���%vJ^�Mڋ~#�\�-�X�b���S�(���	�\�(%&v��tFA��Ҫpfd,i�!�`��b�4Ө�BJ��"#Yx�X��F�،�O�,Rx��~
��Jo�/56!�FzS�u�2F�ɲ���
�N�D(��x�)�),�,��  II;H`�`������.���e#�Q�13���ur�C���.U�n�o������d}������~�o�湗���⫗w��C�����/�0�7 ՠ����k��晡Dn�*�����+}���w߽}��7����o=a�c=�����$�
F�V��TC����2�{8���ߟ�{���לRK�ɡ2����5x��k��yB+~Q8��_�U:�T��B.�#{���}��/>!�((�������o��St��z�-!��Ͻ*�B�̺�Y��>��_M���|��B��N�]Q�W^~�ٗ��y���7����~3暯zD}�wo�S�~����+q�/�D�9F��NUt-2%�9����3Т:FƦ�BH.=�-1���.^�2�-"��~�&C�P�d�������(�0��2	��I�M%Â�6�a��S���a*D �P��67���؍K_zg��4�\�q�w���.�C�}��)V�Q3q�-��v�S��-u��ӵ��K۾���5���K�w����g���G�7NW~�����S�sӅ7����Y�sc	����ßxC�|h�s�YZ�/�VGw�y��y��]��rL)ǽQU�q�=:w��y��P3=[��q��#q�9�bs{�u쐺�b�r�!Q)O��f�*T�����'��\���@5�lW[�u��ޞ�KT
����u��Z��6Ϸ��߸r���h���_��ó���w޸��?�y��:����:�Ԭo[��}�U6L��8$�{��T��8g�+�Xg�g.�� x���n�N�8<X����h��������r[�r�:m�r�/�p>��G�4�8i˥8jxz���Xv0d$yz銵�]f8e�E"���1�����ѹ�|H���%bt��B��"��Y�:��)	okׇ�Q�s�<o��KĚ��Mv!���+��RaR �����9x�Ĳ�Q�#���\��iu�qJ�8���-���UBSY�\�q� gRa����8��W�D��]Y���>�@�4(1W�&�0�P����_@W'����:�@0�E��X���b7��>!��u%*[a�2Z$Nv��wC� P���#� E:{2b@�햬cF�[��~2��sS���O��3��`�a�X�#ʰ^��b����^Ԡcm�:�ڤ�c��O��2T�b�'�ƺ��m,�}$�X�Ά_�� ���uX���YQ4A�;*�N�QjwKc-Kf�yQ��U6 #*I�`j �ת�\�<����px��h)���l�0���"6���*X5D_y�,�*�5�)L��!�I��5��$���-�d@^���q �*0O |�\���tR�B�s-|OnJ��Qc!mi�՟1�iK(��^��Kg�B+�1�p���[̔J��۴Q))�uɒO%�Jm��_�(�!#x�Q�j��*��3��˓�������.�V��Y�� ���T	�) ���M-�X�\m��	|�&u��ȹ@`�1�@S�0����UӍ �,���BS�):����2�G��F
�2��r�զS xu�NZ#NvJ�(�b�
X���4m���d4�6��g7M���MI���7Z �&�MT�#d+	0 �!��,� )�>�J�����(�x��dD^H�s�t<�Q�`���H��pU��eQI�Q���M�z����R�Rd/�c:3���B�B �MjS^�UU$�b�M��3��BBV�RF�a�ԴU<a��)q�g����(�F�3Β.���(�(*���(��%`2��RK$� \�ó`+E�����0�`�|z�P�"x��#7X������T�%�$�r��.��\�e�TP�; b�,b��R����b䅩�9N���
ϥ�,1�~q^���Kl�@z?��yuL�?N��,`"�p�n�X,�:%q�Sv����(NF��g�+�+NFH<�!MU+���) 0�TH�P�\>�ؑЍt ^lD8��؉p�F+;�QTU�����$\ �0SF"�,r���SX������Uu��h! ����0,�jZ��*$� ����N�5j*ۤ�ڨJu
�\�4-{��P��g��R(��S��� ��sM<#������-� ^v=����Y�A����b�D嚀h�rQ«6fә7/;I7��)��S�a�f�b[��tF�B(�浃3c`���    IDAT�5%�8ڋYj�4��\�\,�����J*cE��j�^`�E(xĒ�+K�9Fn,���a��4��������i���;H�X�x�d�WyI��Fa� V�+ �j`dԢ\M�1�֢�QQ��G��U9kc���<�L��Vm��QG3�xH��K �7�Z��*���T,F`�0���Њ�}���N�a��)W#�<�����,h�T�Ub!����	)��ڬ���bI����>����%D@�[e�����ˈYL�X^�T$]I\`����RR#Q��(��|���kLbk!�B�E�DN����B���&�mQ�$- �p?Se�[�Ȃ܊��!I#/c0#�)#�>���ȨOG=q�]�-���y�����n��./��9���Sw��,{M`B[������㤃�`ʎǊ�Q�F6�앇�.06�a������f�,g� �J�N\�����7.oo���㓃�+�W>������37n<��G��~���7,~i=��L� *U����{�y�(�?Q面������~ �Cj/DEy��$�F�a����jSx��|����كe���sTY�(DOl�z,�ѫ�2�a"�Λ7o���x\�	B��-	�E��V~O�=9�㡥(0<8a�߿��[o)�K����2Z�Ԩ(�I�M.���P$Z_�mo�n�oܸz�����S_����\�q^�b�==ru����n_>?����7�W
r�CM�,��l�%F[`��E�cF$��=���	��_`
KP􇀡�%!�w�k�MԴ-/��]&[��*Z)]9t\���і �s���HL-,;6�E����Vg�P�7��W'�����#-A�F?�`LHX���fZ�tW��1��c��~v�~|e�=�o�}�/�����n����yiu�����G��⪙x�ݻCk��g]��#Q����)ɧ�C�h������$Vs=������q��w�Y:���`׀/��NB�k�+�6ܽ{�ׅ$��Үo���eQ�m�\�.	�z]�#G�f�.�p`�T`5�?]
ۄɯ�k}��ש}���{����������������>����g����{|�w�����~�7��¬+�_��~��V��~��9	��W���oi�(1�����[s�[��=;:���g�|zx�������G�-��_k�ΔX�Qjb�d1;�J� `�]���4e4�S�����T��8~��h��~9E �9	�8	���30��W@�`b������%=f���l��)B�+�Ҹ��ax+	��:B�h!����.'�.�Կp���)�9r<���E�r�cp��e��/ʱt&�����˛�[�nI�
sհ��?�q�Hg/��@�Hg<8��R���pE�V�E��"��'��t��0U�����˨���,�-t���wx�,_�%�.��E���t�b�4J���N -�Qg�Y�K�.�u�/#�K��Z�5V�
M�+�mn�M���{���0�R�4��/Iea���Ks�t��a�"�Q前.�XK�K��ޞM�4�b�u�{Mb�|`��p٭�{����E����I��/��[�R��R��+N��Ś�S�@�My
��
�1��	/�!�� XE�tvv#�@F��\�b�I� �p0��`P�@y+L���`��lJIa�a�`��#1��R 3�D��C�[y�5�E��HT#���,���XWg��M�)���5�l"SvJ�1-Dy�H���Y�7F�O���4Q���"ET�bf/��8�:f_BR���!�فŖ���W�H�|hN��j!���M�d�!NW��	�����H�E`��⢨<��a�eɋ����8�/Ț#JFJ�;6xYb�+	/����9��%E����ᚴ#���Q��ZEF$8�1��\Jj���YK�፤��G�$�p� �H����WƋ�錢Վ�*>�m.���R,MH��j�ď�h[�X�Hx#�T�)ŴΣr᭝Q.޶�΢¨da�j��t��I M1"Og' ����d	zrA���s�o�0!qr1��s)��,t��Ԫ�kJ��y���^W�	#��>ښ���Pfm��qVI�e�E1��t���[C+*��@�b#��H���ϴ�5/��\{�6y�H���XKxH0�i!ט.�S,紈��,�T	#��I��<|e˒@
��z�1*�hږ�����R�3�!�����.0�&���U&��,m�(�.��
Yd�F0RTJ���$d�*d���@��`N�) �e��J,�:` �����(���!=< �(Һ*Ɉ��` �-:��EN�bo$��QU�D�z�|�X(�!�b�?F��B�LDS�
����@����X�U��N�U�`,JTU�a�XV6	W=�>1��(�X!
�,��^/`��$ e�* �F(u#0<#r[�EL�L��֒���=�Y|�B|M0�"u�jzc�e��R�#*�	�i�i���F�$�f,�b��N��*#+#ɲD���d���ﲲm1�(#d��<<]��~H�Ƣ��ϒN���"�䦮2JR�\`qD�TH F�8��ˁ7W5�^���QAb4-$L^
~z�q�.R\���PRv�$vX.#o̒R�,!��UE2�s	�e�\�)c̢��S�L�� 
B�b�U��XL��h�Z����(#��b�,��c�`����<��|��"/Qsxv�D%��1��E%��
QS:d�h�������&#�(:�HX��
뿵]5t^�td��]�"���)��FAI1%ca���tHK�`$pS� ��$*�B�rEh#]y���G��O�e����gT�@G��0�
I��D:S �،�e2R���HAU�f�@�($;��0J2�@Zo���� !��ظ 
�ƈ��b,;dT���R �!�*c�R[��p`�j�
.$��:O����13b��{��H!a��Ffv�#c�)r�5E�Q\ed��b�g̋�W�#f��a:�?s5��\�_�{�����?��|u�sşѼ�i��������o����z�'��^��#���l�"���#>O��~�my]�� �/��/o߾����Q�FQ�O�=�p�"�}��w��Kv�\�%�͛7�ܹ�9��c/΄��=� e�O��z(�랶��#kea����{<6�{�����y���/nx���뵢������A
��ˣ��D���;_|�9]�B^x��k��<���Oݽ���o�\��y�چ�ENּN>�4W�@�x��C���Ϗ]�kO>D#�͵�5�3S��B���q�(DO�A,
�o$8	#$@��+uT!٥��E
�.J�w6x��v��Њ�i�0y�m'zn3�S:�t�a�S���L��d�[�mL��Q��ʷ��L}����tc���j��3��~�>��ž�2Ӆu���A.j����?�ч��7�{Ƕ^��NN�����پt�ߝ�z�����������^>98�����s7����/�v�����R���9�{{{�9[.��S�-X=Fo4{���՛	�-�֭[.	0�h�X�a��,�qeq���������k�Że
g����G���7+
C�L�=��V�S�۳{�2�`�]�v��}+��9���p?z��'c_}�5�5}j�ﮝ�����O~��h�_��پ��+Ͻ���_�{a�y���g|M���xl�景��^��h�Vy鎞_%땴W�õ�q�fڱ�?r��eNB�߬];�r}�����_<^;���e`_ u���W�~�P��^�|`�K�ή	��bٳ�,����Hg�H
�KBH�z�)A2p�O�������ڗOq��,��M]�!�.����RP�IS�]�ۏ ��VpQ�uk���D-VjGx��.� VW��0�Ӎ�E���2���3���d?hb.�	6��(.1n���,����0�t׈�j,>��[.��%�@����Ũ!>E����ߗ�
������	��+K8�Jԉ��U]FW�aRP�� �=
��q��:#�U�.s���,�}@�T��Q �,��H�w�H����%�k��b�X>< v�[նAJ25��M�č%�;���"،�x: K��(�����s7C��.F�%�t~b�׏��]�*Z~��k�v �
0����n�;!y�ĥر�޽{��=g�1 ���[�o�
`T3��B�h� )� �
������; ��VNH�v�����@ ����F�^~|aW�@v�·�pzU9�,�+C`k1*�p[ 6+�^l�*���G��DWLy��e��0� ��0ZZ�PX��0�3��`�BJXz�4%�a�Ɩ�����gRe/�b��eCWX�@�W�D�ώ�+}�ĲT)\����Uj�I�/���t�v
,ݨ�������#$�e�E���-D������:c1��
7r�����@������ v�j���8`�V��� S��V
:#p�����K!;<]8)�d�WH^0:L%1��	�.�Ύ�I<���DH(��Ue��$c���H`�\Fv��#AK'\�,RS�6嚜��a��(����倱�ј�Q���[K<�p�6Hb��B�����s��P�����,�� ȅP��c�*�q6ֱ�U*��5	0FR ��SeLW��S)HH����c`1"�5�g�Z�t
���ð3��P8 a�w�Մx�b�5d�h!��T	oxJ^S:c@g�+�bR^��ur��n���%�m1ox:A�R�Q���_I�Q�d����Y�+�Ύ&*50��P������e9�)�p�B��^4���Y�ت�b,��TC<���ltI%R$�O$FR�\�춛�!J$��	�Q ����b$tR�qbcmz�F �G	oJ��%�ᬐ����F�N�b*�� Go�(]�e�V,�,d�m�0E^m�`�(s�t^$�)��]�5�+FBW[UA�Yr��\�'|�F���V9��HŘR�������=o�r�s���W,�H �鄫��1�4#/)����1�0�
3��d��GF�O�[���eT�<�DlH�a�Jj��������������y3�[ h�#�30M��CIY?� &x�q�U?��G2p�3��Ϋ��Je�/=�ئ�Y�O�"8�f�o�a)*�RC°H��Y�*�켃n��c:N��R���C��^m���8`x �,�3#��Q��D�b������Rx�`L��+B��x��$�
C��F�R��2��KG��bWa�Q0e	��
f=�W���L7%�M)��v.�D%�8a�x$;�X�i:W
rSZ��B<F<)F�,�BJ�=]C(EI���	W�Y���1�ʑ��a���`�Ë�)*��VV~�o4ej! U��.d$2Vp��E	ig�F`�x��y*Q��c�V����\�V*P<$�L�2�YF�DE��� 
0˞��/;KK�U'Z"\=)x�c��Da��#yt�OH:�H$�P��C�ԅ�j����*�}^j�6�"&#~%�Y��f�FT��J�� 3.�iT��l��m�U�p�vF�rQZ;f-c�!);�m�t�z=��������tTT���+��(by�PF�S�]��%�Yo%5�Q%V�;5��I��_v��:���-rA�R �`f!,D1t�F�VGa����Ǽ>��vzx����!�~��x/s�w����W�ݺ��֙w�����[�3&���W�����V�k�~��znt�o޼);��*�������[�n9ƞǢ�B���A_�t]ԍ�qh�����b�|u:��hw�"�M�'�?����%�gJR��ޞ���^��a�$W��<-7���n�t�x�jQ���	V�$���?�������?��o>�P��������_������������kg����x�9��v��ٴI������������6f�H�Q1��x����L���돪2N�(�G�M�E� �Ǵc�YD��U(~��+��#�b;D��G��i���c��'��	v����J$���i��˄��� �՚�	�I���u|tv��͓co/_��qx��o���٩~���%������/��E����˲�����uW�闏��mn�^��W8�\�Ƶ?��ͷ������m�:}#p�/Y����O>�\�T��Z�s��R\!����At��{��;jw�ޥx���HX��8Ц�iWZ���8�����������`u
x��p� �u! �̕�����/�,��ѷ�bY��b����֛�lw�ik�U�+V.WH׆Mqm��G����6S����xp�����������7n�:;���_���W^xf叡�?�k��}�x�i�����~m��e��I���6�F��Id}�͏���l����d_]_|����7����m�G?(�;nl�휞,o������v茞t8),�cF��@����ԄFݠ�J��i�)�͍��:h� 1�lZ�`BP�������K�t�!�
4ڗ�NXN��F��tW��\�����t!C�rf�(��+�iH\����]ءr�0��۴c֊��c.�Q�N5/�N5r����w��t���D�~8����3��ÇN���3Oԣ��Jv�I��� x4�?�� w9��b ,�����$H�zb V?����]�Fa!� ��gv��.�S�T�NT5kE"Е�Pa��-�)�@��~���X�8e���X,J:S�s	1����@*�����
�?��&e%�Q�Q1�u���E製[���h����g?�YI�th�|���P����`0��%�D���D�v*ԩQ�h4�Em��b1J�01�������>��+�HyJ�"�
L��S�e���0�	Z�Dx�y�ɦ$�rхб��b鎊@��F`J����?�/�H�C`:rb��}yMUF�j��C����ҥ��� �BNE,{�Ӎ$�ty)F�Y,r$�UR,��	{�Wv���x� 1OB���C�Rl�xJ���z��23p�Z�؀SJ�c��WT����퐄�³@�)b�"[ ����su&�UnJ�b�RO^Q���R

<X�B0��VCR��_  ��
ff��XF��F�e�NT�fx����H�s(�"�@ 
L�M�2�B��Vr����HFl��R�"$#ǲ.#�� 2]����켑��%����;�Q��bJ�o�ƪ�y��Y%�VFQ��\H��Y���Q$N�6�@!,C#<#��%750F#�RQ������ +�[:��(�H�RӅӹ�Q�!��
o���gF�0%�Zz`�bSOY$-EK�H3 �(�(�<�S:
Lޚ����PD�4�0�'�p�Q KJ#0oe�D�f�%��\ VD'0�L�ffxH���r���II�>��Y�p)۔gL/�($0\�����N�	f�?��+�e�ڐg��tY�(�h��c�j�Ֆ'���?6�t�X.�u>Y4!�(5��v5�&*Z˧�i��B"i�)�M�O0��sEK�e�R���\0~�b�Ӫ�c�Z��S�!��:���d۪���Q���R��p.S�D��'BFl�`FR�2���򩈪T=	��CN�4�e�TS�[~F:B�V#�	�S c�0�[N5 cC� �:�)��H`��1�+��B�� �p�8��rl��T�ԣDU�!��̘n�k!�X"lT`Gk4�H�E�R����b�u0F�� =#�"P��Yd$�Mٳ�R�TC��(r���z�(��'��P^��F����M�@ұUgvFV #�
㟕P` y��y;k�f
W �@r1g;;S���Z�$$R���Tm)�ZW��T~��e���N�S�ty���"��U�TF�q�#�(��`#b��2�5C��Cg��8��rU��g-y��|HQ��qj	`�����4�tYVK�.T,��k�)*^�j0�;$�����R�$���6Uj����,� %�0/]�y5�3-��XHG�RMu[�j�I�/��,�_�j+���D    IDAT]�YIN�@�-Vah=��@ϵd{r�e�q�(+"S���(#�S�~�񬀋T*���;0=F��D.%��|���`�����{ϣx)��y�p �K��e�� �Z���Ig�9f�R�x,#��ݿ��	�n!D
�������<m��O��EQ����-�빊Fq� *��Q1����L�X�!U��~b� �x�����㡀!Â3�X�p�N cS0��R�h�ؘ�"aX�H�$(�S�qiEUa�@Z����vӴ�ˎ
8	�tb���3|�ʅW$~O�V���Y,��v��<Gu~�w��z*�$�%x�qH<�3vB�I1HQ�,���>�T��R�Tƭ�����楥�5�q�d������K��y��g��X��ӳ���o>%��Wm\l�<����>�d<~��M��@"wxTFQ�[;��-��e������/*f]�ԑ�A+\\�.[����{MxMï'��=������3��?�f��S.e�\ޞzF�UL����T�Sރ���~����l�[o��+mRO��*]�X���ŏ�2�Sj�&R�j�ĺ<���V��x��䗿�����現x���ľ��_�{�?>���ֵ�1~���e�n�>�Uyzr�~|�f<��̵�vx|�M����r�l�v���F<��M5';l�@ˤw�0��� ����Å͘�U�0Jr�
t��30E���@��,��^=y�3Z��-F H@��PB!��H��\Y���	�('/�^��j����Ǽ��G�>��������Pz�u����x��o�zm�}�}?��.Řtqsc�|u���~��3��t�y~���������+;�����sO����������O����|��^�-���A�z�褺��;w�8s��W���{�����5:���[�^Y����}w����۷�6��G�B=��SK�K��6����}�]!0�5Y��*�Y�g�R�0��R����(�Z�	Z��|���ҥb/~��_�Zݗ���\;=�Z;����͕��kk۾�}����ۯ�g�m��k���OO���_���5�e��������f���e����v�{^��ˏk�<�����A��\�)x��ߝ<�~��y�K���EU{}��:��+=^������z�l�\Z1�N���C� ]B���%�C
��K�:.*J�[/�*=���ǃS�a�m7;cR.��t.+"�ME� �.4S�ҁ)�^�t:r����tVŢƹ�*7�G��efg�^3{.�"��z�ڡ��p��q�dt'r,�؇��'�~�s����!1-D]�.Fx�����rp�pl���(@�-���\����G�h�ra�E:�J1��2"�HFW����\����$j�\}���	���SD�G@���bE��ĺ�X�(�� F�J��4��Ů*���"��åxI���X)$��	 ~W:���]�Tk
&���R}Tx0l>k���P�`�gT�*O�*Q��^X�d��HFe�$�e��l��U1�����[Ӻ/���
v]�(�(]��bT��aE��tBBR��5����y��_��_,��"ko��vb�#���(
�@�)� 5���Q9;]��:�!4���o	����7�0�R/���[":c�F"��H����������tR�0��RC*��Z0��Z�T8��a^U��)�p�Q
�]E1�$!ņO1�j �BR�2"�c_����0eiʂ&�8�ZE;�c@�X-#�*`�>c��L!��c�-����Y��,���X���K$ٛ�]H�03X"�6RSFR`5D�H1b3Jm�i�L��C�1������Z�������� 36�pJ��Bd�Qو��3VWHޢ��Y�L��@:|H�uᏁQ	C�WU������V�F̼\����X%V�T�h[�� SL�
�����(.���iv�,J�FaX�L�S���C! B�KG葔��ئЫ<�ʁ"w\YJ�K�K��F3�5?=�!�X �%��o�獤D���I�R�/���(�v�gy���H!�= ��J&	p^
�>P��0R0K32�e�$��Yp[PCt�Ec�<z��Z!��Y� �i��n��%-;�i���a�N�,��Yj�\
���"g��n�i$8��j�]�O���R$��B���X%�� ���+���0m7�H��8k����V?��	�L�j5M
gH�����Tj�,!��z��`tȹ/*ś�<M�����[m0)��ň\H�i`H�'&�LZ��E!DF(v�Xl�g� �@���-��%��H��!)@�\,0��XL��*o�!�"�-��?׈�������(�XK��/�B��x�*r�-eDB�x�<��]��V���2�/�%Z`�e2��������'�K^�F�yD����jcɎ���$���`
c��^$�pgQ�(#{cFvS5 f����y�'��b�/*�(<榓�U󒙅�mN��0���o��[�)��`��ԌQ����t�\��JX�Zu�Te�O^��<<cˇ'�"#�`��՜����Ei	b5gzc�")\��E��a��2��!� �7����0� �F�ƌ�RF�\Y{^c�e7-��F��n�;؊�!2{L *B�� 0F>�U^c+��{���`zeT?c^�B�������&[X�����<#� �/ӎ�i�=K*@C��hj�r)�(��,d㡄J��%L���#)�z��R#'*����S�A1��^���g�z����_.Qbk��t#
QI���}�����xӹ�>�����-
F�%�~������M
䣆�����Oz������wE�|�������t|���GNǺ�v����y�+�J��o����������}E�o��$wݧ�_�'���ɗG�����Ǟ��M�Xnz:�>�R��.~��+7Z�R� ��m��C��Ǣ��eQv���]�b�J,�T�X����N)K�A�� D��F�9$��/�"	��f �M˭��`s J*�'�!�^��J� ��
ٳ��$&q0���R;*Kԓ��� �����a���cQ!� V�ʛ:~��2޼y�;����۷=Os��ݻ��ޛo��aB�k���ă�۷�h��
ޗ�2����Z�jG�Y� M��*��E�%�jL��}�rt��?_���r�v�s���z���}���ّ3��;z��������_|�����M�%�Hꕕ����ǒ,ޞ�F]���x��LZo���Ly��'Ww�l�u�{~��F HIђ�dQ����r�R���<H=H���QW._TEX�����eY�- ������w����i����1���7�93s!s�Z%�Px?��,��٫^��N��䨱j���?����L<P��y����i}�i�ATU	3����o��TO��)CT�_R��kM��-CAb���"���r(��*� e�ծ���K��@ܻ��76�n�~����}���KKN���3�w�:���y����S��q{�|r��8w��縚-�
J�#���Oi�۬az}2<���lSh��6q�T�JJ��X#��
� Ux�r4�����S���6r<8�7c�n�P����"A/}&|G@��0�1l�!�������_<>8|�r����g]nF�glz�<�:��Uo�����n�cT҅��ť5�ؼH���p�����[O>y����G�� ���٪�዗N�f�(�4+�rpdS�ة�w7\��ᵽ�P�j��}iG�(�Zݹs��`�)�B����!Ve�c�ۿ�[Ur�Q[�G�r�Wz��k�l#`�9Ë]��/CAb�{��G����[����m���C��%G w�G.HQ�M�������dbc}���������+�>|t���j�x~��7�����g�v�w��3���g9��:<���Ùk�K�s�˅��
�@�s��6v`��f�.���x��j�Ӈ����g��S�K�NqÝ�Jǽ3|p�S#3��t�N	#��ˬ֪�T%�MzS��;�s<4��r7l��z�MḨF��!C͐Lc�8	8M�iZA�a�j�,
C�a���a��6���j��SFH��Ff��C��ꅇ�3[Ú�5�d��mT�L�4��V�a��}/z�v&~ە�}H#`Y;/��z�g�y[W$v�݋���&Gʇ~�M���w���R0G��.T^��<�v.E�6���'l��ո����#T��C"�x1�q���S�"1۳F̼3׀U�Nu�=�R�b��}�e"0���?[Q2��:c֔��c�;z5�/VÑ2�� �����C~qJ�#Cq� �8�0-����!��D/�+�x$3�4z&
��^�E�)Bl�"Q[[��0Y��.rֵ���[%�TH�+�a��w�, V\�?_0�C�	�,A�1��ʠRxJ��Z�X�<[�8?t���C� �	��!%0��٦�5�PM��������� T9�XY �G�0���c�P��b&#$�����-�8�����)���d�����R�04��E`��R.J��oƏD��^3�#��a�)~�dz�i�2,�q
�lA�'s�� ��K�x`c���O�4҄ᔜ2�ɶx̪�h���"_�uo
�����&4�s��!�H��fh�&A1Գ�>Zah4�qd� 	¼�R�)�4ůw�� e=�����<0���}�a�h|�sQT��'�A�WH�i�b�����5�a�L��Q������YQ��0�� 0iD"Sz�(5 ��&�4�37D�>�klf�ð�H�LL�C2��Ӷ�{����>G����z�3��)`B���-+�.�6dR�d�*N�L����Ή'��7�)��K_���E.6����a��h���Vs S��BV4�2�&dHSYM9ZS)���a0�#�� ?���J - + 2[}զQ� ْ	Sm�����&h�+`�l�� �0ׂ��鈞�B)�2�L�4�T��5`�.dzM4��% �8��Ջ�� 	 �f#�7K�'AO_U��q�ӳbB��S�h�dT�EF��'J����؀��* l�FO)*T41μ\�rm)jH��LO��)����ؓ�F��n��'d�'��҇Ĝ�\rJ��D�;��'� Qa�2�� f{�)J�6��Kf��x4�j�\�oJ_�z	�/}`�l�Ė	�Y�҉-�LҧL�I�-fq�1G�r��S�RCH��l
L��4�b�
���i 4S��Ő܆/&�YÉ_�-�V��,M��Qr`(M}^��>+�b �KC�Il��	9��x/S���Rq�m�구L9�
�xO��K�!�%U^S��� Y!�u�(3'&���,w� fH�\�.�EhJ�ɦ$;�Ǥ�3$=�v�֗>��+���Pf��� �&Y~������Q�r�d���+a�F�I2+YࡏS���U�R��l`�2��LM!�Yo�LI ?q�#�ӀM��l�P��i
��*S���]�������k��T�)a(5��b���4��@4Z��� a4$v���>��N���S!I0*��*���Oi�5�aȅ��UC��,aCj���9��w�ţg�Q��w���ne�#sCwH���o��L�?��>��2_f煩a�۟.��綻"n� �)���[�`܅�V�ԸF��#*���O��s�s��?E.�>D;s���tS��ͅ���o�(�O�}���ne��k�]�zn}mm��j��U�������{��έ������a��g����<���~�ϳU����w����?.�*�;{��V��A�O���Ck��8%{l�F<�e2%/�24d$8�O��Bk��)W+L����Ŀ8��5��ÈA?�y���T�2C.���F�,6<��)��﹔y?}i/~J~m����J��l���<[<dVf'B���U���ן~�ӟzMP�<�A<z�Յ���������x��18|~�&�J*�b�t�oH�]�)k
"��e��p�9iya��h�pyfa�������,\[>��������?w� ��8X�����dC�祉
JG^�(��WB��Ϊ9��E�SaiK��t���������?��?x���_�B���.��qd���X�{��'�'�t�mFS�<��w�F%��/�R
f���?s^��)�0$%V�y��������V��]�۷oS�U�͓��Sw�����?��2~|�37�_�v�k��,̬���m�}�>;����+��s�V�t�X���RO#�J�8�X�oq�+Q;���l��NTd�q
Іf��v�Y-��LOP:��7U{C�)�*��o�i�,X	�h�6� ���,E���4=e&z!V�f�ǖ�j�t�|��rxtrv~���W<T������}k���g61�8=�Z���t�.N����������������y?,}<�6�G�xp�����yԛ+K��/>B�z?�}�F�v�[�r��F�8%!��A��e�Ν;J�y'<�@�40lv9= N�u8�C�B*^5 �*��Y�u�h z�!wx[�&pa����*���{O0f=�����<g+�9@z���6<��v�K�͛7�k��C�!�$R`06הbau�����痮_ݘ���̮�4.�l;��{ח{�hV�%������/���=K�9���c�i�M�k�gb��g�/��淶WNW׆s]:�ϔ^��[m��S��I�pt�տ�M�w��6�"?��%��$T�!��X5KPXd-_�2T���`�	�:���Q9H�zVZa@��-�Hj��̱�ML��+�($�H���	\`(C��9�H
��;=C��`QqM��G�>~!_�3�ѕ�/4�z<Rڙl�]_92+ ��YH�<ط0%g(�*�3�:�)%[&�j�I͙N:N"�d��rt�E���c���!G��#΁�
ؒ9�89G�sD)l�l��!6V4\�qɁ����18`%ůB"t�㔾k����;*�`��z�L�(�����,*A��d+2�ƔzJ�C��;���+�j���4>'�j)U3+y!���L�����q�AH�Ʒ
���+��}��ه-�8R1�
��c0`��}P%U�lʥ,B����,6�\��OB>�����0egu����*֐FSC&� ��"S��)=��QF.R2A�����ԋ���f�I���K��PqA�*Y�Vc����G���R�1S�e�e(r�m�x2H�nL�!~r���/ #�3S��	B�Kyů7,�"�,6HC�z�z95�L�F� ?=A����L9bR�s0$��@f��4Ť\h�TI1L PfK?�B9�.2iց�7�k=fS�G���Pݐ�L�������;Y�M�Bƣ�� 9�t4E[�z&Sl��9�U�(k�Ý���N�n�Ta0�d���V��bdz-��0�i���]�fq",��� �j)���R�s�g��!ٙ�If����:��6��ɰ�4J}��@�ǼDU���+)Mk����%��K�N&��@���Y34� 0CJ�3~Sɑ��)�dV�z$z�zx�� ���0f�I��Y�!�Lq�o
�kH���4���j��bƣOI�7�>�M#�<�<����V<f��T��r�b������mK��;�H �+i�z.���� ��洏3 ���V"�b����x�PTiC2ؿ>��tp����'$0[C�����ӻ!~I�9$�4z@vbh7N$L�`�L�K�Ā����ѣ2�m�� ̢bkX�-�a	�c����7sS��\HfM�Y� 8��h �D�?C0C�	�ڦ�Yi�r1��D Ĝ�h�HP��;��T:=+�a"	P�<r09��kz�Z�է�8�SHd��4��rQvz�����Xl0z0$�WT4�O�x�3��' ��`�ţ�1? �0�h4ra�ũ�(��/d�� eM�hXi���ܙ5��rM�NojZn~c3!/�`�ä��\T`�f 6E� �z�2�io��    IDAT!�Y��+a�ԣ����a��!s�em���.9�:�d�I~Ʉ�FC ��E ��Sv��#���c�6e�d�R S���Hh�I1���\zmʋ����I��0�)��0Kp�% OTb�]ۆ�����55qq��5`���$L5���M��UM��W�0�̳j�Y4�NHJ�40S�C٩9=[�J	f���:�3k*=|�ţGH�W0<����ڢdB���5`H�C��F_�l5�v<Y���	�8�j��lɓ��2M���FO�������R�Ԙ<9x��k��O�9��h�+~�.}J��`���x�D ��>�a6[ PN�	LV� 䝹�����
�fM	���ʵ�7^�>��87<�ttv�����gep�%��H��w_y�h���dx���w������nVx��F�zy��wrVI)�Qj�1+�����Sk���U~�k��-��Ι�q|���®^�������~{xQ��-ͯxڡ*^6:r���l���>�����EOe.�������?��#�o���u�9;{n�$D�a���œ�����E�D�nF�֐^y��:O-��p��6-S�z�瘻?�,f9b����n{�sAO�ah�jxdH`�EC�'��=���8���9Cza3��R�27�~��sC��?��?�s玥w{��/�U�Y��B>����L�ш<���WzH���b�T�����hi��ɷ��m�ֺ윇�`V�Ńʪٽ������WԾ�A���1� <YC��)}��M`8��C���a��..�9.ͬ�xQ��٣�7/l�-/�~�ųG�?��Ͻ>3�����ͱ����~����Q��6�Z��ss3�R(8�jxv�$[���=^����J>�X*��)Brq��=Yh���7k(Y{�z��ӟ���Xwb�M$V\H��޺.T7!�a��#�nz(ˋD٭`�% �^lu`h�)e"fo�J�'Av��ǂl:��>������������/��j������K6�C(xK#W �e�/���DF���0�$��>پB�����H��Ԙ�Bn*0���lJ��C��G���P� �H�%=z�����έ��	�%.�"�H����w�aj�l�+D��Vq��w&ϖN�?���ZΞ��ҹ�_C�'O��&=�#���Os�$1��w�b��l�a3���w<8;�Y�=;Z�2s�Ǘ��ҏO�<���[��O���rչ�7n^_^]��Î����'f�'��.cNFr;��a�ٗ��N�^4v�p���V��q�W�W�SdG�%WX=��tG��x4D�_���{6〴�<�p��߾}�2پ�c+;n=	3s`����; ��<E����#~��� v�I�C��ێ�߼}�k(Ƌ'���7�]���7��k�o}���|����ӓ;'{�.d��Y�_�[n�� ����ĩeKe? �Q�N�������y�ڧ���l볗�_�.�x�s8��ѫ�K�8#�E{a�5�x�4z�~���x0��	�Xi��4fs'fkA	C�@�⇴��e'A���< �&r.XaC�A�?&�M���br
��Y�͘�S:�s�G�M
zNYiY��}e
�T2�C��	�����>����0(�S-��@����uZ����J���DoʁY�c�J�}.$��������b�ܕL">"��d�p�p80�O��pS���_W=%[�2�
�!�Ҽ�(�z���sRq*Ύwu3%<�T ���Hlκ�%�.技���9��D���3��P�-w�H�T�����a E�A�0��䋟Sl1��\Ye����8m�B����di�a8���Y�L�����Y�bh�-�v�؜<!J�۬Ԝ��#�2�^
�� |�������R5�c�Y�f5)��0���!��4zTL�1���1k���)�hb~M
li,D~M�-�dK���	A��'�!/4����V���8M����d��xPE�*A����/Z�d�!6�S���Coh
��׬5��V04b(f`CA��H	C���y�@.;���1���,e��|��}��EQ��Ao	���Dk*��� ���4[j��R�C�Oȅ���<R�!}���[ch�@Ӟ���L����+��_��,~}��m��	��v%*�|�0�VzJ$A��!����)}�B����eHЋܰ�(_b@Ӑ���C�!S��m��E����Lh� Yx�7d�G=�F����%��G��PraVOlR�∞�HG���LB�ܡb��!+�l��9������*�\qJ�&r}���˰�&�^àLA�G Ō�Ո�j�8*�)&fy,���B��4Ux�Jiȯ�f̄a1Pr�I�胙R.H-�f۷�V�9��-���J�WJl�� ��"�L�Yӓ�Y2=�4e��K��U����R��r����Q��
,�jE���k<���������� y�0|���ZH%��U�B�1L���4JەgC��i�Y!�,�YS MEb�(�i`��8YO_�mBR�հ���D3�ƊR��/~����!B`��=���i�a���Ҙ�L��&G��)�����a���K���e��f Ρ(�
NT�0q��]5������7-�$������+�YT4y���Y1!�$@�Tz0��fqf2���XI�Ua�g�P�|FL�DN֐h��lQ�7�4YR������.��Y�b��Gj(�����R&G��>��Z��YqNQ2��	�a�	)��([z$�!	�aW���xh�``�g�E1������I���c��Rs��'[r�0��R`eJ+)xS0%K0,6S|��'6����ʤ���������p0U0ʷxȚ)1c0;��=p��{����� G��)�E�!AR��l��TX�DkHbBn�k�p�l�b3l����0r`C4�4B!�ă~ #É� x`� ���:�c���"4;�RKC�Đ@O&�eů��-Z=}�mV�B��4��B�'~C`V`d��5�M�-妐C��'�YHWd�s���2%pT�5�=�^�ي��,=��%dh�!�]7�DBɋ����_�@�|� ~�̞�=U�7�m^�t���y��'g�t���nq��o���@�H�D��^�;T�x���� xG�L%7g�?����p��əF ֋/Oe����������Оs#��E7��,���y^<�����з��-�O���ﮟ>�����??�{n����,w�=J����⅍�ŕŹ��7n\���B��z��_�ۿ����*���M�wW�W����KW.�y�-�`��c>u���K��Q��G�#�jg6��OI�:z���t�0�B�W�v�t���%U�aQ��	CC�TC�����5c"a�A�� �"��Jw��]C��DEo��H�ʳDҶ�x�_�:mSŀ�fv��ל��65�W��XJ!C�j+A�~i�fY�%Z�|���������,0|U���h���������C����;c�^��6��/>�9�x(�&~��л�'��2S��r����L~<з��y��������o��������0����~w�����[X_[�?;x��m!PY�B�2�g4�\�� �8���B8�D(S��ݻ�Q���e����ΰG'8�I�/N��f��U�����z�Rs[�9+�\�ܹ��2��G?���~� 6C���X�[b�[B��3�_��&�o����:��*s_��Ѭ��coHV����K)j+��>���`gmy��Mq��o0|:s}�hnf�Pq���xJ\pF��?����Z�F�C��F�	z�4C9�',h�3�� ��շLE%z&q�b�*L��Ƭ�h�LA*r�	��1k��/����jd�j�Y-g	`L�.0C,�#\�" ��`�7��x���5���@����o^�pV[^X�U��ǲ���j��9�����>���e�ÏО���k�����������������������wVn-�v�����ƹp����|�s����S8)�P��@�K,���T'e;��,�)IHL�L��K�=$M`ǉ
 �e��>�0k7�2�i��Q�Y@v?���=|aSv2�1 �̵K��Co�;�T^"V��8h��+OL%�0p1qY;�XDxV�z����/��@�����͓���>����~���wn-�mә������W��G3Ç�����#_���GP������x�<�n,�����wXKk�Շ	�`p4|8�_�9xq������7����k�{v��V����gő>�b��]1|��)��Pjy�՛5�0h֛���)��@��T�4��Ɣ5-H�H�pJ�3sM�4j	� ��&Z&�,S��0ْ�֐kLl�\���?a��	$62G� Tr��Ɛy~��`���xv����`�иЂ9��fH���y�w�mi�~EŻ� ���x���ЛE�7�#O�\EG U�^jj�q
�'!y1qh�RAA�#� tE1�Б�V�2����\�Br�
�, z��(�	��n�*)~��C��N"ϣ���1-0�d��i��C����F�G�:k�r�"����Dl�0�<Ҡ�h�PF)�� *�J���e��!0[�������PH*l�,��#�����J
������Y�0ʫ�8�B����$���� P�9R=lly��|�	�`شrD� ��0 �h ȑË�h:t�Z��RCUj�	�Ь�PT����DΊ,*� T����cL�)�l�VS�JAoH�-<��Nʦ��y�#�tD����rכ���e��\o�k N5����V1�aQ�ę�>���BRp��b��QRBɅ�$/����4��#׫<٬x�"-�)�I����Y�m�_�>��u4$�@9����_{C<�m����PԤP�����~,�jBSj���c�F��fS�%=�/r��׷�(ɱ�,�xX�ȗc(}�_��J���*zJ$%RѸ.# V���!��|h�!y
��)&�A�d��fy�R�;�y$L�d+<��E#e y� S<�);zC`�M�c�1����x(C�b�M�����l5��X[S��Tj=C����'��X��(�D+�B[nTC����F	�kSʢ5kjJg���	lHKn��(;����%E��B-N��0��Vs*;`���Pr'�764+6�C�Tsuc���`:�h�Gf;d�)k��L�\�d�S?d2��
�l&z��)�LTř��'XQ������1�R�v&�Ŗ�8Y1A��2%w���8�rу���HC&ȶ�d��[$0l�Ii6���Ȣ�f���L���CH4ˣ��� eM�$�7�6[� �� ̖#&�����V) �>P�p�טTY�./4L��!0Z��C�� ���@�#s$�JDP4 01��G����#}�6�\<�0ŀD^4�d)$����`bHF�afBS04B�5fTZY��g'�li�<���]�M��ڰ�a�U���B��Ä���t������Y�i�N��aSFC�Ĝ,�`� ��I�
-��l�"4,<�b&�x���	s����DHY��8�L-�!�}��̤h͢ʊy��Ő�
���|�(�B!��'1�g�A3,�<�M3dnS`��EN�S0� ��I_<�	z���P��S�%�Sƣ/[�H�Z V��#�� ̢"ä�
$9��,d�� -=��	v��V��&wz ҁ�g�G�)B����&XB[�/qT�����m!<��|���;^4S�ZV �a�h��'��  9b5�`֐>%4��0y��  Sy��'wR"�+#`�hsFI��.�d��*]��� DE���]�  �`�Y�g�?L�,C��J�� � lXTz2+���C�L1t�9�4�40S]��0�U�nY���)�[�1�i w' Yq]"C�3~.m��O=���w�[�x��/�]�9�(�r�ocm��<���������5=�{���3�}������v����ڕ�"�w��`>�Q��ݒ��������F����^ڣG�ڹ�x��Nػ��y�η���VW�}1�)[�_|�tue���F�Wv9�,z�#n�e��o�y���w���k<�����~���Ϟ,�6Ĺ��y˷�����?���������s+�3�g'�7޼�r�����G�>����~��;}k��o�;����b�ӣKW.+�{V��ml�?7�x�k�����R
/�i[ l��vw�x��6�	�J��%hݠSpoytda�LkM{�w ��n��2$c�4f[Ȱ=i���j���-�������o�CeK�k�4y����ׯw�`A=j�y� q�-,���Bn��!6U;P���;@�\}�$E�WSL41��=�QXuO������Quk	���o����y�o~�/�=:<>xxogw�{���q�ⅯS>X]���[�޸p���,�������կ���'��O%��CC���v�;,�8GA:�<�0|����A��N���έ_�~�½������s��g�a~iui����׮�y��	�Z4��//�<�5T
�=�s ����U�۷o���������Ql=�w;�)���E�i���ck�PA���[>k-/[�;h�sa��Pzv�SU�6�-��m<���쬈0,�� [qJlR�r����)�얩��!�	��N����B�~ʶ\66�Mo�?��a����wp��4���jw��a�6|6~N�����.r�λP�R��S�V��>=Y�dj�� fS�k�joJ/�S�4zS k��,n;���F��K�Rcf˄F���҉�z�SLUL|���{+ZX%b�b"D�J�Vy�03(+sO��o�]x����|�쁘Rxq^sz������O�~�)�pxT�g6=-�Uφ�F��?;�<�l���ή_L]��d�/������{�������?�z�JE�?q�(l�Zq�e/}ET��w�
۾����2����A�� �TS�1(��ߓH���P�k�g�zH_��L��������,*�{ą��_�E�6�5�dK#~��-���؆w���_�^��L���Ǧ�ݬ���ɑ��������_�^X�yv����|�����/��T���]��f��F��H�������@�kݱ�l8�yx9�d&��8�9r��'O��L`nfok�ɫ/>���?;\�ˇg��ϛ��s�+k�=�,�b����� Q��RC�zHr0�jx� U������*)wCH���䚀!���4E`H���$���8��@?�5�V�ДI�\cn�G/T�����iL �0�©OaB��7_�U`xz�����vZ~�F~)���FG����)g[N<d;S0 z>7m]�=w�;\�:BE�ɋ_N]Hw�������9ά�+
��n�4[ѐ�9��8!E, k�_�]�ˬ\rDE�0#q]�&e�*H�K��* L����z�p$���;���xZVq޿���� �!�3�?�y�Bժ��!��9�SMZ ���= 5�J*5r��KGMD"^4S�i�Z_�IË�#$��ɶH��Y&�(D�0�`���^%Ek�l�C�SJе��S4hi��3�,$���)_f0xّM1�=�ϯ�RJ-Y����J/�6CsJ�V�F���))qZ} 6V���,�6 ��C£��)�BJh��P����e��Y��)���c�mj�2���x�2}0��f��� Zr&0���#��oC�0L ��g2���#����p�@��z���LQ�R�5�ӷ�������1�z
�,�Ƅ&�ߌ3%���X�dE�b"��3rW�\4�osO �o-s 2AC���D�����eE(�ֈ츰dL;�0���E�xIc2����.5CSB�7Ć�!r�z�hM?[ `C�,N0e�·���8ױ��\epʈF�l�6��"G���g�/������"� �Sx48��B�    IDAT��҈ܔPi�1�p
��x���#��у�L��W&��&��%Lyh�6%��Y巡)��)C���% T����f��,$���t L�a�(grI���0�l!���\�@T8�4�k
0L�`
8C�%�Fx l5+�l��&�Rj`yiJ��ll�k��H��UC�81���ly6�'vK�<�Y�hQ�db��Po6z��edV ���J �@���%C��L
9JB���+���8����)!�ge�	�8qpv��IJ=Y�C� ��KJ`hM�
̔�L9��A_��'�bk6s��G�����f��!��?�@�aЪXKCY��M��J�ǐ#�(J$�$C$Y��q!-%Me�ԔF�'+�E1!�R�T��LO���O1$��W��oG�K������ N�,w 8�%ް0dD ����-�0Sy4D��f��|��F�5s�f���������a��+���/�l��/*����r���qfBi��c�^0Hh��@s9Ҙb+�0��/lJ$�ҳM����C1�*�,���2�JO���;����0�3�#k�4!=sxM��7%2��YV`��T���II
�T�����1G�/��;a�����@h�R#�B��EO)��К���Ox��z&�����3?0+���+*�4� zWF��2K�	��Vp��=!=)�*$A2�F���-p�dX� �U=�8�����y1�Ȫf�>G�"���q}l
,��0�FIh�9}AR�5x�H��ae��YSe� 2@Ϳ�-ü���!|r����V$�Z<l��g�����&7D�!r��1A�a��̇�ƃW��`�����hb�4$빳�Z�`�ʑ�1ԃIĩ�Y��f��x�i21d��$��&!aPj����d��)۟Y10܇d$f�
�EEIփuZ�㑣o�R��*<�.������s���r��O�� p����O�W��Y�v���Zם�m߬:�������J���������.�u�Lm@��[1�';�{V/��T�_�f_ÿ��g�<����ݿq��������;/^m=yuzp���"}�������o�v�����l���/?���[��}����k7����.��S�Տ�vNN�O�_�5��ã������;������ҫݙ�����Ǘ/�=�X������Ϗ�w�_<<��z��㷮�]���l����ӭ��[�N��j��>;�/^|��ŗ[w�?���ko�z����K��'�H�o����Q��ӣ��/�^����~u�����׮��̮��fK�	�?�����������ɖgW�Z����)a�m �5~Q������˱%f�ʲ���z�.8�S͜?�ûÄ	��+W �h���;�NT0!_n۽�޷����5TV�3��D��m+��l3<x���+wAo߾-�n�I��?����&��l�ۢ���H���#Ѿ���
�tneyo	�O��|k��,�{�?���|�s.��?y��ٓW���m7�.]�tq�{�|��O��}���W�8��e�M`�)�;�d�u<z4`�_Ou�=[#�gT���6=D}����������_n��嫽���g[��V���6)
%)����f�h�vx�KJ��'�Y���Z�j.N�U"1��H�=U�t~���"�Z7o�D{��]�ܺT|������!%+�N<H�ۊ���O~b+��`�������;�����5u�Ӛz�))�
��R��>�N#�+���_��_��9�{�b���̼G<�����q���|��Eq�ݛK˳�8��x�"�1��	j8#�	�n���]^�O>��$ȣE��UOk���Lj�"����4J�>��&BH&a�V�E�DM�����L;���E�/C�JO��w�<ҳ��QP�*I��"CBS	<�FBC&��7k?��$�#�������g�?ټ4�Iڙ'�kެ��[����ea���t��ħ�A;	X��g~�o0���3s�<xvꫫ�w/��έ�-��̬�:�z��ן?{�����1��¹���+ގ�H4�-�HS�N��m'r˾��4Y�=��9:�\�ؠz[J����Dͪ������0X��%B��}l��vmkC�h��J*B �吀������8���v��bm�cg+я��b-������汇�s+˫s�7�\�~�λ?����\��qnvk�C��mWPW<���r�t���ȯR{�ii��=�۹E'i+�Ӕ�E_?^�p��9;�=�B��'[�o=9{��7V�7�N���!51k����e[��+r;�@iV#��4�V��f�2��ŰWi�҄	?���
�c/�a���������_<�k�B�|V.�L1L��H�f�ZzC C����;�`0ˎ @��@
 C$��EB�y���ƅcDj�����m0��/����I���裏d��1�2���B�R����nW =|�_ �2���`V�/Iy����0ԋ�C@!�!�h�}D@N̲c+SƔP��˪��
9��g��r����O�?��\%�V��q��N�.�̱�[8�7��+���T"�H"�
 Sr�/1()ך�S
�9%rC鋄RRzWz'eG�M�`��D�� �r[Aũ�r��uW/�B%���Ʃ�C+YT8��\�����i��3g9�Ί��ӑo��q��Ԙt�&��F�dx���P�G_�A ���ȅ��t�S���9@+n�����`���QxJ��Yz��3�4}��"�&S=sS�U1g�hfy��7�5�)�V9wrɄ	C��@Vfi����\���,
)G)�(�V%CzT90��,	� LT���)Z�M��V�	Svf�S$�01�@��%r�De
xj���Qh���J�MA�A�Iy�)TJ����Cã��S��C3�ա�Oc*��b`�u$N���i�1U(���o��1�:e�x�0��"sG�ߔ�C�S��"�"�r)�8җ#�̝6U'���`�o�Qf����CV��z���`PjCV�4Kl�2Sl�k	�d�bҳ��r�kfs
�*t(A���UL�	�&6�0`�h�$N��95�)�2�ӛ%���!Aϯ)x-�<BN5*�!�m C���	rJK�P3d�T�"%�>U�k���I�!+���- `���Cȗ^&�`�����D�ŀ*f K@� ��)E!�.u�f�5��9_L ˎ�t����O��'���BN�?�\�wP�RJ�#Tv`Q�]k��^�P�4������
_���B����� F�P�Q1Ә ��H��4HD��>�' C� ܱ͜�GHJ��hŜ��Gʬ��@h;`(KA��eE_�y�,��Li	4E��D�cH��'Fv#�p��;M`����!|��2d�_�1�2W���dIER0��%��>�[V=��91s߰��y��p��ѫ�d�U`�D�S�>&�4����* g!��,~���/M�dH�bf�J`J]�NM4�	[2<Ac+�b��GH�7��F�4�d�|��8�DU 䊣gB϶���LS�0��P��" &*Z���	 �a�` ��i֐��f�dSH4C�l�1�k
�k &���)-f=C���ya^x�cЪa��I[^�)NCl`y)BC��&����V+l}��3 ;gZ -_ �"�� W1���)0_��W&�Sv�yd�������4������B�����7�����P�/�����"�l�^��"��Q��'0�c��F_�`h�D�d����;d<iAra��*_����1�l0z 2w�6 A�\����	��|�i���9�`y�4���J_<�����1���8XN��L�m6�"�nZqH�\�E�_HS�YSN���a�d�Ac����,JD�M�HۛҔb�5N�`cvd�#��f��:�:VeG��Dk��3��!'�J� �x��Y�d ��$��t��d_�X�v��8
��r�Ǐ�eH�aY:��_��������/�}�`}ue��ox�sqmiy]A��#��!qa���\�t��non���"^�[^pW�w�͝�,/��//�s�����z�7o�s��K�/�R��I��t���[W.]9����?������l���k朻��3�ǻ>оz����o^���w._9�k=�t;������ֶz���7KpxCŦ�_�9~q��b�ŧkKg��z���5?V7����G;�{��G��|�xN ����89tc�`�^��H�9�[�Jmo�6~��o�;�}�uqc���w�nm�z�W�{���ض!�2[����w��X�U{X���P-�e�+�󡗔)�Twȝl��<���6�&2���~��Ex����_�Ce�*�bW���e��u�����w�^�rI�����-k�k�y��5<<Z��/���?�Ƈ}h3P�7��۷�jWx�鷿�W0J�)_���A�ҷi��Jͭ<���[�b�]���է�|���ϝ��vu�ו������:������񃇟�����G;�'/�|��|i��S�k+������0�C8Α��4<u��7mݨ��K�1�D�bx����������0�E"$J�x��Q����Y��dnq��ao�-��v�������+��+������o�|�����˫׮{�RU?~����H\�I���[t�������+�ݢ��,�J�Yu�ޅ{�ꩀ�`�&!6w)��\-~�Tg&6�����������/=���e��m�N`Y�MqFƩ�Z&��!�|�����m�9B�G%�}S�ƀ��1H�96�y�/0TH�@�S���W��F�G'ǯ�q������K��_[8�.����e������P+/���_�b),��b"i����.�����5ÖU/_��`L5+���mJ�a�G[��|))����Bh�v��*8ccpk�T$��ʪѨXŷn�/�.`��P�E�^�%z�0$畆�czM��8#�������Z��T�T���������Xٸ��qvp6��0�����e?b:�������O.ʟ���̞9IX�u�wz4?�|�������E��}D_Z8�����畓���g/w�m�����T,�p.����h�o����匩n�8�)���r6:<�	�`s`� �6��:Z�0��*��
̗�i˪3=�ho�xlP���T�Qs�	C�fOs
��*��m�ǀ�#��p8���Cf�|��m��}��|GÓ�}_Dp��Ņ�������߾�b��F�/v^���'��H�xp�>>;Z���3���X�`��zb����}��GóQ�q�w9����߱=����?}�p��ɕ�����eko��=�F',ⷝ�-����G#kCE�a������@`�9��rGf6���p`Le2�S掭0���> 0�����(i$�!��a���*r[�>+�YPGn����"�La��ԋA_�`H��1�ܶ��P�0aho�$��f�����5G̃�'`�7ǂ��%�3�����=��{�]W�q7|��hr��nW;O�������x�*��ʣ�e>����2@���Ѻċhyq*�Eh�����Y��e�w�1�ܬ\�xW(W� ��W�G�l�޽�\4�U�+ �����.f*9���I�?�9��:Zq�V��eK`�VB*G��5S��x�6S
�Д9Z������Z�c~~Y�8����j��-+B�����U[0�ȭ~~]ڑ0ѫA_�Q坊Uå�ǣ��1!}{�l��#�ȝK9"g.��_���ѩǊ���6l7��2�^��44E�p�I��`d}Tl���Q�ԘS�3�4�04zM�8!N������&�G��`�����)�)/������)��L����f���*F��X�Eۮ#���00�j��zT��͚�b�DT�	LY����;<�[����, h2+SͶ���y�����FoJ�#ZH�2G`���4��w
�);�GB��T
VH�USFi
3~z����1t`:,�0s�# #�z��y2_4d0=��ѓM�]�� �Y���1c@��n�E���\")c�)0S�BV�(���1�E�ɯ ��Q���\�]J�2	��8-*2�«!����C�dD��Ȧ0�*`�b.�ȋ֔�Ka�n��CO��(Y�����S��3+��1[��D�h�L) ���/�{Ō�UF+G��`���D��DZ�@(�b��E�������Ȑ5��Y�h!cN ��'$s�֔C	X��V�H&0s�<f�!E�5�04)�	��V(� ���
�3���3NVe-�0�B0�4�Qi�&K�eZ���
ȗ/d)�� D��g.��Sc�7��&�4�`(+#��@O��4e�/S��)���y!���d�|�� IN���V�T�1����lcTzJ�	!*����U��I���wS}��-w�3C$Ӕ�0/mWz�����坌���!eTy3%0�RoV��
3�)aW�f8��:��;`	�dV� ��Ԑ/2ap0V?�Li�aB���P�ِS�Р��j�0K�9A?��Gh�j�E;4�( �t��{!��)�jŖ�^��B�sDc���̚�.�`�@c"#)�WͲ�s��?� ɐ�
�L`�)+�`l1�N	# `z2=Al��jL�eW��T C=��B
>�8��1��g�MI3�)$	f�k��	x�^^f�`�vN+!p�H *=%N�|2��	C���J,��r�<L$����@3L��B�8�Y� �=� �Fx�w�Y�8��&����⁤�N��*8s���UC�H�Dȩ��a�1����\�*��9����֛B-Yݚ ��T�� ��iF��I@�>Q��B�#�ƅ�xp�!�+I `f==/Z���G�$M�����\�G�g�/[�`"���,[�\�BH6kX��+fH&����pM/�؍���J\<���#�G�5Ҟ!$�"|����9���Wt�)wz��K��o�'f}��9�����f(#J�'���1��*�ri�ţ8!Eȶx�A.�@"2u��� x��!����P�t����'�|������X^[�2�;�{��/���=�y�������^���n����d��u�_�t��ga���Ά��<r�8�KI��{�K�s7^�znc�_͙��k'�?��\�ܕk� mim��b���;ݍu��p��$d^�v�S�O?�b��D��[�7���.{�O���gk�q�b��\_Ey:|u��CVN斶^�8����������ř���Ӆy�$��l��5l'���N._ؼ����x���98߫�O��o��`e�����W��������}��;~}ӗ��UΥ����U�Ɯϯ̝�y��ōe7=V>��Ͽ�.VVd�E	�۷o{��w��|��N�"RVv�@�p�Cy�n{�81��h���E⹦����Μ+��8����Trc��qO:v�O.�-Uco-��A�㳭g�yWZ�I}ծ�|���;���=�po����;s��:\i4�j�&��}����!��7{��҉Jx�s���������2o�9(l�����/�����f���&ݳ��tɒy���9�e�lo^��vzp�psygo���lu}�oS��� 70Of�|��%'��k)���O�cT��������_�S|gu��O;�����iLY����W�x����?��o����ϟ�.���g��O�~���@�^�Z����u+խE�]1��Ŧ�O�5`������=V���~�W%���a�z�KnKb��ݻG��Ν;�&߽{�o��o,+��/sQ���S���w$�&��Mi�~�!�7n8�}�S��ⱦ3���&�6l��-a��ih��Z������t�}g��e5�������g�V�<���������N��#�wO}�����CM�w��A��븯]w|��x�����W��b64E�xJ���D"i����pܨ���T�)-w��ʺ �w|��ϑ�ݱV�YQ��Lc�!X8�V@��Pv��ؑ��T8fP�އ�����1R�@9(1���o�I9Tl��D��X���hԲ    IDAT-���������=[�H��h�}�" .�xɆ#��_O/�x�铮�Ϟ����=:9�9�Y���z㟖���N���ś����G��X9}����?�9��lߍ�	�W��2>�䡝�Nֻ�;��}�#qR��9�U�^���:*:�։�.t�I�����*9���@�Qٚ�:�lk��SY�-���``�����{�2�9���;��ǌ`85�8���e��9�i�7��_y�?'�������̣�{~-sa��;?���k�sȳ��E��=s<uJ�Qr����#���dG������OS�M���q�_��n.Z�ӳ!�9�g}ڰ�'GW�����Y��:p��]q�;�3 fE�$%Ҷ�-E(�����[�I��!}bH��-�ɢMQ$���ݷ��~�^L	�D�ɓ�y�ɓ�U�U��K?M�q�̸��\���4��'�Ԗ�!g��(��-ej��	%�E�E	�����zF�7�X�U��xa�3]�Gn�u�R���0! �QW��2����8a�iࣁφ�#1�']�&0�
^$M$��[1h"OM�ŻN!)�4$
V�}��a��;����w�}��o�X�V���=�ڑ�f7)\*����`�=	ﴤ�6�`+���l1g8u����&VB�}��� ��}��kP���s�_Fmth5�V�Dm2it�[!#r��xl[�`5E%x�rb���4����ɰ�KQ����e�[	�B��6Q��F$�bk#g%T9A�P��z��qကĹ,3˯���y��ԉP
Y���2�P `�Id�7.A�O<�&@~ �90�@��~�#`���@���Y!����[�)��0A%�'H���b�"?jI��D`��0��՘�C�"��YM��BOVpbc�h��fNCO�X��tЈ����^3A�l�Sǩ�kfCO��fFT��E��'�5L`$�.�� ^ovz�=�Ŋ������՘��#G�� �(�
�����
0li��"��?+�Z| o�)��Ԯ��/�4�Y��\����#  �EH��(-���BN�Z?h�GŜ@���dU���0⚞ B��u΋��(*J*�]o-�ER]�<MBbB��Q�^1��cìWM�[�&�`&�������0< <��ũ�>^(y�į&��iNÜxb"{��ҫ�Y3� ��%�aK��W3�E� "E�]��3�N��Њ�� �$�d�`����f}&%��z�`10g&��eل<&�'*����6M]<��,BEH��V5s��P�[H�\ӹ�!�SN��e+�C�wk�4� ��w4�h �!�R���3G  Q�MS0����		'=�����	�ϔƢ�%��.�G}�bC�
 ^Rk�+м�G�+60��Cn�;1��S3cgΖ�ѫ���̋"xu�	9%*HN�/ 0z��85a��ؔ � LJq*�`
=*cQ�T3Q���%w�M��nƅ��	�`�9bZlѨM����l��X��p VxĖoU����8٪�d|���.E�&��0�� �0�3�P�3:MV ���ig����(+']e&1�e6�Hȶ<C� dl ��#��R�>)b��I=d�C`.D��k�Ɛ@/ �`��^ �		�l a�-0��҅D��d�xPS��c� �A';� �Gb2NC��80T�R� ��k��Y����#3��G]S�
��!���NW����!�q���ER�L����I����J������|�.Ny�8ϐa��,����	Y-����Bf�7��T4���F w"r]4�&�b�a=��Y�t1�|��$���@�CS�0��J�?�hqe�d��H@E�N���\ ���HI/�
C�lUpF) Ne�F�1��)x�x�n��C��w��}�,W�������؅d�h"�e��*����Hh2jV�b�?�ԅA�4��: ]V#*5�f���Gc�`���;�2XxbV�Ȱ���	/�.��e8����-�H�̑��� ,-`b�I��_������ ���<0�Ph���x2��*�3��#A/0A[M����i����Lb<��*0$��vJH�D�d
����(9�G�����I	/��Y)4>�C�d9�g�G ���Db��d�ǅZ��H�dH�xT� *eF�6�z)��D�Ʀd
�یNF�<.�i�%�o>>9w������YL0(c�Ӄ'���������dv�ӣ���b<�wF���`�;�u�Lb��]�>�_���i�����G_��|�xk������jG�u��mtʓㅟR[�ĵ)��l��F�c�#������������Ӌ��6�+ݲ���7/��Ӗ�yt4�B��Wق��|�r���nw��g�������֔g�7o��}p�յ�o-7���n����;ۗ��lz6��
���yNo�Y�ݍ۰�A���u���ɸ�y~zҚ�G���`��GE����/q.�������O�~��ܩW�����x��|��W��~�s������^�Ƌ7�+wE^�O�6g��b�Dݚ����\H6M>�;��yAc��`w��U��ݪ��QUf|S���=�!L�ec�04����o�%�͛W��V��F񛩞��N��W^���ý��qrY��t�w�<eh��s��f����O�J�=�u��t^<z�իד���2���?����fܽsx���չX�ֶ��u�q)��j%�$��rW�<?0u����y˃���w{��_���X���"˦?��}e��M�b�?k�O`fG������ɛ盓7GO�c�F��oy�������Z��kh���a��r|,�����{���}�n�O�/��<���Ϻo^O/�}��W�خ�(�5Z��g�_��Wd1��.�,GH��LBc���c�RN�װ�Kw�ړ�ů~���@뭑���/�[{�,����_w{m?��N/ՙq���S� �;4���]��k��"q0�1�nb⛂��A`N.�0�S'}75�|,A"lw[4��|>Dhs�K�u��c�3�:��	����5M�`���Ç.����JṰ�/CQ9�s��q�\����L/f�Ծ_�s&��F��"�����G?p��'�c÷�����L/nK=��������ܹSn�_v.=�11�=_�;��}S���nY���I��W)i��2j�!(�i���S����,�^�EER[�+�0!1M�g�Rgt�%Ա��!@�Q��9I�8&kv\�6sp���A&^�uXF����j�p���8����9�Ƅ>M�0����r1?��_ݙ����3D{�>���ۚ%S%��H[�J��BY�V�:Փ�����r��3�����V�;*��n��k�����/�N	�Ʋ��@���{{;�����/�y�����<gQ�����Y���K��Y��*�ִ�@�}��W_}���5F��fS�n���$�>��oݺ%�4���%�;�rh�
��r��6�li�^���\]��&=A-*�!�Hp��ѩ�U�X�l�|���=��`g��k�G�����~�GrG������zz���k�O\��a���rN�l-KS`��om6-��qV�!�r,�On:�����v&�x7��뗓��y۟����QV��P�,.�dJuӡ�, YxU<o��ޕ)�3]��f�^�R̶}��8�'?x2<!VH��ƦI�W�p"y�K�U&&��Q�� o��`P���B�t�J�|)�̙���d��yDn�́�k�#�7�!(L���lQeDl�
�0 �^�Ġ�k�`��R�eԢBh�(Fd)�A���#f��!`<�'��1m���>�u����	L�+���a���������u�1
�~��٤����_�8ǐqV�{����8�^rİ>�#4|a�#D�/�h߸��D���*{V<0�6Z�����ַ��tF���B��;_d;��q�r3%xxp'T�j]1����-�{��9�hJ���_�$�Ƽ@2w�B�)���5a�s���w��8,�ĀP/�oh)��>�L�x�2�2�5��+b�,��L�o��Z~d�FΓv�	LК���S`&�$0�2� �Oɣ t)� �*M�1�a��@ҤЛ�g���0F�T�s�Ef�l��i?�&s9�m�hR��H1|0���_� H$��h��
&M5�4�׋
�.�dOxd�[!���	���99a���*���f�4Q�k�቞�$SL6��c���%�^���QM�_re�h&��C�~zɤI��or��\��@���!��\cY���i2Q8�x!�E�cEI���w�&*����g�_�T���U�D�M"�X��I�ԡ�@�3�K��� OCx��
A�����[���
s%zM`���-9�f40<�B6�
*y�w<�4�`��&< q��L��#�H�)B�W�MAH0�lx`����O�-T6)�`)!����	AΕ�BM�P�Jf�d�����#RzY��Z<���k� D ���Nq�'$H5Yؘ!s�
�Z3.�04�dh�V���K���AAk ٪�
[��LL`�<a�h*�xI01�J��/�FA�d�t/�-G���,i�O�Dmh� J	��5�˿Ŝ2��7Jx4H3d�FaiD�f b �I �Z5CzV�&9Y"�bD���)l�9�$��ɡ����R��-��L0����`�
���|�I6�` �F�8�|6�QM3�Z0*��o�������Or��/�%*��.J `cd��ģP�[I/$���X�Q�2����D($]䄤	�6�R�͸�Z<��`�aBRj�?C�(����$  ԛ�eP1Q"�Rbet������D��k�^c$�4zQ�u�3�(��-M3Rq�II6��Ӧ��H�aaH/[�{ ��S�q� `PF�UM�-�m��:.D��5��,6�:L�����0����)i�!c�{�ZS@�&M�B�<�8՜�+ɧfz��������0�A2#���ĐI�	_�����6THb�Q�ѕѱ���&0�ؐ3$�5�C%���tdi�@�`5a"��:� `���P�f0�2?�"00%'�)�&Gs_͘[f��6kI/�!c�� �KH�41�Uh` �㫇�L��G��1͡�z��Y��Q#�4��O/�%����w[K�	*x���ģ&`�c5�X�[*�t��4T�����`ScC�YL3`-�`�!R�z�GzM�
s %�4MAK$���b_��P>ي�6g%��'�� )d0J��L�?�	X�0J��+�jx�0W*u9��襉������;RW��pM��2����k%�y�@\d8�N�Yq�S�-�K�Ux|AP���1�yP�����3j��5s<I5�PK��?�b�@		oh�7kJ�
&�'�S�z�g b�
�4a�*0�	��Jb�$몛$`,�z�`³��߿�,H����w�'㽱i�l-&��{��"^�g�Io�q#`k�����V{��/�Z�����/���֣�����捫��������t|��-0w=)g�O�=A7�-'s�Ӛ��{A�Y��UPo�t�qv~��/,Ƕ[v^Bk��Z�����nv���M�7�����n.6��妥�s�r��w�[�o^�����i��]�/��ӓI���jܜc:��o�޾���+�]5Nu���rnj^�X1;+�H��q���l~��d:[���g἟����vv;݁k���ۿ�?�y�r����	Mw�����E�-*��6�V���F��7��;����/&�`<���i�z�Ѯ=;����vۻ{�;{ۍrɹ�]v6�w?�?��#�� �:^P&��k3��r5�[aLݮ�C�x��s7�������o�7���ꦦ5�O��~u|�j��.֋�'}V��;��W�����ټ���lq���^����h��ǒ���kM�jw鸶,��`��o�r��ͫ������u��*W�������gLMw��C�$���Z�qeޕx7_���AUKn��k���_xB�7ض��I3\�[�n�������xp���=���������Y���9_�����/��Gw�����+������U����Nf叕mLyP��c��V,�ň����S�ǋ}֘M�Yg����������k�tK�;l߻��;�������Csg��Y�jU8)8��>|�~$f�����'� z�����S�h����n�^�q�dG!Q9�2�l�]�t5U��^rApv��L�Eӑ�ٙ x/��!�xy�w1�����?��c�n�<~����ݻ_|�F?����	=��K�ly's'qa8 Z����cr]���Y�$��h{b���d��³���������~�q��5/�޻:�[�^�;]�/VSo�-�X���D8�����0L_�Q���/q�CѕD��k&`�����bF����2�M2A8i����=^l�D"3���bHW��<yR�LZͱ��Xc��F�{u��#~�M���f��d5�rQBnc�/&��G o���1Ņ��	V�W������'��[?��.��`�;|c'�t=�,�I{6���{���l�������?��;�;�g��ngy0�7�;`�Ӡ3�W_=t�t������ȅ����<>=8VJ��Y�`7o�4
�ܨ��M�M��ѣ�ϟ��`S�S�\3�����:�U~���{R��̵bR���m�F`�����v��t�G��q/���-zLȆf
`�# ��h�f������{w?u;u2?o��\�:;��}��>����r��tvt�X��eʪ,��w!�3�VK���uY�,9З3�_?5a�r�X6�20�&Κ�9�T56�����tt�j�5�ӥ{��A�m��Zʲ!�0W���k���I%AR�L��*�@���U�R� �c����jz�L� 
!z��5�*J�7� �K�8���n�Bfe�����ʆbB	�$��N����!/ ���5I�/ �H�r¬�fB�6�j�8���fQ�S�>�0��O(u	[�<Z��5L�Jm)���8`����%�_0\[��(�3�5ﮘ�U��5O4H�	��9[����m�pQ���͐w{�#��x�W�#���s�e��=3�v�	��ͩQ*�`�pmP��	���"a'*zC�)v����.y0L1���+���2�?��?3R�N�{+//R�ȃH�D�C+`T��_I���v2��J&��Fi�D��ܡBN�駟:�8�(b3.<�6|�f��rNϑ�J���0�ƴ�x��H�����X1$�`b�TW�
22%����)����a�3��a� r��G0� 4�Ћ����ᎀ!�u(rm�.`�5|l�x�9��J%��#ȬyJ��#l���(�za��RFD��`�^B��IPh�`	A�`�����OT�t��L�C���2�����rzՔ&����Z'��L@�Y�9%�^͵�Đ���l��Ŧ,ESH
+1hJ{� 52a�e!a�=���.�![�QC}�rX*��u3Hl���!~E�xw���nUg]Y�<
��߸�GH�\��35�^���3�`�0Ŭ* 4��'�̚!$`~it	2r�4�"�Ӂ��.��C
[M�����@�įZ0� a2@J�`��4J@0��!�LA/wa�U �9.q�WG��h�	�a��� P׆5N�[ �F�a�)�C�^�h��S ��rB���`�j$��!9�@�a�<ZH��T�*[���<�QP�ѓY�$f��Ix!��4��$����Vf�����i�bS�'1@�d\!����p0�c���)��HـL��5z5�Cap�D�������
���<fʘ�s
�&+<�L21�F%�
�:czCK�&C��Iq�>#�e%�� b�VP��E�Ar�P� ���[�<���@���̵b\4!��Ո�^``���^� yK0�<	&x�.�� Q1���M<I�`���5���%0�*��b-w�4�u4QEF�l�u�Q��;C�Yc`�� �k����<xzzT��EC�Rl�N�fb��!�t�cK/_��	�
�PG��%V�BŶ��^M@L���N    IDAT2<��a&)���Q�0NsDV!/��^�,��	�u��'Oz�}�������.��$�#C�x'(��#����'KƘ"+�����Za�wH�&0�I���:2}	fE$Z] ���𛘓C��9���f�����9��%BMr��٪��`��0��1�t�b"��$B[XoE�6�0�ի�G *�%N�h����"HM�0���/�� � P1IT��=%wLdLԨ�:� ����<l�b��̊�7'�XQ��iN�������`�oI��� %u`�lE�I"�-��3�^'_�2)��Q�&���4�0��D0I��D����h�{:YJ3@$z��)8	j0u�1R�\8\HH>���Tf\����f~&�4���:	lɹ�e��I��&~�3%ל&�!�$����$����0I���ԓ�'�+��ul�1��.����EB����9�F�T�yJ�B|�V�l0�K�<0
�V��Ê� ���v� /0� &AW�4%�oN
��SBl��G+��+�`�ux`D<0C��V'Z5%z�/$$�%`�`��P�ٰiB& T偞k���GD3"��g՞�����K[�Ak����~�=�n��ys�F�I��A���l|6�F�+ׯ���ZO������E�����#;����ܫZ;���ٞ�Is<yy�����;��b����2pi�o�� WIG��'v^,���ތ���5�9�U���})Ao��ks���sGѝ��>G�Ng��s��2�< �w;�U���ɫ��t�q��� 2@Ϳ_s�ק�1���{n*Y�տ2��Fυ�f߅�A����?�*����g�Mv=��n���X�v���:��b�����+Wo�Z�[���/��b,�A��ځ7���ag��Kk�]o���������R܊�����ϳ2J"�E⾬c�h|Bp�"dߙhz�'�墜;����=S��Z�{��(.��6�$��wmˋ��x9������{����-oٝ�{3��8ݴ>����+^3�pq8��G�=�\y�]��^y��[�N�N���k饠/�:����M�ݽ��z��-���tm�:����d�Pѕ}Tk9AKª<��G�hʹ{]�6��.˽Q�u����_����|��U�	�Y�]�n{6�v7	h�Q9��s�ޛlכ�?��7�,�ak��h�^�_���^L�_�8|������O��l�uC�m^��9��0Y��NP���#��U^=�ֽ$sm����xr�7����^w������|�{��[�������#���˦3�:��˧8�u��u]g�U�s����`�>}��rZ��$Mx>7� ��N�\Ծ��i�!4@kC�a��q�r���~�����,"���߻/��ѣ'O� ���`�����GX�#q�S�a
�R���Ļ0$�%Mx?���I&?��s�r�TӍR�D�=������|�;�ܻ˵����_��Uw��@p9ј$#2RE�
!�DƩ��DE����6��0L�Lq2XE���w��0�����d3B	C&(`d����DK��s�`��"�΃6��KH9��cs�Tb,u���Kφ2gb�1$J5 ��L�8	�Y����D}��4��b:����Mo��m~@��W���~��c]�/)K�S�C�_V���˱U���+O���~��N��F�;�?�kW���7��W�����b�f��ׯ�����[�e�G��F�5�)��䞰��_X�����oV�"	��ݓ]� �����U�##����ҔXɔ�$���/�o���9`N1�fj�����8m!��aF3wj���1[�a�'f���w�-���P��I{gx����=��w���Ã��~t�ÛF�^?\��X�Z���s�������ѪL�=ʷ��L��W5Meu���|�(�eїW�:0o�݆'��oZ'����sʯvvfn�V��cCE�X4�1)��kB�hƤ�e�}R	>xz%M�c%c���kuL��kfʒa��eK���	�=�F��2�j�5�Q)�`�
^���b"	�gZtQf�b���xdC]�l<ڀjEW�&*��R�)-3&	ɨ���\�<&ڄAFh�	�/�������w�u ���I��@�+�tq�_�ӌ���v�zmC��};g��C�x�ɨ������Bf���MS�v�$�؛��BPl@l��!C�_� 7
a@f)��4�Ċ]�a��J/lc��%�R�����y'�ŅMj�bv��4)����|��1|~�Ĩ��"��w*u�6�|A��%�����Ǉ���cdk1I�0b6@����1А��R1���C$&�(�B����  -���̅`p:�� �ua̑^×��j�C�X��0�	�.ME��w��'���4����`��J�4L��K~�Rs!�j]f��5<���������5�R��X$��xͺ�Ǚ8��)�BE�IR�)<j�"0����M�a3��l	L �d^�x �CHTjx���ۋP�� S b�8�Jҥ� �hf욡�a��,K@��ĠK0NJ 2+ӧ�Th&Z���B�� �Ta`�D z!�PY�
,&|�"И\Bb��Gtq��E���Ze�Ҷ�ab ��M��Ge��$;7&l3G�̑h��꬗���������0�Z�L/f ]��AH�"��fMK�<y`�3}"I�h9�Ǔ�dlQC�\�8�������LPi&Zxl9L�J�axtq�`2R�R����R�ߡ�\Y�� ��	��F�Du�ӰJcd��&����ڐL�\�@������6cLx�^�;I�=k	����g��   �dE[T�j^R@�^���fʱ]>Td<�P�'d���� ����KHH0u&��R!�c�:��*�U+� ���������	�5B��4�1�{�9��$�-6q�!3F��BT\�RK>H��)A���&��&-��2L�.x�	��C��x��;z�ir�P";��M������P!É	6J���S�p�`�T�$p2�e���"�Λ��i��,6��8�ă������G��q�D��8� $�%�jjb�R�����5�QhZ��ؒ@&
dL�P{�V���E�q!ZTH�%�"S�d��^��Q�F2�$�$G�,�� 4
�h1G�	,���2@s5Cs�+)�����ŋ��84�ECF�d�zu�.���G\>4�z+]� =+~-�����,T �Q�Ya�K���;���BF@A���_3�52��[B�f�	�3��@� �J2�9E��KbH� `�������b�1M dC�P�WC�
y��
f+�@)B5$�B� 0�Usd��Ψ�H]	;�D� �N����	F	�0$�x`�� �
 YnI�4Ȱ� (�adL!���#�k&T�� )����'���/C]�a��L��RM�k��Uԧ�|厜],��5�\ aN� آJѫ�S���Е1
�/0t�	3<*� E��̜!_;(3˝1f
'����Ml�3/>���k�H�&��	�ƨp��#J�I�|A$
�0B�9Z`�'�b��$�H�0ܱ�N��[Vzx]���RDȖS�Z4yįi^X�A�B�f��h�L���#|����Y�h`Ԭ`$!+0��D.Z�Њ-2f^�h�1׌<x���TJ�ߜ�!i�I.�`�$h�7�P'�8%�����W��2�L
[��"�4�B�xؒ@B� z��f�K a���H�/[�pR*a@��� w�P��#!���L�#w��<�z3X��\xe6q�nk�s���F��������'g�O�$v�����Y��]7���9խ���t��*hϓ��Fg�'-g���|}~v����ʻ��;��<�LǥĖ��`4,�B��a�H���2R��yl���f���5�X����Sx��t���ρ����&������}�7{��a�O�B�ى&�_.O������vf�G[|�*?7���.���\Y���v=w���	��߻z�=ou-W�;�B�[�m��]�z��i^^9�x�`��^7�ư��t�w酴���'�����#��2�"�V�ZEaȗ�2�n-^.W��;݃�Nwom�d�����Ϩ`���f�pa�͵MAp�ZJ�,�^��ެw{�����ce�^�|���W[��^kw=}oȊr�{�^l�3m��;�?��^y��$ݙs{���o�Ζ����Vw��r��`��ꌼ��Ko}++�oO�)���r.��[�R�"�z^��u?éر��أD^*fw%��u�r��@�+����Õ�!��Q�F^�e�v��U7��nTK��V{����+��;��gnj��/._˴y�������p�=vz�b:9?�\o���`���l1� ��t<y�ҙ���A�]?0��$�ռj�݆�J�oP
_4�pْ�d>w����g��[��������?�����j�9��/&>,/�����d�l�'i�q�+�����#�>tM�����!ȁ�RsT����g��d�z��4\+fh��(%����b�"F+Jae, .�������tS��Y���'�x����/~�<�)g7�����?u����\�u
@�@�6'~ώvd�'ٜw�@:��<{�sN[.z{��aZ����b�f�����[�y��j��Iz|�8�^�WM�9.ˍ��˅�NK�a:e��Ӥ�&!���|%MdJE��P��ԛ$0��4�`160��ZH�<4�R���d�[�]�XY���̲t�����έ�in�I$��RDX��$�(G�v� ����^J%0��e�0�8��/&�f>ݿ���C�l����$����ߧ���w��-���|���k�w��ۭ����i���<������r�����ɯ&�z����k�����|]�9mȣ��ϟ�?�.���_|���d�ʵ-A�-D�����ʂ����_N�e�޽+'���j̳8 �߼y�G��q\��4�'�d#	�#&�?��#�&�L��x���
Ä��=wX�k�����^����p֓�g/�����_��-��Ε��?�����}�5۸�w�����1ox�ޏ�.g�f�|�0�e���v��~�ߊ�����y�1�̘%x+��oJp��ٱ_�>}ٟ���4��ڍ���oYu��%CȺ�!KA ƘH*��������d-�%_m�`b��b�6[0�*4��V`�5�qJcUX-0�ʢ�-�^����,NH�^���&A/�fJh�Ci��,T��i�c�{e��Āٱ�2 hl��&�	@���I�.�N�Z����0cr�z�u��MK�2N���\���>|�Ԃ�҉�S�6�÷�954��$�Y<�����b=��w_τd$�#�"![��31���*�����]#<NT��#��O�;*��q#";��il|�A.\ۡ�����#N{P/��{���+�'�{���	2RA�b\I&����v�X�������h \3��Wb�s�<_�4Pz噣��_!7��x�%�bh �|z0Lg�����:`a^ ���q,���e�'�J��u�
����t.r�%��"	�N�ĩ�ڠ a�D�S˺�&S� T 
Y�Ɨ C�� ����	�D�fu�����@`��!�h�S3g���7`	d(rJ~@F�8 }��		&���, �F�!� �S6���+�	�b��&����"'N&��6A����& HM���J <�0�'s�PIV�f���#I�6��e��P°�&I<z�bB0@l0jEo=k"�F��m�5 ��+0�����D�#�P�� (ã+	����$u�c�D��E/M��J�R��E����׋�ߌ���BV�%�EX�*��@	�D�41�'&�@��D� ����!HIc�DI�����--3E�4��j�Ic ]M.Xe�L`��^�1�W�3��p�&_�2��js]�H�`t�(�ez�؞��]Z�X�B��d���)��B�.���J⯯�E��k&��M��1��_�0�,. ��`�F�&f��:�(����t�3� q�2v�!@&*M�Qð₠���x��X�FϜ��-�dF/! 4"V\���'BM� ��Ta�	�l,�cw8Q% %�	^<�L��F"Zx���`1D�`~�:�0�LBK�L���FA+6]�Ȕx�x�O<���y�� h��R��&���"�'�`�� 4�8[f�	X�{ �ˇ&\�)�d��Ĭ�$�ꅤa��%`2�z���/uBş�5����G`	��w�ԋ��0�d������� P�oi�P0�3�p�`�"��OT� �>M�:`V(!��!M#��$�μ�W�H ��Ȗ�*xcLB�$r��}f�/`$
=L
 6��$�B�K�� ��Mo����8}��e!]�H2F2��0zM�
A<�q�Wif.�*=|6�Aetz�C2Q4S(#�)�h0��h����L�Քz�(f\rR|Ts
C�2���^r��ţ ���fb`ȗ&+ M�&d�!h�:1�9��@��ܾ����"T�9@�M2�fi�����%^/B%ׁ�;]��i3��ҥ�J���Q����ppZ��3��0�Q�D�'�{�F�����H��ɪ&�	;᱂Q?{�L`҂���Lv>���DA�Sx�����D��a�96��W��e������J��j��!Qd		M�F"׋�	F��+���!0_�bNo\R����d��V��#���w��	l��H��RD����`R�f���j��|)4��pS����;�R�B�N�kY$�bL1�G�K$�S���<�Xac�Hf5����	�,��
	Z��!!�͊Bk���H^�hp&�4�DΑ!��z��)! R\S�O"�@�m��Sj�L@�$<M�hҥ�
�)�\�#�Il�b N$�x��/C��Ⱥ�c�6F�rQEl��0��te����\���K�n5m���e���Ek2�/:_�x��tn\�+���|�Wo�.��xz�<9+�1�������ȫ�Y�g���'������M͝�k�ݽ��3yy�x����E����|�qo�cs6���zzW�ԥ�v�ܡt��|L.����Ƽ�2f�.7�z.�z��dQ}�y���_�[���_���[����E��
�~��|6���v�w���9� �=��h��Ĭ�{������br4�x��hh{xn���7�s�-��5��s{�jHAs�l�\��8z�������;��n]���<��������7�^C8��ۻ+�o=��ŋ͆W�zW��jte�3��9/^t2j���{v�n�?Xq4��;�z(ǩ��Hͬ�w�Pw�dwӡ���[î;��7�o�����ZG�rk�.Xo�6����v�S�ד���~6�HP�c�����w��s�����3�����!�[k7�~�hˍ�3S�ŬVK�o���]��BQ,ZG��*i[k�N�PGnk��d9Q[�~)s{�5�vs�O<6h�l���vˮY�<<���_�z��Hw-�L6wߑ.�K�Ϧ��t����r-�?���������C�������f��r��n��������O����k���Н�ˉ��w��u�Nܫ��Eh1Tc*�2;W�ڪ���.�uX������9ݺz�{|��ًM��o||�Q������/^[W\��6ڏ?��]C^L�Mm���QTqp�O�}�2� �<yB�qㆀ<x��'�d��S\p$�l�Ǐ�h�2�����+�6���?�؅_J'<f�`sN4;�n�������d����9ѝ�����>�Q�"�1�u	�X�xz�Γ����ڦqQ��\���/>����#+�s�;^}�=\���R�b�<�.ϧރ����pIs��=D����2���MJ��^-6JL�5e�^a����铮(Y�'(��	Cy��'. ���O��0C2O��LD>??}��7���4*K��~�jbR��ZIX�P��g�4 �^Mϊ^�`䬤�usr6��rgg�^�vo�#���NX+�9�K�Œ�~�ŲYN�Nd>����q.���g�Yo>��뚽�N��������߆����`6]���=ڲp[m�W��5M@^    IDAT�J���S1|f���4-V����_d&ц��o��ҧ=�K`�����M�-V��Bi���k�/�?0f��m!�۷o��ϋ=	/0S�po)P��=4��H��~���1��;�a��ל��>�-&�U���#ypc�ַ��?������^����yc��� ��w/�ܛD�t������ZO�zf��Ѳ<�x����+)���Y�lz�جN7g����d��g��?^�0��Uo?&ʃ�S1ѩq�y�zC�Z�|`@�d��Zoe�S����1�$�fM���d��{0����̬��*�L4�Ĝ�F�� 7M����x5�2��C-��+���A2�R���Bwz���i�'!�h!5Y�[L�\$~k�!F�!��D�AE@��^$�e��̲$d��t�IM. -Zk������N`n��VuS��܍7��-rwԀ}'t��I�fJN�٘"w��̑��D0"F�O���s~5y��cR�g��.M{�XD%My<�Q`6d0l�%؏��W�9L��g�ۖa��̑Z��p�p�cfct^�Oِ1HC0X���5B�0�g�{f]Z���~<��	�N#�p�X "t��,HN��D��	�.<L�k��ӒH�M�
̝;w��@V3d�e�P��§���R�#��"`a3�7 ��T�R�ɏ �x�E�V�a�H�4z	zE�t���Ǻ�X<h�h*�@jzC�5L�E�6J�u�0	� �-�!�Ny S�Պ����.�b#ЗȾ�<��љe�����C��(r��_���KBeQ�f�D�	����;~��"���$��k�q~���oza����&����!$ Y�QZoi
 <�K�z���6a���ԥIP`�rE��h�2.J�l��i2��腚Md2
T���g���6a��@��%C#`V���9�l3"���z��u��/�.lH��lu%z�5�U���I_7��c�9 M
/ܑ!�*li4ui&�4i�R\Va�N�z�XT�9�@L9��S ��� l(�L%M�$���lij~1��;~���<� �@��a�ɖI��K`KC�i�L�ɲ��3�სa��2�)6�}M�Z�H�R�Gf��*��5N��GS�I���2M` Tx4�L��Ѥ6F',a $����q���=�Fх-��d%'4�1�넍_d�m �\�35=|RT�.�-!a�ԥ��-�,ь���'NT\(F�8��_0r�Y�`�h�ń9Y���_Qe�qJ)-�&ZN��T�;<�`�ui)E��B.s�ϐ�<2T#��A\b�V�.E�~V4�0t؄�Ucؒ�QbKl>��B�B���I�
��l��G�4�LC��h�U�}�F�3��-׺ �dk�z�.r=5+z�;M�ǣ^����\���F�|03^�@W�&�#��~��RM�G��ɑA�)�h�<�BQ���2u\ӰJ����_H�z鹎w]u%�Y��G$Jr�6�����$���X�L�+ɘ�p�D3^�\/�ڗ�3�FH�0�ҫ�G�P����iB@ /!'(�������^�����>0�T�$H�I5+/�GMh�Km�=s�%?��B��i����c`+�&��kMã0���J� `�43|HJ<�4	l��*��C��o2_4ɒ:�La�B��.1;��$*��5�x0`� ���i�	F*`T5��%�z,�8}]�T2Y�8b��4�pG#�P�@��E)0�D��G+6�Ô�m|�Y�������On=8e�)��r˩��LZ�&�5rz%If.2MQ4Ɂ�8=���T"ǦV���Q��H<�ژ�d������(za&�4\ �A1Rx�H4�(���+3E��Ә#^��3	��<���K#��\\�D��`a�@��!f��U"d�>�%h�9��"𫗡�M�ތL��fz0l�����X��͑��B�Q�<$H�3��JU�2�V���z�ܠ�o�l�_������:�[�;�{�N�\~x���x��˯O��n�����޺�����7:�\�÷�Qv;[ݭ��Ek�h�6ww�_ye`k扞�z�]��=�zC�wT�Ϫ�)��mv�q�pu�=�VZ�-��t��{y��z@�N��J�<隹�׺�����ڜOǳ�˪������7����IPO	y:�<��8>?��n��eE�BZ�>[�so����ƪ�*W���5��~\�b9��X�{�m%��I�'��s�1&�T/�ݽr���ܚ���^����=���^���wv޿}�����oΦg�h�5��`̣{�����3�[����Ǔ������t��/D�ͣ3ǟk�L�KO��[�&�<��x��N9����r�r������o\��z[���U/���$^��S�Ჱh,�<����{��f{�7
O��<��??}|t�L��ֻ
�;Q���|���my��z�l�]��3k��0����^[�uh��;�o�զ�+��.-�����iOOz�T��B=�U��oX�]k������w}6��q>�u}���皼��馿뭮����3�n�{R�?�{�ۨ���t��3���A����z(g����g=wv7����Y���̾��M��:7��o���oF�<~xr��s��kK�g���������-�-�i�j�[;0��n O���j������?y�������'덣���7�[w|^����7K)�����x�V��4;�I�����n�C]>�����Npmَv�US�X��_�N��L,�*B�~B��9�r�����������'����?�BZ����\��QGH���]&>���=KJ�>��ʯO����8��n��@�v�4	t�������X-r��z�g��q�x����o�v�6�z�����~t˻���&��ӓ�d�.�ۼ���tlq�mq�5R�AP#����UҕU�)'�>Hr��w
]�ɐ������o��Y�2|c�!P*��e�B�Pڑ`�d�"ҥ�4�6~��C� �Vm���D���G��[� 8��P������/!�ҫP�ck�����y~s��;�F酿�h�zέ^ ݑ���m��S�Ur}�rʫ�84���_�<f�/?. �6����w��l�{���ẹ���`x�W����B�2F���_��s/�mzP�֭[�܃�#Aʦ�d���d�I���`�E	Ä�K��?~��f3j�l*���R��
��GO��큤آ�Ëxxa��6P�luѻo�� �H0��aW�0��[��}�6_v��}���Ӂ�RÝ�k{α���[�?�ֿ�����K����}S�ޫ������ǟ��M8^��c;=�\�H�_-}�Zi�����l��������h����扷��:^D�����oS�&�E�6"%��DP,hğU�(!d9�!a��&J5�a+M���G�zteU�c�ȡY�j +�\ �D��^>���8	C�
NJ%�j]�2���J#S
&���Ȍ���k��!�^>���Ea�Ш���d@�6��������,!��	$%CT��&Bh��a&k>9L����f[��S��	��+K�1��w�����[�q��}g;8{�2�W��@mC��(��& qp$C�wx��ǣG��{�Ћ��������;��O�T�d�6!�6f�X����\��	�tK	#	14	�A@T|qmDM ~yg"H�Ȃs�q\B릦����λ��a�Bv�Gb8`�P�,o2 B��n(҈�p�
������$���D��`�xae"�i��c�\���^Sc�e��T߻w�)I�����x0(��$zrV�x���7K���%rJ$�4�Ƅ�W-<9�rT4�
d�$�cSh��]s���J�fdu��M��_<���eʢ'g���R�3)d#b,�x�#2MH�<=N1Q���!< ��z�G"פ��D͗�& �:����d,�z@�'�0�)��_i�N����V+I����D� �����"���:KB�$�d dV���#V�H�%�� �Qt�)��Lr��ع`�Rѥ�(�y�B�D��A�kj�	'�޸���-�YKHx4͌!X�H8ҕ!���d�	�I��Ⱥ4�C�Ѫ5)��E�&C��)&`��K�|) b�^S��c��F!�*�k���f
j=���^�p&6�!$�� 5a�CK���:��)��i�&�`�#)ATa��`��$�*c�F��*���I?L���10�"��1�̅�.`��9��\�dJ�s�j�� R�(!Y���x��
�����m��`SGH���\zR�3���- * ��6��`j�A*b�a�+��DR�LRGI ������:x0��Z�Z[V� 
=�Ht)d��]B��RH�<�D�]\~Tz�|��^�A�qFI����B��d��0V���R�Z�՘ʜ�EEP���:c��`,`� Ԕ<����e �����!5|��Kج�8ت�,d0M �e2��AS�7���D�E ���^/� 1��3�Ox2C���9��w �/�.zH��	^f�>���cZ�L�*�L)T1�(�h*�}Ƌ&3N~]�d�
9��d,�P�k� �5�R��^*8�&۸KҘ@V34���ĆC���fiA���`�� *xMrL�yQ�պ2d����Ⱥ��u���X�!�T׎��Q����d ��M� ��KSN�&�&=C��$(yx���Ƴ�K/`z�j�:ۺ(��QWF�H�k�+�0�/Z���0�ĉ�&�e���	$��#���_��|B2�W410��ᥢ,s���l�M<�!a���Q�E���F!��/�^&x0�ب�GJ�u�酡O����TӇ3�bBɐF�a�DN�dEP��:!`bS2�z��z����G��^��C"�%��FG�0h3+�F�&0��!c������D�$~i�"a���*�j5 rud� `P�K��*��8C�?�k�	 I��g` �P�9�4pL���"���U<�8�R�:)F��:!q��Ň|�<��+Q�d�j*R��IdT��Y�G�9�&���+%W�h"T�G�V=�:{5u�a�ԛH��w)çVg(� >��sWJ���"���梲7����n�����V���޹u����A�廬p�����Q�?�?����?����j-\�	�=0��H��N��ק=Y�ozo�b��i��nd��g�r�}y���lt�:O`���D�\�t�q�w�\y���h]�ϖ�jyݭ�IZ��׎���xV�C�4���']����[�V��h�i��)���d���{�vwӘZ�moP�2\o|�v��=pp��ٽ�f~^t>�����y��$"o�++�b�;,����oӝvg���������z��B��Vk3�JF�:~��zr�߭���[��~b���O��۞D����G�N^>2����i��왗�Ǒ�+���[֏�������]�~��m�?\����^����^�4[���2���j�׶�˭�[��Ψ�WL}�k�{G������'���;{����w��7�h �F4@P$E-Cj�H�41��-�D�D��G��O�0/�p��Z��2��! $�����wo��~d�ag �N~�;'OfeUWݪگM;&��n77@]��2����;��l��V���vZ��q��[�[k�=�{RD������B7���jK�xZ(����O7�����-x���nj�����/m���\D�7`;�μV.$j�$�'!��q��]]n<����G{���K��s���_<w~��S�.l�}3e2wٛ��D�n��Κ���n�L��v��>>=ؼ�u�����{M��|�|���>y��e\���a�NG�Y�����^)�r�<�9�YL����T����3�;Owݧw|;>*ux�֜���;>r���uN�3ɘ]�t=���j��U���؆`L	��,<;��eI��Y!�t��8ɮ� +�k���s�Z+��~��nUr�������b,��^���e���c���,�����M����yq}،�ys�T+f���hܝ;w���Z��^���2�ivG��r�j��kwo^���Xy�p�?���ew�$����y&ӟ]X�Q0e���b�L��"�(HE0Aj����mjʈ���* K�$� k
	���:�K�EU6�2 _�1�0�Uh���B/��Թh̶y��-{�I}'l������g]� L��'�S����jx�aBN"���+�:b�x�c]m�9/�՗�~�`��2i�v�)���:������9�1��M��eg9��Y�v��[��5g�����7���՟�d������p�a�Y?�n�eo�n�f�����D��Pꗩ�If(�NwLS�J�i��.a<���
x����=6��x�O�%��
C`�=�M���qd�3�ؘo����p��$����}�����{�g��x�u6;k�.�o^��ڸtnt4۸p����|u{�<k���8ٛ��j������/S�3�Aw�Y���3�ֽ"��3f�P7)�!���Û�����rPYrZ599x6��k�NϜ:fɼєh��u!ӆ��Φ�rBV��Q� ��&p�ɜLCO`B��Xi���!5��,��l-+��a#s��2' gN�a �_�U`iR+�Lba�4�JG��u� $�
�qW'u&	[�0٣ahl�}�����E�MzTvK�&.�)c1E��+�xdb�q$B0ˋÆy�ʝ*���ז!�����/qҰ��1D����?�dFb�G�ߎF+C��5���Q� ���?$AwB�UXu�M�x���s,�HwI��^z�Dv%�4~� �l��d@/�e�k���E��]9�^z�/"T0��Z�w{�^�K��{���K�$����0���� YNP��r$¬�%V���;�`"��H,�x�i:/'�!�H`22C��#�;	�d�pf X���?x��j��̹&���?�pI�8-��,ϝ�; �3�x������B/N���3D�d�	*�"�ф�&�O���Ȝ@+!TJ<��D�	�>&̉�����#�L�Z2	'�R��D����U̚tG��>H�	j`'_��r��&��h��-a��$�`R m�W��H�ºT\�6���iDb�ؤ4�^�֊��BД8M�q�4��w��1fM���
$�h��h����c�M`���a�Bk�H���N�af��@B�0�4� U$Jl8��
g0�1�0aZ5�W����I�/��d�h�0jC�u�NPB(BJ`E����$BJ���@4\�Ш�C�I$ٌS1P����0�MN�+6a*d�ÖR<��(���h��I��9������01h£�8�Ux4��-AM�h�6}�OM5�xa2C� ~J J.,��c��Y�3(�iX�D�=��PkF�^�Guh �#x2}�z�,0=@�U�{%/i2���C��o'�/� B�"��T�S*�a�����B�!0-!�3	[�j��Ux�1�>��Q��
F��!!��$��h-q|>mL9��t!��@I`���:��(���Pk��D/�	��0T2�y� f�SZ4b�^`�O��"Q3�I��KA�!��x4L*&If��Zk:����HB��Z^(Sc0g�wu���`:댂�/�
�&�1�\%'J~)y���F�M8a�u� �6�┞ߤ�y��?J`V�4�d�$��
��Q��i��[��	@w���u��$�"��J�~�0����	f�HhD@��Pf���&�2��kMaCE�Ѥ$l�l���Th�Qh���)��Zr�A~m҇�	��/���0J��&JTl1���7��Z��H��!�5�W3��/d���;xH7�'T0�j��3�-�Z�	IFE�6'� LrM�њbLS&R6B:��&5!����i��/r����&~��!HaB�P�����5��$lI+�FIk��aJ$�0�6`2�����m�i�)�"(�"�K���l@2L�`�2����M���Zz.���$�WB՚bӠ�[#���[��qA�T�+�����Gl1�٤U����S3ON��F�pU�    IDATs�L�D�%�l҄�`�$s�O%����MYlEH6��H�i�VJ9�_	��:ON��A��a�iX%65�:Д.d��*M�0dS�"MdlH��bv�*� B\��kx`0�RͣB H��/�x&`���D�(A2\�}���������^ߍK���aZ�	��xQ�_��
�Į"��0 �ZI1[�j&H��@#� �I�
N�d�̇/fs�PYg�0G��e�\<qa�#�ts��-H�!g�[����/����ŠL�W_��~.x�d�һgS��\v��h��FVw�|�w��ֵK�Vwr�/%ɮ����f��,��n��Q�O\�>~z:�i;t��t�{ݝ�}w�:#��di<w��Ұ����|����^���m�=�5:��f��_5��|��`8�P��Vy�묱�d6�38:��KmoG�x�d|:q�ҳ��'���q��>u[�3���sثR�%q�^�ti쏼��Zw~�㟵r6�4�MO>����K�v����yc��[3��ɹ����2��}��Ǉ�����g������x��k/}5��;q�R5���y��U�b�q�����N����Ɋo��x9�i��M��9M�nJ������II�ѳ�;M7�<�囖�S�)��uT)����kn;��d��g-�t[n�֭!����lt�4���g��]�i]���Z�5빆O�g{<9�P��^|��?p:Z�n�3���L	?�Q��ܺ2��ٸ嶥����Q�sf��j]��<�|�j�{v5|�����n��������4��ܓ�^Z�u�������xZo��G�&�����`4<:}1<��s��< 2@Ϳn���U���gnm�����\7��:����x��bg�����r���k���j=���'@�'������{��YzmS)�zq�CC�Y�[=�5��<�Zt}|�M��Vgn��ݗk�Zvy����Ҿ�������OϢrQ����Fk�sQ�ŗ�������l��3����VJ;�]^ �tuW�4��J����`ma��k#wF=4�1�,xMo���k����W�2���̪�h�<˔˰���� ]>u������?��{�|�����!'`�,p�ۭ�۷oÃ����O�b������g�/G|핻V��}U��l�\��}��ݭ�r�C�~d�Il��g��W>;�=J<u�Đ��fDl
�B�YN�����޺����W���MC�8�p� QkRXA���n��h�����:TRJV�e;���鼘	.�У5�M�w)Y�t�T��Ł�R��� P�A����糙-+�D����Z��l�N�ϟ��x���A�1z�e��Y�O6�e�C�gf���6o�.��;���R��;����5��O(Nz�م��uK\��I���`}��lrs����������=Z?�)�H9��1����Eo�>>�M���ݵk��cM�䮀<ڻ/�?�ۼW�gd2�����nؘӲ����do灔ÙkUre�����W�4���!V$�kǻ}���u��.G��.{8���6�������g;���k�yksC'^N�~��tg�/�G߿릦�����hit</���r�Ё�	n����-�R,Le���E����U~�R&�_�h��7;�
���c���G�G���~�u�m9d�;+���1�U��y���D��r0[�l�(�4<���j1��)���46�CIX[�x&2AS
%H�P�WL�C�I͖��Ch��ᢱ�/��X�f5pL��aLia"i��_��
=�̑7B�ΪN�6	�a8x0X�M�'O����1�x��j)7s�ɋ��.c���,����E�F���Ç�&~M`��L������tv=kT�c�pn�H�D�av�
h�]���.�G�g9�Pf�a�;vC�Q�J�#�r9�Y�P���Z���;�=z�f{{�F*��G�"�G�1-�l����x�k	;���#!r�<94���$�w�ꗅ����3�P�#�=a˞l�2Yk�i�OK�䠒� ��1�5��Y�N6>��#$�R��z���Ԥ�)� �N�6�B
��3��w�ܑ�̄���8]�7�'ZC���4(������,3Q%B��)]�d,�G���8�L Ԋ��U�Z Űf���`4)�:�&��*�IgE�E�%\��I�'<�_!�a�`x�2CO��V
&�b������P����>`�d$�N%$��!��V-x�Φk�\�1���4�l3aK×:N���� �}F�\Kc5Dh׋��F>��� a�)���L�j�%i `�P��M0����4���L����̱%�dQq�dz�(6��ő��0�(���9w���B 
NM��N��#s���(6��|l�#pMIF��`��l���N��m�D �6�6�[�!�%Ŧ=�k���.�O���Fϻ�r�< ��V�(?/��"�^�d u
�M0��#����]kR�B�$`��D�x x�`��w` H$��`��0q��J!���IF�B֪�V�� ��KlY��&&�dH � �I����`��&<`� d�XD]F����\d�$<��c!$=LI�MH�)Z�Mw0븒�/�X� `2r&A��Fj�!�i"GcO䗬V�h�;2�&�����@CFL�M5�2}���x4���=A�z��4
A��C$�J�|�U̼$��D��^$��0��i	9����f�x
r�����)=C=
 �
[��M`0r&!N��VxJ5�����I%Cˎ:x3�
#Ye"�!+02 ��p�
@/��sW�m+ �&�
+)Uk"�?	2Jz����f� 㔀�/��;��:�DNPb�f�I�
~�Ԅ��G���5̑B������24J��x�'(ऩ���;V6�y�!�V�D��"������/�x��L_��x(b $�iP�(b���0��:jz5f��$��B�V���	�>���R�\M	�]4 L��EZ1��L��;K��PC"�tG�a�F��Ԥ``���&�^=��1�����B"<�`\���S��WDB�(�06�I�0� �5@�M\h�����(!'0Z��/�*1 ���R<l��IX�H�Px���ë��(a�2G_����|��O�3�2��ɵZ�$��D!Ȥa6���Sxa�ӄD<
�F)9WC�
&&H�����$����k��)i�M$��b\��]6����S�£�-	@�ү��<�FH�@�I����rz�
�"�O`̑��dbĤ
	^SL��`4a3J��"=*�-�����f�1ɬ���8�.��)uh��L�ē.���I��ޅ6�a��}��"AB&�x�j��0d$�IEbpD���Gu��d@��`32�_$Ae�#hu�b:.?�v����-�x�r��d�ۊ���F��{�k�V�(\�k\�XM�ñ{l�Υ����˕���յ��ۉ�(�i�x䣏��sɓu���=U��J������=͟���ݳt�� �έ��zS���޼>������=�w49[�z�n�8��m�[�u�sևy�{<�:���z�h�y��ŋ+���+[nx��������;='����y�lz:���E���|i�֭�����11zTs��V�L�W:d{��xY����m���>�f�<�Y��_y�qz�>k�c�[,>DfL:k+7j��N���������v�����fS�l���s��[1>Љ��^�͞��/�ۭ��ڪ{�+�o��F'�é{6��K�Ϝ՟_�(�5�.^��h{��ttx���g�Z^�j��;]=�c��'���+w�}US'��=ͺ�Ys��.q�H���\|��y���\��^�l;�6<F>���h�����wzns4v��K�:P7<��(�:�wZ�F�Ys�9\oeu?Ռ=�5Fgc��C�eϘ-������#/��IG�n{٥����Γ�/vη��|���yɥ�~�?�����6ګ��-�>����h���u��"c�'g�Q���r��Y��Y{ٻx�~�����N��>����Eߕ�yy����`�6n���9ܛ������:rw�Lv�f�a�ص=��[�����SR��Nw�e�^�=ȓ�;��Qt�}$rk�3M�U����:����gG���>z�z�.�D咣?x�^������{�}��;���Z�������ۊvs��s��m_%�Ν3��u�R�8-�;����Ǐ���#�suZk�!��芥+~��P�b��K
� ޺uK�s3M.�b�����w���{��Dc⎭�O>����%��޽{:h��[���n�qn󍯾�o}����h����_���7������Eͧ}��f9s*G(��l�,�����k ��M��MM\k%(���@�E�M0��5�dJ��0�4�gU�k?Bá��']QZ�yLM�ӹ��Gb-¥`��4��Aiz��Ev��|s�X�M� �ԂK'��L!D�dS(�60+�t)�Dl��ĵi�3��{O{����t��ǚ?�-��+7:˳���E��_~[P��('�%��t��:>���+m?Yqô�t�~��nu�\��a���9��=E����:fc핕���#�쓾W��f�����ɌZ�?����q��F��E�%�Ff�F�n���k5��f7T�3���r����%Ma��%��+;O�����W ����ˡ�A�)N	�dG�.�hy����qn��ck���W�m�����G�Q�Q�k����[?���}�V�{5G��u���?�S'��rv�ڴ����oJ'(ܩ9R/��wX\�K��J͛��>b;��ǳv�[��p�����g��|�d�����g�_8���Q���FMY�~�������&�"��f٫gc40)��.��++��g/�7x�B�	@X�X�u��$Ju.T��0IB@* B`�h9͞��F+0�T�MII ��9�MM�x$$r�m���D���/�2�4�r�~���^mN�H�/ �f�iO# ���j����5���n�-*�\�P�P!��D�=�rG���a7ah��T���?�0;w�4�=lX�����7��@ެ�"�@�������}�NTN|CJ��l�ਃ�wHLVY%tD���0����%vs�x�ҳS#��2#0=u��>bC�PƸ�D�	C���LجJ��{��K�ȹfEIc�_Ţ�J���X[(�2v�dR�2�6�
ZM�mJ�J�~ �!4�j��d���0�g� ��(�C��ȁ�p������Nft��������G���𘩅[�W�hB��	; ���"s&������?/�T�� �a�	�xl��*H�s�AA�N+���lZ	J���"���`�IJ܋A�1�8"��/�����	ɐ�R͊?9�\�����#Yb5J^��쥳&}���HSbX����@	 w��/Q�#�/�)�)Y)��4��k�y!7[�mbӤ_:ȵ���2��I�,2=&��W���$�]�a����N�O�aJ>�À?A2�,�jJ�`
@��D|1�Q�J���Rm��� ��(��a��Q�� ��6�
Rn�m*iDh��d����ܩ��#2!5�_�	=�\+���'�A�)H(�_���L!X�0X$��rJ���*i���%�8�/���	�	�;#�f�^F��Lm�*H8�_$��q�,�A�`��&EڥE08�1�}W�Ɗ� �i�'3��;޵*6F(����F�Q�:$V��R/h>k2� C(~��Dï� �J��t �\pMV�V��8���JbfBC��J&��^+�܅3�$H�JV��P����# iv��	��l*�V-ɉ�����@��;�3ml�M�b�FN�A-0�`�}�0H�r
C`3�&1ךnjʬ (�L`�;��-z�)<��D�-}	�!ƦZ�H�	Q�g� �ٌ_2��	��H�U���fx Ҁ%�S� Lp$f��t�!��mL�QS��I�O���B�!&�p\ӄ�R	g+�&��l�a.6V\���Ca�$��@���m�0�DN�0�D����l2���J�D�8P���E���,Sq�x� �c�(~m��H��Y]䜢���>d�i�ƢĴ(�(��Ր^<ș�9&f4Wl��AN�E���2�a�'f���xA�/�0�dk�`E���U ��BK��Q�`S8e�H��T! X06�g�.�x�3e<��ZU��%~M:G	#�6e��L��8�Q�Q���}d��Za�L���*w�Ͱ� ��69��0'����b$4��D��	� ��cS�	���!Ġhb��&0sr&A1�LH�U�,�K9�z��2�BS��ȦZO!a[���P)*�
������sċb3N+=s�ie��
����_� 5����Y�$`K�4EH`���󘄄�^1�C&$6H�`��Q�*ƣ��U�,%�j� ���r����F ��0�B�s��'0���a�m�r1�0S�$�T0ËP����2NKFkW�� .ԚhR'9�y	~���L���K�S �5�,Đ����E��q2��/H%$�����H$Z�5!�1��h1�l�d�b�,��Ȍ��<���#L�d�w���6ԭ�'#<���bpQZW�J���!f׳4�5un�u;��##�n��D2��`¼��x3������j��r�wY�ʳ�����;�o^��,g���k��<z�dwoP����9�[_�x�k����޼qk����~���~y����>.�y�]�}㯾��[�.]�}7e��p�u_��ǂ��������j���Jz6���/��	Q�N���g�&�Q�S�.x���]���.O���/n����|!�N�5��6&O���g�(�5{w�Z���z������{G�j�Ӎ�^}���y>�Tm9ztk�ᒗ�(l�ϼ�Vz0L=���®'	����}�3�k�ͣ��?����g{�n��[v��s�e6��X^^w+��O$�e.�75�^��҇9ߘ����;}�L:+����Ps�ElaۛF{3����i3�v�yôvT^�:l4W��w�,��,���m�!���\gcW�[��q��Ҟ���=QOK7�V�Ƶ��������Ҳ��BL�K�����x8=��`�㙼r�fH�68�y%�Wc��]�/>�r�$���KW�[��WF�CO�Jk��:O?��ɳ����'�������u7��b������z	�rw���ўw]=��l�c�V����(ź��jy��a�(Z.�Y�P)S�&�,�^��d#��%7��n�{���_}}���O?zxt<>�'���+[o]������q�[-N����?�����_t�A�\80����6�߿�B���VW�<������|�;׮]�裏��_���UDW�-�.���,u����҇ş�.��d��;��M�r�����~�i�[<z�Y�frdg�� W���ƍK�h)݅e/{6%
�k��(�®]�(O�������u<�D�������n��*�'ǃ��lp�t2,�>R�U�E[��W��2��7uPxR���
0+`�(�C}6��H
��O	��fSS���R4��8�a�����q����*�;E�]����\m�2Rr�t��ʕ+l�:����
"�f�@�n�@-G�N�{��lZ��e�AV��sN����@��:�wp���IM6;�e�=%����Z���(��=�C��M�vuK�EnQ��]`��\�|䯪����{���Ƭu��5;��ϫG��������p���=?��FkXAs[[�݌p���i�r�%��U!�K���\���d*&�̘�Z?��2"Ókd��;��`�v=ɡ��24�����aN��S��y�)W��`P�A�&�w�=*w_�ˎ�j���u�"�k��^˟�~bଢ଼�Ο�������Ny�@m�\:j���#��.��~Ub�-���M�~.R�s$Z��c�������5M���n8�̴'m�����\&����O5��V=������g+~���[� ^f�4�I�1�}7C��ْY�P�-v�ē 0 �(�d�L��x�&=���m��$ ��i\��	?��MB���M���̜PY��2q�^�͓�    IDAT$&,�J���:B�' �� �`0�saWΘm�%-`�0�sO��QS��x4����l���m�a0EQ)�����s!i�Az���o�g����V��Y|���p;ThJ���8�8�����m<����۷o#�+�� v��;��[���D��;w�ꅚ�U��&����M��T�d�9�=|�0��}�Ϋ�w���ʀh�@
�G��Ʉ�#Niܰ�_��_�)r��꫒/Z;��[�D�:�I�}��@H/�'��J~�	E����`���	������@<d���� �[�Qi�:�ǲCi��Gy�)�cG �UA��Pʉ Xp���H�8��L!�TX��C#Q��G+l :�I�_Hz <�&z�6R�����t!�&<Z� #'\�Bx��蠱K++����j&�n"��S�+�"j05�V1(L������Ө��%��Pfe`�wZ��'�J8��0��3�M����+����F�	�$	���x�x27���ޠ����1���/r����n�A�)c�PSb&W�sɑ ��$T���FOf�ȵ�~��b���V~� ��J�5��0��&<���a��rz��¦0b��q�����)V��\+�c+�dI�ME��h�Uι[2$�	I���v� o�q#^tJw��1�G"i8�$N�`HC/�h{
~��>Zk�m
U��Y|q�D/��K����.�9	%�j�jM"Ѫ���*�-��D�Aj��4 �<
/l\G��dΐ���J>�f���&fz0�9^� #T�1|�i���`�Prt�RF�E��f��s!<�Z*�~1�j��BQV�$\`���Dv��F�C����P�)HJF�^@2L E��0��1��&�h��
�5���08��*� I&� :LHTj���!�+<�R�$��h�Q��YM�U����+��i�ʼ�X�&�d���/6J��Ĝ8��!Q�h2Ka��t��V�(�ԂA%����τ��x���]T���"{0��EH���:�P����&�6���"`_����*��w�8��Y�0���&x�pR�M��L7�
e�_�x�8���A���4��F����ީ��
O�V���S�P�! zmf	 PGHG�H�:fM!�IlL8UkU�s�wv
�&^z.2��(�C��V��J�F�,�į��&ʄ��h�M`|�h�9Aa��&�)�`��d�"1�4ȳ��	=�����+M H��D��E�\#�L�d��G	�,xM��Z^~�CfK��%.����ːؔy0� "a(r5��)=r�/b�Sgt�&$���S���k3��$W�V+0%޹�T�`4��M\/�%�BHz�SB�=�6��>$Z5)�22[1�?0�H���&���!c���xlf��d3�`��V�l3���x�]k�I̚� �G�jz��cH�BAI@�SU��h�&�bK_�VMl!��� ��RB��!��1 �D�' M$��Ü�˔�<f�<�*��$C�P�y>��F�N�G���"OV	����l�i���f�t�s��il�e9Y��k
O���0��9%!��H*�Q��T��U"W3W�C��Ql��$�B��ɚ�(��`0�(:w�Ѩ��{4)6C�0�4�+�j���	̳SDiSw6Y˘�2� 4���� 4�L�M��l T�Ȅ�|���³"��T8YQ"L�j%.�䨄��&8��Ԫ�T9Ktq��K\��Ƴ�c_��VW�{���ӽ?�{��������ry��EK������Y�.��q���#�.��_���D���?7�\�fW��]@_㚞��+��l��*����������������a�����t��������O�x��K�_��w޾��W�^�Ε���y�`�x���>���	�{�Ɨ�����-���x�.�Z���+��ǹ��v���;n�fx�3eFq���_��q��']��c�s��:���s�ư��q�C�nڹ�V����ng����30��(��O�'�,Yv]��G�> ڨ�{]���ֺ��:��'���u=���}�U�Yu�4^���f�U�fk��3��n�����_j����޳���~���Jsy|:?�.]�ܺ�i������Ro�.]�X_�t]y�|M9.7[egY�a9s3I�7[�񭻞�v�8[n�h:�N�����h<ڙ������ㅍV��_y��W���~����x�S�zq�������_��R�y���_~�����I��b��Y�9��O����vg�|��Zgu^w�;�~��k���h�O���7�7V��r/ti�T��p�--'�C�V����,�X���2�,[���wO����~a�>==�;�YY+o�O6�7>��_~�w�����h���<O:��`9c�<�y�¥������y���oק���鷿���t��P��޵�).�r��ˆR,�:���jy�)�$?�>+���7;���Vge��͗�;��'�>v�>�a2��\z�ko^�t�`��_{�+G��ߞF�Bf�)�_�z���Z�G}��V��؜Uxh�2˖�k��X:`n,���
3�+�����?��Cx�P!y��w��藐����֋���J0N�R�Z;��|��'?A������ƝS><�>I����~���8��;7�%p�������������W����G�'{�>�i�)˩0d�F�#���w	Q������2(�`h��6x�%�4
���|��2��r�
!��9R�	F�(y��tD-��Z� ��Eoӕ7��������gHAPi�&�ʽ�h�C�(0�+�8H7�&hG ��U��.v���餷|+�<�퍳^�=x�x���jn�u���G��(Ip��^�K	��Hĺ#5�{b($�!{y2���S�J��X~�W�f�Q�>_���ʵk/?��l����7_�N�Νow�1ҥpǧ��"W��*)vwA���Q6u-sZ�LzY�\��E(����K�?���*�>��޽{;�l�`�������Ȩ�"Qg�r�Ѿg,�{��K5Cxy@`y�Rlx<��w67�y�>x��������|�j�q��?�o�uk�6��.����vw&����t���;0Q�!�|_��W��o��"�馅V�g��g-V��vÀM�ӁG��f����ӏ��ɺ��z̼�����e��/���e�4�$$�� �/���oA���& "�)��@&P0����Ui�㎭"T����Ė	�V�&}6���s���0���E��
��>�W��]Z%99M0��< ���`ԊV1XGĦU*J�����p:)4���\X�s���kw��&�Ml���o���T7{�����mB`�<��-�c�	w��;w�8���b�k�ap�;{����Q*�; )|����#;�{NKtJ�\`p��T���cⷷ
8�9�Y�9����J i�����B�5)U��t��ًu�G��H�͗>J��%?Yj�#��$�kH�"@�:��!�ƅ8qZ��޽�4w�F��뾰��$`&}�E�\$��FN����*0$#�hү���0�~a�*+ن��L�:)�d������T�q�4�2��&��$?N/b��S�@�����N����D��L��&5 �M�l�g��h�M�M�7p�+7{��1�?0��Vlҫ1�#HG��皐`��X�I`Z�(���lPt3�b3<����Ó�MPc#$Tr�)����'�	�P�!B� T�};�l�I��QkfibKVt�E�b6R���ox�+�UEb�7Eyǆ_1pBk��8f�N"=�N0����gRi2-��$l�%��H�ؒ�5IV���Rf2��� �@�_ld{�� �_z�2���b�M��R��)��LO�%����f�+����$ H��1P
ɾC^�\��L&��)6a�hz��}���3��Kl�hy�T��$M�)�"�n(*�EhF)�"�Ĭ��H�9�"�Rx�e�Y����,��"�jC�E�eFi�a�P�K� J�� xA* H41�f�T(L(-Aat\�Ԏ�ŗ�X�����C�5Z�s*H����_B5��R��%�Ո������k=�T�NZ4�Ȥ������M�M�Բ�6�Ug�g�@�l�`B*���3M&���9j֊�b�B��C
R!G�IHj���W�bK��(E��+M
�
Lȅ����H�qA�`6Z��f���AȐ@C��o4j2  5�¸��B�K��1�d.K�Flj���ìUB��UfE��?Á���P�*i��7�C0���1�i��ɒ��Z�)� <�
��ݤb.��D�DTNƤZ߳_�H�9�x���dB�Ha�,��� ��B�`��?��𺐹'*�4�@6��A�)1��/2�U��� ��͐�V�g��w �"~�x2��m�
�2#�� ]���5�M H{D�#̔���P���_kH�0::k�����@����UmP��$�@`~�9��j@�O���-�I���Qa�^����J+5N!����dSb�&!�t	}�&|l!a��S�<��ؤT8-���ʠh2W�B�>���y�A+��d}�Ƒ�HoZ13�&}�ă�� �d2	 LC�xI<�"DE��&�j�M��*ޱ�U��PsA��/��9!CzT�	L�i0��)H^��)a	�*��凹�l�M6�f�ɐ�hē� s���/*=��%Q�}��||���v�䓜x� :�0)��6rhi��0+&"4(�h'p�'|�G�0�Qbf�M0S��G����z��pg_�G5sz�, �E��٦�j�aHw�pI�T�s[���M%�����6M��ïP�Ʊı�$|���GH�D�̈́�4�hi�M|57�������"�dJHz���%~풔	3Y� �jy���� $�6�K�)%��UB`�N��(��-s���V.P��Z�?L��+�!O�h��t�	�*�� I�)<�x��V0��RG�]�w	�M05$�F��2~Y����L�_2|B2�63ID�ͦx�BI��p�{Z�/�IC���%(4)�Q�!��ì#℡_`K�Mp$�qs5}�R{��Ĳ��J��x0>:��W��]�|��h�d���坙+������G��JC[>��1/%��[|GЎ�N��W�UԌrK��tr��b���g����*���w���_�ƕ+bs���"n�[��w�=���O��������曽ns�֩���M������l����^��z�m��m��'��dV^�Z>vܯ?y:�Ŧ�gD=���Pc4�9��W!wY��lq�b����.�W�:-��߾3�pi�c�nj�|j��/������E����绋��j���V����������؇Ow���t;�._������?#\�wজ��^-ؾ�oϋ�^�q��FgՓ���g���]�����zb�>������4y��#ץM\�_6v�.t|���j/�u���L�Z�%m�s��,�ܽ�!6gZ�������-�,�|�<[�y���ӿ��~٦�u���B����@oܾ�l���ӳ������w����6�-u�{%=��Œ�=���<n��soc�{?����~��沏��?��'z�����cu�՛y-���JK�ݸMF�CY+;Bɯe��Ax�Ny���+�Ȯ���u�+>G�?:9��~k�g�֝�v{���>��^��{�.��݅��o�z�Ν��ǝ�R1q���A����f�w%�5:�Ӓv9!qJ�[Y_읟-�v|!���>h/�#[	U�*����a�\אַn���Ǡ��_��Q~Ҵy�\���(��xjau����;;�)�r�qqstp���6��?�}۴�T���/|��Ϋ���7�$��?������A�������w�CZ.���g?��9�r���0,&V�w�y��{�����=*6xl�(0R���I���H��"<�����������f������'õ���97h�>y��ҥ�_��/����{�v=�� u6�̇�e�W�A �)�h�e��Sc�Ҥ.���N���P�TZ3�d^�i%�è#�;Y!KHE�&M� 7ax�%�d��){ժ隉Aq�#і����#G�L(��EL؍D�,�9=e%�F����f��TH�}�֑��B&����{�|��r�Ȝ��Dm�<�'Y�QM�mΖ��X�C!P9+�Fp���)����HBc�����٨>Z����r��=�n�}ir~�������~�2�s}��O/��]�����޾�M����s䪢?�pvsZ~tP�*�z�HO9�kJH��o��Q����;�7H� �}^��(����AE�g�m��IвR\`���w5mw��� ر�S�1�w�<=�^��Zk��[�]�輴us:���;?|��;NrΖڎ�gӃ�g��3/7� �_���;S-SzV���Z�����tGq��A�ф����l��O��~�"�T�, �����3o����ć�[e�5[cX]���E�E�lr']�
�F�J�I<�E{٣*� m��)�3��~1�X<�*Na4)L$
�:�x�����j�ÃU^��Z�KOe.N`�%3�*�]���ʄ����P�̙(46�"�6�j�d�GMJ��T�L�5 �&^�6�ZJLNWd2E�0q��$��l���. a6	�� �:��Ŋ	� �PGP���mK�\�tu,�@���1 �k=��]��=����Y��B���"��V����*�q�^&`Vzᰄ	[B0N����N��9�(<r$BiA�C��h��,9�N�"xXuy��/p.���G��&0�w`K�%�#�O?�T``�apl�$���i_���^�^��;��/)bb��U"��*0�8���m�O/hشj1��٤�$�,9*߼y?%���2fJ���fb��I	)x�K�[E��Eµ
�	~�RD��c&o����rG)H NC����@�I �[1�Vʨ~�F���t��L�&� ȼ|b��b��#�b��G+apJ�M5�����FV� h��G�i��1ֺ�@J0��3�D"Q�ך�&�8��J`�9���3�k���4֚
�!_�^r�M0��W䉐��%R<4��6����EK�`�UL��"1��FH2��/)R�^�yZ2׋��ٛ m�I��?�	 �HK1��-%!N�@�SҨ�cS�Y�ɤQ��0��'�~afM��T���*q������oݺi��Z�Ni�=YM��]C&bH�Bi+�����&1��p���&!���O5C!A�9�#K�`,Y
Ic(����LMVW�����R�gVs�kM	)˔V���kve�k�T* D.0����9]L�I<N�b# d���Co,��"J��B�)[&�L�tʦ�t'H$�&	��dK�^k�=��P�r��Qꎒ@#Tux0�.^�9��%�YH��Aʱ�>x��*]�%1 !pj�d)I_�X�`Z%3��!=~�؍y�Ъ�
xV��&�P��i B�6O�Y�*aB/0<زa8]�ؘ +`�I�֪)B����)�Ʃ�o�aٷ�a�R]�Wx�8���M���׸�����2��9�<H�M���פ���l)���6�'���W�\�"pNfb�z�N7a�<���B��(��R��a��Ј��(����/x�ï��u���D�"�V@ꔮ��w��j������0I����y+E+6CO%�<����\�r�ۮt��m��.��`1�VEed03dE)xEG�Yǋ����/�j3�/����*m������s��$*�RʌK*��%b�Z�%\��̳�^bm"Ħ練�Bl��1M\he.{�3���%f�V��B2��h9�.��J+�N�y�43�he.]��JG��c��#sx�r�P��/����5+C���\"kRg^Q��;�m����rj�H���cs�&J����`�L�X�T�4�Xi!�����<l�
 �������l���5�@�*�ab�)�Ic30�BZ�.�p�仞    IDAT�0P`VQr��i���&T�$�&V"�����&0A�	^��&Bz5ג&0&Z�!�`8)��YE�*񄊹�Jd�K��s��2LO3@�R����#�)���3C��������2��&u��h͂��l* ��M����.�D�V�=lZ�( ��0����W+&*Y�+w\C*���Y��P����ӗ����x��*��!�C=�a�0qG��&!�!ÉV1�0G���)��x��hӔn�m*0& J�[�F�|��	X�j��N�uSJ�m�
�M�M%������"�qD�.�AT�C4A�C�z� �!3�QrƄ_ �j�<$�8��Oi�� ?����8�0@�Ǟ��G�2Q�%ωD��^�3MLl��h���=v������e�p��[�Ӌ�[O��lnN��}�2�K�^���[ea΁K�|V��8\(���u.V�MU�s�ˋ;�	������x�i7w����[/�y�Ð�}�CWa'n�6;Mm�]>w���j�kX7j�x�Z��z�٠?[�O�#���JS�P{��������?�L�"]-'�GϏ>��#˨;~f�+��?f�r��g(3�J�|��TޙZN���!
�����^D���csŃ�n�ͽ�o�� ��-fBɨ�-�s�d����#�{q���os�ꬶ'�ӗ���ҵ+/v�=�b�qwp���o>W�.ڵ�6n嵭k�����l^�R���ٰsژ׆}��v���+׷fKY6����mc�<
�]7vJW\��q����E�"�㒫؞;tS�M�f�2=������h��[����L�ڈ�4��ڗ֮]i,�;�)ͥyW~� C@��v�a�um|�z�E��z��Knѝr��ݮ���o�|������??�t��7��w~𭗮_�IN��o�n^�y�6��7�Ξ�|i��2a�z�y�lv{����ڊ;�e��,e>E�\���vܶ6-��k�Vo�t������'*���=v��u�E܋��n����R����������6�߾q��F���|n�k/y%ds|����u`8���⵫+��~��饜6{tvX��"�e'�F� �4d���J�K:����ݞ_B4W��ϭ?��+�.n��wr��G��_?��騼���Ug�Ne]P��ű��z�y���2�$�	3��k�'�x=����޾���޿ߩ�?���������?��k�"�7�0.0 ���l:�1�/�:YY	�ݻ��Se��,q�:���Č�3v!�_����l<�\�����r�q����aq�ya���[W�]��=�7,��N�{�=��Gz���uRH"��-���Z�n��25�h��4	����FA��ަ!+`Ŧ�&���AJTP�_rdX/�	�Vm�7�z$��&r��a�����e%�Z9����Ł%�)0���pF�䒹b�RV�H�tO�����-	�Q����+�Z����G���������ٹ�5���o�[����SG��/�ː��][�G���t��hׂ�ظ�����:�;����ow�o��~�I���r�/w����lX��?��^MfJ%'=�?0���/.�!l�ٞ��`(�FN�W��k%���f�Z ��J�1���lo��%*#l46�={�՞�����˭���Ň�Tc�Az��6��?����`�������Iݝ��icR�̼�����Kl9�yp���䙲�����\���&��-`��9�f��a|6���'���>8�̓���jo�܋u���֝�y��[�H�d)�'.`~�fz�j2w���"����ȁ��I[Y��R�E'J�=�!�Ha�r��`�	�a��Ԧ+}�F3zr�H*N�׊VH��S�iz�
���!`�+���G�
��	�FX:(�&T��Y~ʝx}$�x�H~��;�������[��&�X��F+$��Yꆜ�_�չ��
ئ�e�e)EEiOa�Y�z��c��S%�0�R�*̅�&�`����I���� ���� '  �	^ݎ�&W�A�\� ��']�̳�e��5I+!1Ql��!���		��L0��A�eM'
�r����/Y�!g��?�)Gdx̢r9�2���-6H��.$�L,�����ʃ��0�˕5K�i 3
�2���b��I�}�%Qx��8� �1�,��!p0�^��u?�Kx�����-���cVl����I��Ҧ��l�A��Ա�k��LQ;�Hh��%
��@C��l���Z��e61��Gz��b`�_<*�ЂU�P&H��_]�(�:�*N��Pũ�]C�5��FI���hbN��S����VB�I!�c,8"�a�(:�M �DR�Ux<2L_�b�0[}�T�*v��ѓ��x���6Hx��*a赩o&IH`6E^qVB8��W�?r
�G���L�tDh���;T�$�	fH��	���5ez�#Ob���I")�߄a3& d^�-�R`��q��PS�$#�;���y�Tv%�4�@
=Awx��f�v��O�ȉ6�ì5�i�T��lG��lS�k���rm��R�U�U�+隚��I�`i���Z5f���8=eK	�U�I�a�¾��Z)�����@�"!`�O��#J�"�A����fN�h��T�HB�^�d�P5O�h�Uƀ��� �QEɩscŁ�¨;y�@[�<�9e�֦�^6�j0�%&lM���ԣdF+=~��3T���V�-Z�Q��h1+a��� �5q"?9�����/zVU��9�����"�q�	���Z��2��Q Y��ŬSa!*���X+�b�h9cM�a��ᑋÝI��w;��=N�#cU0�7|��$ !P�k�,B��ƅ�Rh��O�T �4̅��"�O<9{t"�D�٦&h��,zY�V�Z60H _��U����Z�%uz�I6ң��	������+'���fz�[̩r�&	� �&H5Z��͘��10��!̙���
&��]��3�ܹ��L� ��-�
9��*]�:��hA	cb��`�$�	��,l��� L���$�ؔXa�/q� X�8�	&-R�A�)e��^2(4h�:9�-NT\#��N+B=���Dꀹv���t\s�	�%*� ���Cם=Gv\i�G "�Dn$E�d&I���*���ٔ�ʬ_��i��zk�z�n���X�$kIU%�[f��o@b 6����B�{�H��ǿ��������m�F؆�E��$@�%Di�
5G�\!��L`�hD�i ���L�˽N��#�)�&f[�|�c�Z3�UK�L`̓Iz��|�=)% ��x2�l�$��@L���/����ϊl�uA2��t���lJҮ�_)�X`C`��^�Bc q�l@�`��<�s$D�U�M��c����)ך��$J�Lf�d1�̗h�\�.�/��a�A�y��4'�EB�V���b�d�\K��YؐH\�4��3��	_"�H�,~� 0�7
<������pGFBH��aV���7QD.��9j
+��>��&]�Mz�8�HbH#�z��2�l���o8�)��f����.M=<~��I�T�k&����-�9=0���E�QЈ!�@Ra,�l�Ys~���
3!� ��xf��9�͚^MB����_�!�(�<�0B<������FI��Gh8|��߿o;P�+R��^3�
@S�� �ը��@��&]�
ۘ#��(�>�`���W���y�l�!���Uah���г�(��"0���Ԛhu��͛7�\�j�x���8/��B��f�������Ƨ'�<�)yΨ���>�y�N���xg�4b,&�%���V���xO}Hp�AG?hiu����~�Q:&���Ve���憔�7�/a�e��U�G�	[Y�ol<���x���t~0?X�1���)�JCϩ8����ݭ.�>��7�ﯞ���;^>��09:z���~��9�-�̝/��M{�2��y�խ˹�pb�ν�}�+�Wߒے�rZ�+��]sDzܯ,~�������R3/eW/.�C�������������n?���ً����g
�!��Sk�߄��n^��vy˳�K�Aoq�G������N݄�-��ƥյ��;�k�g7�_�"J!�}N��&��-q����������I.Ot��?ݜ���zӑ�h΀��Fc����=w3w�^]��-�<9i�g���ۚ�4��S[��Jyiq������C/�]쵹��Q79���7w��?8���V����>����{��Q�PY�K�ŵ�7�o=��湳LI���-�P/^\���6Y���巔�࠽z���Ԧ<���?��k��s�;嶷I���.�B��j�'�s���~wemu�
�Ŷ�5�����ƥ�����`��~{euc����|�~����MO0�p��ʷ4e,2��$�D��9<�NL�}�<5k��&��٨3k-�w��[���}���[�����C��X{�Ӗ oܸ��)H}��`�vB;RN�vBt�:�`ȹ�G#z:�����Ӑ��a|�������Č�k�.|���Y������/=������ߨ�U�����?�Ћp�_P�3B;�?%�
���O�B��`���;�۾�О��u��{w����O�������dxpx��O��C��'��Ȗ#NC6"E`�n�ɶI���gs��gs6GR��J�:]4�f�-0y�s\���~	�!C��D[�����uEF����=����|�1�N%\��ۑ\a��N	�SN������L����7"z1�㏆��E��)+����0�����L0;�ʹ���x��Q�I�����9(=��+%/_�`�r�ޒ*��紙B��ѹ���~vSJ=���j?�ܚ��;C�����<��ݬ{�6�|���͍�׏Z��.�4�����y��$��ށY�"��@���m-H>���3j���۷-n��%f0�6@��Ey�g,wǃ��Q�h�Iz���R�{O��M	�b=B�D(<S�yH�y6�d�Կ~�����z���F�t�;/��q�����ޏ_{��rJ����G����2�įT��|��Ҳyvʣ��`��RPy~�[���SBL��(�/GB��E�+I�~�h>?���=;�=�y���#yx�Iwi���mg}�����%�d�9/�a�`�H��V�4G�EE�K<�W�-7Eӿ�,�PifA��b�:�X��FI�A��0
Y��wQ&Wa�=���05u������ɸ��҂���Qҥ��.�0ը�0&�<9]z�(�0�f�e��� m֭ ����>��#M{�->��9~��y̝~���������6�/F��;�E<8�s��������hrz�׳"���l�Lb��F s��U���!%[��JH؜A]/� ��O>qh;��i�rı?¬(��FG]{��ݸ9B��f�eeBP�������܇o�jM���*�x� ����g�yGH���@J/�<=����)�� bSM��X�F
�iϱ�X��Т��(H$2v��&��ي0<�_5/2����B`�Q�R-��.u�߇���{{�jf��CI^R�i�lQшжLCV� ��(4�EE����B��T�KEk��F�6XJ�B_�J�\�	@-!4� 0!��Y꬇���z�Q�����B�a<�)>�&��)%f��_�]���Z*^0d4qW|����)%��,�Bw�6R2ApRI���.��� �a��CB��T0�B�ZWU���� Ԕ)�\�FV�@Sk�!ã֛���������2kj�F���P4cŐG����O`H4��v(ӫ&�e�.�����^y�	�I��&��,�S�xa�����cV��	��X�����X�?��LDNPf��b ^-��2��j$�sCC6S�jM�̩�8��<�J�vZ��ccTB����tN�0`��Q~2@��(	a�5���8a�*���W���8uY�1OHF!0Tj�X��R��Z�����������*�Q�Qlw`�3�� ��� �xW4u�	��Q�E�n�+�^Vd`Jg�m��qҧ�,r x�X�x�	d�KS���!	�q�_�T"�w������$dN���D͵��lhr5����Wmi��8�$B�
eVB]J�24zx�s0�䁠�7��,��hxL���%�-~�	0��é�>s�(et��86������'C��� ��X�|e�
+0��hF��p&Br��	�xD5Q)�ƠD�P���R�K��'!0������f����!��Pr$uj��j`hz�F͝P]4�Iߙ˒���0uF��b �a`�Qʑ���B)���9eǖ��@>M�$9�D���kƙ+x|dU���taHAB0^a�J����(�@Gڑ��r�ܲ�!�E�``"?�5�"�1~��� $rz�Dl�BF�A���H�m���3�OW�D��1T��}r�"d���x���;��1��&W�u�%�)�5��X	���?[�b�/<��b�����D�6 �0�0_�E�5f{����`p&x�cK�\-�ŠXlb��^�C�F$"���W��Li*�Iu��_sz�f�ۨ�l\p�����Rg�&`�<R
^����~�ea��ch�\0�S�5�d�.Hid����K`�Y�0.a��)����)z�	ƈ�-r��Id��/C�ũP���,,�\`  ��ʆ� 6
�P	�;���C��( R�`@�$��QA:��˟��#Hcѥ&CJ���	LI�.����#J����v�~y���(4h�g��*��r�eR���`4���A�V��o�4����k5�8�X~FDo��c堥wDp���+�F''@bNf�L�. ���F1�:/��Q�k"|�w�q��3��K¥Z�H�j̚bF�q!�.�JRD�� Ȓ/-)����`h�cV��`좕�۷o�A#��i�0�Uit�ăP�<1����o�J�&Y�B�P���5<��_��������7ߵ@}�t�3��?���{Be�OO|T�Z�E�(ν�ӽ'�+s�����<�Y>���!9$˺��d���;�N-�v�W~l��'���:^��g<%{Ǉ{O>���������,���.��������o�N[K�Kk��ƕ����������#�I��Μ_,I�w�=��Ξ��}�'��.}t�����G�����\G�e��֓��VɃ;�n읍f��}咵˾����ȥ��"9.�S6C������7���@�r�(�G7'��_.��U�x9�{4=[�Gc=
�zy����t\����9���.�����R/.,�����{ey}�mei�����KS��i�6��+�m]��Ǝ���cwwg�+^2��&���7PV�[�s��~�{}�Nz�������1�Q從�sGg����>�x�\oi��N�@���	��O���/[���+�������V�7.��.�m�V�_P�9;<?��������p������޺�����������;�w��Ov�\����卵e���أ��/�[��������?>�����Y��˧������V��n��g�,=*�r��-t�1k3�@�_������{�ğ���_��;:Z][��m�ӝ,N����p�qw�]�ŏ?��:*��=|:.����2꺬=8}6�k����wO�N����k��q��#�QKBxrn�r,�:1v���W�B���/��??9��/����w�/]��:߻��qg�C��o���?����_W��?�������������N('Pa8�Ԛ�G�d9@D���s�%[`<n1Z?��O����9O}��Θ�Ë�Įb�ѵ��ϋ3�;wX!�#C��s��|��W�ы���s��<�e�vf��N�D�����ւ{��A��?{��?�^�vin�>=:��N�<�=�bj�`v-���k�d���H�d��d�$����Ef�^� 0AR!�E��y����t!A�0 �}^�0����o�Л)EN���(�@�V��I��-ߙW�{,�{ �!C����]#`�4� �D�I�dz�u��    IDATEa��}q��e[���3��r�����M�Vgq������u9�����פ��en�W+x/Ƚ<�����܃�s^�<�zs���#��;^���������ܥ���,���O?[��?>>���?��Yw6��[���r��U��A��0���Ȁ�9|Y@Z�?G� �^�ϋ���\����6�"Q2@�=N+[���]�	�|��%�`>�[�>	�oN�
η�~;���_���}����.y��=�n�8��s���4w.����ѣ�g'~�z�K?�G��L�^�ә󧬧/ϼJ��B�u< [>�A��`�����s��=�ۚ��>�;:��쟏Nv���?|�<�u��m;���>S��/�Lrs:��N�Y�jM�"�x@��Y��U�`%���ɳI�4l��"(���,��a,�Y�L Ք)��d�x�Ѥ���	�a��mlu)��U��8����e�Y'��`	)~�t�*̩�Ro�j��o��������GA�)��X�T� 2��S�3{�-¡�&�}��E��ʖ4���,fJVd;�C�H&�x�Ǉ{G�����d����j�Cr���#4�"6��#O����AvR��kt~�.��Ëө�GpA�Q��El����oC�F��'1���#�;~$l�������H�Qĵq���5O��E*���y� B��Ji"�`5!��;E�j9�R�p�P+���t}���o�6�Y�)X�F%�̋h�����L�IG��ƣ�J���#�٠h0�p ��nݲ:���@���KT̹��gh0b���sgR$�`u�)0|��{�yx2����̤�M�d��Qû���T�i�⑌�&���@�I�fY�$8��3Lll�K�A�'r���Ia�� �J	�bWd�.5[^�4��"��6b�(6�rcEfH���f�Q��.�Y�0�e"��GVg���@�����^]1'� p�T=pb +�õdr�<���m�S0��FЋ$�Q&��-r��1�4���2���WZ ��7�	C�9Ȫa�d�C3$1Qӄ&�8i�
Mh�
 `]0�3@^��ɌSƖ��C��C_������5M0̦�S����C�����%B��Iu�bC���ܑ��$���$����1�k2���	3M�f�dBl�1���h�a���fjJ�"�X��W<��k`�(��Lp�Te�]`q�&�ɼ��L�O�1�ԋ?]5�tQ�K��FI؉��7�x��0�J�Ҟ̣^`5@0�b��$$�h0�P�R75Zu��4�/���C� Մ^I<IK 0�	#!�$�R>�:'� �J��!=���fJ+,	ԕ�QCr�_{	��e�\�f�0X���	N�V�4��G&�B�=C�g�h*���@�ćJ���`0HN�0!P�G��I�.�^��x�aP����[!�4�^~c�	G�Ü��1B&�x�$��$KTrKH��J�S�S�ܙ4]2 N]��A$�ؘ$	bP#�R�,�C�
���X4aH/}F�Zo���VH��R���`�3p�$}�iـa�F�~]�D�YW��GZh�+��\ZI`�h��S�8¯��,cx�;.�� �G�b�FX3LH]���!/$$'�`�T+���bH�s�!aT=$]�����\�<"tPcV �V�M����\`h0��.BT��|�L��*�E�L��O��Ê-�^_0��; �1��Кx_���d���1�	����8	 ���`Hf��#T.�[J<�+l���3_ �Ԛ���"�q�+��
L�2��4�ΐkBҤ`F�V���R�/����C��J#�ŏ�P��T
w]<�v��N�..�"��E`Ν.S�Pa��-�z1�ý�%���63 l]AF�D�j%̬�����K����4̉ʐy���q)\гե��������u�Z*�8}F�od�ʸ����#r^❀�_��s����B ]�ӟ��5y���;�H��-NMWQ2}���0!(�I~��p
0_�l��#ݍ��蒮FFNl���S��&ȥT��]�X	^�b��1@B�%�ʟ�g.*E��+�6�j�1:iANVooo�u��}������'.͑{�.2ۃ[����s=]�g��������vgAn'�*���d�4���b$݇���}O1z�, ������^q륵���f�Nya���s�������	���&�Ý��_�_�r���o�_���E��^�OΟ��[�/��uyރ�����������9*G^�;�Z�\����oO�Ϯ;���z�3�|[�ެ}l��4�wў�{b�(�c_J:.���^]{??��]��	7a�.��s��cj�'�G9=�b��Y�.K��}DO�(2�.O~�=Ձ��ƓSo�{��?X^��x�������{'�����m]�����2N��s9:t�u�zecuc�$L��d��/�m]^��=?]jt>�xQ�.75��|���+�6wV=�Ꝺ�"�2G/VvY=7/k̈́z@���0��7��7/9۵:^j�Αy]�S�w~�/���2���>敍u��o��yѴ�ˣ�{�;_�yp��[׮��օso~��ѭG���yHqnimqy���ʲc����{O�=]^^���Jo����I��\Y>>�w�������Boe}e�LnI������ͬ�f�X9Yw�~�$��.5��B���ۭ���n��ޕ���\�F��u�=�ǎ��Zc��ͬ�ߋ-G�~�t<*'���Y>�w��������M?��٬�?������O��-xk���bVK�����Y]�b�BXYo���q*B�۞۳���d�b^k���~���{�]�}����l}m�;X����-��&�羴����v5�S[��X;�
�,i��;�PfRg���윾�˶��0����6(NW�n޼i?��%�7y�����d���l\��k��f�'p�SN0�6y��O
��s�R���ɾ���;���]�裏�}����ݛ�wG���^�����ړ���Ω�C�h��i9ۺ�iO��8��A�\`��,��l6y��ѥ��I#�&�#e0a�,�9��nhʇ���c���_XrKV��\�!�2�x<���m>#䙡Ӎ^B�#lY���	��gM@�8����`��3L!��!X�#�� ���fx颌��{:��; j�0>31��O�/]r̞.�N{-{[���{Z�
�X�/�8Ku}�3u�Y��{�*��v�~o(|�L���^#��7�ۘތ��ho⇕�ks˫_�h����;�<����Ү7���{>�����u��7�����z�W�}׉�po�΃{~��@|n{���B�W>❖Wk�}[A~(2�����l�ʒ$K�iH�KN��ֽR1���:I[�Ϟ�E��uf�3r��7~�I)�������������h��r�_<1�^�蓏o��F�MMgj;��������HN��~��m&��o ��A9�ݐ��c̦�*�y���A�
I��s}��}~��Ps�d�9����=k������W���Rv^'��v˧<_�qPg◜Y9B���F����U녹��R4 0�9ׅ�9���&�4cN�i�$9���	3=@����#$���*��z��� �!�r�`�:�k�Zu"�"���*+��I2FC�!-@¦! X`��`���x�ݲ�nm�l)S�c���*a���B���̑��_��Hl1;"�SY%Xɶ*Nm��1J�5�r��]��K�����+����p���41s��Gj��I0b����z%��R �����A E�z�BZ̺ ��w1���N9����.��d�teԒ�p-$��%$J`Is�	�F�N��wIs������&�\��$�H���L��	!Y��P)8)Q	�|YW.�
,.�T�9���`64rţH�����zm����qg��́���_� @�G��"	��!(Ltf��I��@����l
 '��Wr�m2�&���W���jJ�4%@M�A��W�(F��LI>3�4�`B9ލ�%�r��H!yS� �(�$�M��j*�a S
>�07v/m���0u�����pU�Md�00�T�C�*�ф�^-u� ��@�9!$�Lãf��
�ZW1~u�i���ĩ��<DC �0O��P�BͶ�9+H��]��r�Q���7��H�"�-d�	 4�$]!T)������f�1�2��#�J`�����>�9!�a�$���d8�qJH/Bj��fho�P�pQ���qZ��	/iҐ!	�h&�5��4���j��E<�L=Y�j��渋\�2�Q�_�h��В��	�,u��A�9� ӕ^r��d���be�v0r
�Wb�`<%+�J �v�Bȫ�+�Sg��qCr�$\�'�uENV�)�$ȰŅZ��1Cj&�a�C�+�j<��U�4C�d/�	@o������E�Vb%L���k3r�Qg���jE��\z�W�~&�dV��Fb���8ab$9�V�`�D�H��d1�/��l��U��p��97T�@ �R0ĖSTi�� b��4/�c�����C��қ�(	H(�N�4#' �����3]L 1�R��9����a��[�*�!�J9����T6�`�M`��x�=L�t)q�o���T[��� xl>IVr�ڼ��)N��LI��X�EH�А�ĦY\1�.u�◭&Y!3�&��[l��$60ᱢ$��Z~J���*,$	�>��J���ʐ�t�	#9l,���I��Tfhj� ���r��SV*Br��kГS�'[�}��&
��LfX��I/Nq���d]J��I���,< ���M`���T����:gi"�3Yу	���A"Il1W��Jl��"J ��%+iD��G���R/*`z�8U+ 
Zx�B�DM6|���LJC��sx��x���DEC�g-͚s����x�ߺ62������+#�ָ��!��Uz�Z���*E��Q�U���V����  ���b�^͸H�/ٛ��(hC���%-zAR��$<+��^k&r5�u��3 91'NM�R�	�v��k�q��?3�����;*M�(W.���g�{ｇ!C&Q�b�!�P�l���I%׫�u_��z�h,*a���Z��~����K�����˃2���fU� ��qɁc�E��=[QY���WEJ\|n�/W�ǧ�%3�	F/`=�j&c��Y�C��Y"��罿tlc��'���S6�Nk�|~�3:�'����]�u6��=7�q�����rs�U���r�x���w��+�ք;�~*ڳ}ӣ�d=��ݲ�`r����'��^�
.��g��ã��t6���g��u�3k�m��d8�ݲ*���3��L���Zl��<5�gy,��VѸ�*V�32�N��~"r��]{�ַn�����|<��٢ŭ��A�����V�yg��z��6��6/]]Y^󼧬���<4k������Vg������?q���m��3_e����f��I��.�{�]n����Ɠ��NaW��SS�RG2]�<��w�������n"�\�>�?oM�M^4��Ϗ֯�c����:_�|e������~�rkΏߵ�V�77V���W6/{M���s�[��kK����H�3��~���^�������^_�G^;n�;͜�iv��W��-[����Ȃ?�df�u���ݏrs�5<�X�v���u��;�y�Y\���Ƶ|���B�?hM�'�K]��dYq�z�,%A�t��o����M��Z���^����w��=8��o��_�;$����hpؚwkD����3GSVks~ɚq��r��K�ݑgS�ݓٴ����37e>�����O��/O��c�s���B�˗ʫ�vv���\*<9)���-ظ� �UP�پ� ����m�E6׍�gq���Ke�߿okr��ɛ7o��2Z�`�4��\lDbK�w�-	 5�{��P�P]|	��m�����?{��?�����?��G��+������M���g��;<?8}I�&�N�g�ʛ���&�8�Z- �o9 _}�=|��W{>@��d����J��=g�U���������OV��P�������u	L� ��S�#d]�l����S����s1A!�(,���8*��2��[���ƌ��30,d/��3f�,��� �D��'�Oy��o���ˎ]~���P�eq��S~Uy�
���򕄳�Y�x�yu4z^�%%MO<����T:�P��[R��Z[8X�C��G/M������W�{��ő�=�|iqtޞ�-�q��n����hqr<<��sK����⻉M_�!�t�1 2��	��Dkt�l�lP6�f����euk��rwVF�����Z].?�t?̤x�;����ɉ����OG%^�������O׶�S�g�k�n=��>�Z��%"_h�<ooVy�p�d�3P��L�q�d����?�ܬ���J*;oy����d�����Н���^|}��͝�tqu��m�
Th^E�,��.˃�,z�X ����+�
�Y�'@IK��3��� �mGx���$�f�M�W�gBH��S2�W�%��j�T��)��aքOl��
���%�F�4�)Zc49TC��ӻ�c�ƅ�pꍌ��F!�e�P3d�s��E�B
�!�tY�>bz��.��FH�ܾ�����}Wԉ����H[jAr��=��A�D��7q�u��c���q�S+A�GT��:p(���`\j�x�Kf��"H���:!	;Ǭs�A�j(08CIH�p�-��;�����8V4�W����5m�Ð��$H����#�;%��o�l)��̢5(�!T�H5	�L��8����O����Eb����&F/W�b+�H��i�M�̝H���_��_�1x
��ƫ��K���u��#��Z��|��W�F!lc4j�*�7��Q��M�GHj�,`rL"���d��`�Ԕ1�a%Zr@�jzd4x�B��>s��ɔ`&є��`�4�-pB� �&zȔ4�
p�ѐ	"ɸ�J��3��`bK�E�!�ؚ8��Ef]J��IVk2$���I�q���*r���� �6� 0MB\�K�Zo"9 ��o��ٹh�Y]$x���ǆ6Ck��y4��I���p�!����&H�OX�e2Y��⺦"�Z.ƏV�	�	I3<I;ZVBJ�Z��
9C#��$(3���	8+�Umr� A3QqG�	!r�(5�#ċ��[��%��Cd�_t@h�)i��!Z]��IH�a]��OO�a4jGP0��*�IH� k�Ȕ��?|�g�K]9	i^�-�8*����Ey +Cz�,6���L[TqG!�L7�&��h�R�	���FW�0g�+��JX��ti�PG��ɀM�d8G_��x�9�V%YW4��]|���KH���T�.��7���t"k�J�d�;��^��D��X�&͗�柋����D芦����` �e�I&<�B S�KoHb��m
}��I41��>�!�Iਚǩ&�X�bUe�ڬ.�Z B�@��J�a3�Z�]�R9}m�T�^3VU��q�I����{�H t���F3A�\͜�.M��l�d�
 ���Y�Q&H�I�&�E0XJ�������=|��JI`l�+$d&�c�Nx�uQ#|����7���kf�a�WCB�6M l���D�v0�xh VJ�!�M/!$����$+a�B� �H^3�O�`��ȉ�P�f�� �;M2d��-M�Y���!�	�6	��$MS��G�.M�!s�&$�/�4/O����e����Iژh&c����J�#�� Ù ȉ'َ,����+͜}�6�a�PK�zS`Вņ� ~�^�YCI�f�bC����Üa�$(aS�Jf���ԅJ�-�����E�  8Q��F���O��B��Q���,���F�Z�Jc_��E�@J&�4 ��Gɞ^B��+� k�!�E���b��1V81P&r�I�R�*]Lz����� c�W�y�i`�����5C�yc���	i�����4L 	J��Cc��BN  ���k̔�)���᪫c��    IDAT���sC�RL��>�}�!�o�+1���}<�%閙�r���WG��$��_Ԯ#Ϲ�A)�p�/�I�$�>�usk�uc�s�t2��&Ѿ�I�wМ{I޳���W��;<������K��W�������p��:/Z]�[�0�G0'�3����ʞ�:�k��O���/G�������������4��Q<�,�ng�S:�E��:!���Y)��6�-ޑθ������c��0s��B3<O�H�On��v�-��ٵ̤^�)
��=��ag~u��|��:q+��������������W��i���n���k+E&ȃ����'-q��Q�wt��β�����q��I��5h�v����ø.%Y3�A�0�?Ҍ���V�x��|��;i}� �v�k]�gg��Κ��.��p�{a����W������u�����Ks�AQZ�]�n�S�~4�Tx�g�7��ݍ���?��>>z�x�Fg�2i/�NΎ|dtbΚ]���Շ����h�Y�r���*��;[�q~|�+�+~��![���Y�ٞ��fÓ��q9�ݵ�+	��{>��2(��[s�nzzr�B���}�%�_���֣���{��<���_����O���6�Yۉˍ��S�	*s��b�_���u���:q���	���(?(��|�<!�_�|�悇���}���|\@���z�t:v�����u�v=zbݺ2ɗiʕR�M����,����������.9fIxr����_~��W.rnoo[�6
x��xU��ȿ���s�WB�`.Һ���US�3=���䘝�%GOZ��
�\�����/�;Mqm�~����7?�×��ڵ��}�͝�>޹㐾1���W�7/_������^�����+�v�ۋ�M�'��l� '@ؿ��c��8/��ȳ��7ƿ/Ϗb3Y���h�j�����b��k���+���.~�F�!̚��X9�(M�s��M `&Z2s8��ˌĕeŀ��`Q2�Ժ��m��ХF�S�AO��.3��@S�zK���]*_p��>}�:X\ű���M��ݳD;�!��/9Kq�!M[Jy�����=G�!V����;��:޵�Ń#�h�����}R�.�)ν9{��W6�vo�����|k���i�m�����_<�+�M��X��==]�I���휾��M_tΖO�}3v1��2��wo򅓮'��3���9����P]����kWG�'Jɗ"��۵�g���?��W� ��z|�����~_=־�ܞ��u��������-{��;�����s���{Ϝ��w:�D�㗹���Z��M3��on���'c���,/ '����	�]��:;?����#�d�|���γ��٥݅����d4�v �F��i��/�Ҽ�$�yS�B�Đ/K��C_Fs�	�.�a��f
(����/�4c,{X-�h���Y��)٢�Y�U� �"`NS�IF�&}j��P���^CR�0�4vR���1��FF"Na|�e��70�K�ÓwͰqD@�؝ݛDB�����aӋ���dྠ&�8��%��nbFe��=�
B�w�y��=��ʏ�.��8����|�7
$�T�:�������t��N���:a�Ȳʏ��A�W7��;'9��,s�7�$��jԎV7�d��)Q�&xyp.�Q'��Er��=��ѹA(CkFP��y"t�Ј�S'�b�H/6�V��;V��ݘ�J � X T�o<�T˛bP�lş�x�h��AX<8)y���&�H���V�b6GH���-��}�0����0B�K�.T
<�nI�H��a
R���N�;� v`�9���S����}���ka�ͯ�T�G��3��T+<*rC R�7�  s� Ĝ#x�jE�x��+!'��k2gϐF�!P�3���ׅ2��)%CE%2z�j���_��cLj�6�^��X�x ��#ASf�F�+zB�����S��2��u��
w����r$�1�EP� $�:��'�0W�Ũ�!%T �.�4+8<��' �
�	@Z���X��a�$�O�>��I&�E|���*4j�&͋V4��'L�����
�-�Z�>]a���.���XX�g\�4aj��.$��F� �#`r��0VL�ɯԅ�L�Ae����a%�0�3�+�J�L�l�i�h��5+sS�	gL�,̚z���Ҙ�� �C��DM��N53�ф!`E�f�3L�z�2�̙Dn�K`05{�K���" (��ÙZ<a�L 0�B+ %�Ր@�Z�t	,�
9�&uƛ0����@S����uxB�ZS��	0	8��a�����CV��D��������p�|��M��Z%���ᑜXi^,�ŗ�P���@�R`j㥂�G02�J<C&�+m�..t9r&fJ#�G��!]�N]&HW�1��	��/u����R�J�$�E��KM)��<��(�K�&�1O�	 Mr�E`u�]`4	L]�q�J�4JHB��	%YaN·"2+JH%��;��z�3M� .j�O] U���hV�EG�� �D��Y�d��$H�:Ïw�X��&�$�m0ibH0��|�DV�U��[!�'�aN�&%9 $�^9G�^r�	3�.ulu�9x��*��B�d}�!u����� 0$['�D�'$�~��	9#�kM �R]c&���	s�x�5cN&Se�U�&�� TL"��FMcPJ��8A�k��� $���,��&0�B��)�P�5��0<]8���kM�m8aR�ȱ�L����
N0�6��|���(�[9��G�V$Y'���cG���(��� (5H�(��m��$�����0V��i4d��G�R�Tk�E+��'�i�2��T<+��b[{���2uO��7�qƑ�b�A���l�1Q�#�E�QSfP�s2����� ���@�J!�7�[����q��{1B�J�1��Z}���hpғ�����T����J�K�۸���g�:8u�@qy�K-]p�n���L<=X��y��������X����� ���E�w�&哵�6~5����������r��ehO1v{���ڸt�^�����q����{���<yﺷ��8f}zt������K��{ώ=�����
����~��/'�T�f�?����av~6���}o��3�^�v6:^h�y��un�ϧ�Z�PP�0Y曵��~��t.����)��$���⛧]hm;T��W�i�3?�ZQ��r��w�}改���k��9�˅�r�'?$�Z�|kz2{>�=�������[��������K���������]�.�at��d��^fk*�U?9/ǵ+�mo�u�ᩥ��do���Yw-_-�[~��.Ŋ�S���_��T����WA]d�$�u���=�\�E퓝\�����;���ڽ�E��lY3O�zǷ[n̽'ֳ�ዃ��{~6j؞;�ߵ��^��C�Y��V�=힝NNٖ<�^i��C���;����Ȼ���mΣ�_�h60�垤�)u�f�J�����u��aO�Z�9d��ݛfY�N��9����2���ɱ����t���_~��ɾѽ~u���L�1�ߜ.�ƻ����)��HtY/�i�@v �s<r��u�	�e�QAOWͺ���_8=_*/v^ڸ�%��K��O�����L�K��K;Xx��7��}w�߼{ ��\�	��کA�.�j>x���Q�_�[*�V������"�����ʡ�B�}���/~��1]Ք(���5N���4����5+�X]ބ��0s)XM�K ;�v���K��t���w��zeu�����'�lZy|n|�h��`}���3�(�������OO|Di��/8˩���O�Oڃ2��'��`���K�QЧ��o�d�dBx�t�B�а�! �R�I8&%�L��k����O���Ht�3���L	 �pg{{Ȭ�$�f%���0s�(�Q���{[�hjg���Y��.
}�D&b_p�m8>y��~:��tpޟ�z"�fc��F��"S�A���9tMo��/��m��Wb���V� ��	��_�Ι�<;M�zNx:^-?��_r�{�}y~�?ϭ<ۺ�����:�Z�;g�aǏA��W���`�	�_Lڣ�cϿ���\���ăD僚���7���7Ml{xx쨐m�vԁ�mm��%ۙ]9p�<~�H-W�����h��.��@�������:t�f�'G���ӳ�ѥ�-�����˗^�˟�o���F��b���6�agro���S�d����;��k8e�.�a��Hy��Ta[c�g�7FϠ;��E,	 K����h��(7�ϽI`8rk�`wttp䀘_�a�d���x�3�t��ERxi&��L�t�e}q�QXr�����P�Ȩ�Y�ѫ!�1�\W�f��J\��3C΂���ӱ�,�	��(2�Ew0��5	f� �0�\Є\B �Sm�P�J�	2���/j0	�!��N!��6;l��y��~����?���Vnb�
^m+w�/.�X[^� q:U��y$��q㆛|���(���N��i#���w��x��x
�����i F
��/� ;Lp:�1	���)��V�e��@자n�	���R��^���OOy��	wf��+斞.�4�H|¦���I���<��*i�M^��a/$I3(`a�<_��ىa6������Vb�9�"f/�2�m��+�Ί_�����߻w��Tn��h�Px��2�.����?��S���5M�c\nc'�9r�ɤ�)M.�}�0M��Fd����n�@CV�G�e������C�2zV�ѓE=�&��Y�L���P&<� ��������^�������a%��Q�<�r(!zc�l�s����9BJr��kJ�l�H/wf'1ǋ��&�U8ҥ)05N�O�" �FA��,'Vр�qj�6B�z5z��V3M���y��iL�f�&�$<�G 85Io�Qj��U���
��Jo����Jf�dE/+��B�K�4
e�IW�?՚�%X��@&d����W#��xh���4J&(.$V/�@)6���$���l 	� x�EP�� 
�I�as��"���3($1�$4�U!�p�͐F��F����T+0�ɀ&�b��e"�I��e6L��xd}4	 .��0�d�ş�6��$C &MP��V}ч'�Q�+xp2��hԡ�2$q�#�:*���� 1'�04qWà�}� �WYa�h�p�JoE�2�oQ	# ���YB�B��^I$q��+�2���`�~����
�&]�@8��0&P&� �%�+�D0Yo��6`�ę�%�0�ECX9#�����Ye߆ׅ�xP)0�a�p�f�5� 5k�	 �.zul��R���֮ c Y��F~]`d��k��5�ij�1�Umx.z$�]΃r�$L]�h\t��06�!d�c�,��ԛ�hB*2!<�آ��'׃FS��I�	  �Nl!�F�X�;�  	`h�Gd]���q��^SːӬy�_Mz���%y�0�`%Mj��5ßH4rjx%Ni���^B49��Fm0)I�^^��0��7�.�0$���T@�4i�X�xg� D��X%���TbH�S	���K�2�4�2�I�ESa����)��DN��"��\G S��EO`\���QdjTq�l��$���*T�)�ʫVq�Q����C�q�
�"i��s ����ǅ:����
�!MC�5���,\�<��m�����K3��/0Z�\�MT�
X����J�M�Q�a��$.
K�@LP)xt�g�cHe�����4���
>V!ץD��^9aK�0r��U�g���)�(�2k�2�V�[����q�f��ǻ��KMs�
����!|��D���b�WB�5��&x��"$���
!	R}��$3�&��`h	�J�'Xo&=�j�FT�� �/T�'��a&�3Ș��p].��g>����	L|.rA��5_�?�_n^���F/�{�����>U775-��˵Β��ei z\H]\jyz�xh<gVR���n�Ev;ѕ�r]�<Z���Ci����O���<�;���w�=�;���GG����q�3���������l�|������N�x�5�rOs��6���5�x�jI��X�k�n�|���f�:-O��"�A�a�*7���'��;������]۬��~�џ��oN��	�b�ePrB4GHK�1W'n�xۡk�J��L	֠���e���W�{���
s�w3��l��b��2��B=Y�-]�w���{ǯ_�^]�/�i�M����]��jnʵk����a��Z�- ���S �fɹP��y/�/�=niC_Zr��l��%?��U��׼<�Qy���-t� �<��*	�M���jI���-?'t�~�������"��b����}�����;����do�I��&�������x�������Gϼ���γ�^gx4l�z��E�=.4�����gY$Wz�^��yu�J���wU��`��yd��%'�S^E�\-��W�2Y�%?�a���h�e�
�d��ky�ť��syy���ϻg���7����Ey���t��w��mK�Y�g͌����ʺjv����3\<5��S�a�L�:q����>�L�����+����<�<��{�b�C��坵����(�=<~��(ʮR�@(7��j�|��w��׿�5�V��&m4�t�����]���Y�D�{d7s�ٳ��>�b�p���W_��ɩT���`�n���o~Ö;$"q���c��4�6�&���A.e{#��/���s�����[��6�4�+�L�_��[ooˤ�y�����l�`t#7�g4��F/�z�l���v'�uQ�Le�6a2��)[��J�:���	4 ��Z3����%���U�Ss��I�fl��H��P��&��}zuᇏ!�,����.)C���O�2R�k�/����a��s�7�dA[��\�KS���|u�J�>3+]`��Mrnv|�$�+��^ߗ&��z�E�ܹ��ak+�O�GI���~����"�)�zJ�ɼj�̐$3:��x�{�3�%��O��W���^(?[�I�vk}n���o�������Ŏ7 �tO����W��Gӹg;�^��>>�zV��6֗ˍ�ӡ�4z��1-5�dl��%�آ�GQ�s!�%wK�1�dI6����N�t��w��JW�]���������n{u����A̓��a�����2��Άg��O~��.�_-�xy����k���O�i���@�q��mY/"/��r�*ӧǙ(kH�Y�L��5�b���^�ʹ����۫��~|�{z0�œ�7;�ݥ���I�3��8�p�(^�ԅ�w�L��R��&�'��^&�H�e[]�	���j�zC��zP  k�;zHJ��ę١d�-�r�U4�D�Q�, ӭ	 ��G�����m�%@�R|���	�
/�����"W�.&� 	m�a�-cK7�z�)��;w���h�vG��֋Tx�s�;r5���H�"�k�Ѕ�m0a��0�x�_��/�q!��;dn���.��X��0��ơ�����9]��L�5� � �$�h5��_9Z��ũ��S̘�]���v��/����q��)60�� ����D�N���,c&5{����/��i0
JTE���ԲGc��kvȒ�W���A�642�$�L�noo@�l��Y^蝼� t "�4>48��JB���к�i�
0��N��J)E�	rC�+�)x_wd)2p�)r!���+Tz_B����
-�S�ZSW��Fw��Ԑ�5��;HxMJ�<���� 5ENMz&f�>�lyӤ��F�M�|��kz0� ̻ڬ�/�`� �� �QY̺�4���
$���(	�j]�jV�JlQ���7V�+�.C�z��t��U�e�k&EBB�i
����N��I?<N5e� Oom �=�.M�d���4	)<Ѩã��0�$���pA8B��$�h��A-��� 0��9�-�(H��N���}��J�
�N��Wa���������xH���	C���Q��(��1.���!(�j�B^�_e�I=$�DHI�T�bB��,� )�m�«ٌ-���!}��0 T�Sy�I��V%Ø $(�`�1�4�    IDAT^(��JR#�^M/���J̈́m�i�%����2T ��q�V�Q��!CH	�h6��'�$��W���-��LHH �D�&�`0J0z	\ �@�0��� 1�>r�`8��޸Ќ�:�\�a�ԕ��j�#oॊ�^���Gl񮋠�b�T�i��\@V!�Q���[�tUs��V�M0�m��� '���N$q�� ��N�q�^r��&@�f]�J%D+��a��"a��`)aR���AS�@ʿm\�-�?>!5�%�(SScK&+X<2�^ ��C<hɉLx�C�AS�Im�K��`B��G��(�4���sF�Ø$��Ӱ[B�̊�	$�ꑉ"B��!�eË� �
�|� ãI}4|Q�A���	�4aM���+]�M�O��m��ܦ 
㫩'��W�z㝒��"�T�ҥ!+d5��&MF�)����CL/B��Xer�æV4k�ĦV����x�5 r��#r�	5����LθP))��GO`d-M
JrH�� �	�>����Ll4\�@2���&�	�̅ᡌ#d ߒ)c�-]�1ghvX�z���DN�D	�&������+zVdJH3����Vx�KI�!0!O�4a��o�.N�]�/�?Y�&�	I3��J�4�_�@�1M�"0��	[lA�|]L��e{ITY `J��I��0u\�/L��N��D�$��G���FSja�i��uFbBCP*O�u1	>�P�*"����KH"h�7��!�yx�Q�^�C5��� d�zq~�J�C��*9C����`�V���c�ڈ_�(�"~�N���I��*C�j�(/����ӱ�=���Ng�:�T8U|4�}��`y�ut�^Uy��˗��x⁶���n�s�������\�X����-�߹�Z��w�38��#���]������ѽ����s�h�#��d4l��\L���̓������ɻ׶֗�,O���-��;|��G�e�l�V{�1��ʟl-߂_�X\{���q>Wi]Vp��q3��aGwIǓ�nٝ&���"y��y��)^�9q��R�~�����Ξ$��3�GDƖ�{f��*���6R�$k�Y[��a��C=��͋�l�8���(��A��R��ʬ-����Ȍm~׿*W���pq���ι�_���^&�ᑥ�u��T���0��E�Оͬ��dߍh����3�w���/��΅�.�����O���t�w5�^���k��������h��]Yj����=�N�������d���,��V͜R"���;M��m���#�=7�����f�_����]^�h\�����!���Yoۉqa�a���{ٝ�=�鋤�'ψ�x�U�>�i��C=c����X��l������o�Gǿ��?��ӫg����7�ͅ�����;��v����������c�vـ.����X�d۞.���$eʠ�uI���~"�}zIWW[���P+�V�r�W��2?=����q�ܮ,y�R'����+���Vo/my�7�;ӻ|Ъsz>�s5y�J۫o� �p[��м� �/Q"{7���+�r�����|�v`��+��;�7<�����������O�v��=������ޝk&�~��E?�m�����n�Q�� ݗ�>�K3���K�@�F�[�V3�[�_|�[�v즷���+���-��FQ��P���c�;���\Hjݽ��6�y���O�d��_�����W�e{�����<�e�m��������ܿ{��_r��~ó�����b`��u�-�t��2�y�FCP����ZR�U�ݩM$��5	9Tj��񰢗��&���Zx9�\B%0B.xa@�SF���I0�����F0M��t�L���m�ӭR��~�hD���hB�QEF*�(i�0�0QK�GQJ#itmM�#&��H(7��0w�Ó�/����k�������=�rIU�.�7� ���_.J�HPyݰ�&��g��Ѵ�A�e1�F��������ō�[�J��F�w�����/z��[�������[�ݓs;+�*ga�����ysu`�*���5�.'k�[[7��{Й����	�<h�R^�������YZ^v�P�r��Tž`�u����s�Al����{F��֦�<����=��ݻ��积�k�˟T\�:}�����k�n:�U��6'/�'Ϧv����g�n��_��=���a�^:�4����ә�_�]��8Z��o����/�]����`T65g�����?l����/������t㚵��-��w����輗+��rr=�2�iR!�c[�O��
�\ҟ�4)�Дc��9[ 	ah�3�J���*�aN+�2o+���\c  g. ���8MH0$0�$H�d����7=(Q�8����_0��+��f��%+�*�+`x�r$�LÝ\�&��[�)V��Q	^.Ye�"0A΅��:`��g���v��N � qJ�y�8y �ٳg\���$1�R%0<`��⌢hA{����[�,B�4NW�Q���G՝�4߾�}J� �1���VlbN��V� �����]C�U����ņJ`��E����aj0a�* �'X���*0�l\�@�Ɗ!A�N�\3R4Ω�V�CO��-B�.�lEk�;U�)�t� �-�#AH�oF<�����t�d��-�O�<����G��o��o��&����`\"��J<�Lt[1�u���3�U���M3�lٴ������$Ns^$��W��$�!`��g�ФȄ C9 @bP���ѽ�R�F�wI<�I���%WK�\\���ur��|a�N$r��5Yd2�b�.�_H&�H��h��-���鹠p`�U4j`BCN�d)MॶuȄS�j����a*��Z��	� Z��d��Y�i�*)� �a�(�\H�����n��(J��`�4Oo�Jj��\�5�^��!�T����vV �ژ�Cc���CgUR����r�M=8�)�BE\�ф!!��Z"��!QL�i2�� 0K�:� ���J�B-+� x$VU��*e�)�)���a�"��� �89����4��&`�@��#��U �i�LC9�� �^bRwQNH.䙷� �J"K�a����5�9���AN��"ș��Gj�i�4��Ǒ<T���rI-w 4ROd �?<0MB��T$�Vma�]��ETR�(QVV��i>��E�*�k I 0|�(W�DG��S�%�ؘ�����P���$V��M0�����E� ��)��LN�r�T����>�#��3����$xBT���8#���Z��OYX%`E�!I��"�����J�/�Ȋj%�aa���"�y�h����a�Ǒ����m�xUVgvw����e��kG�鳴�$����Ti��B������
�d񈄬c���� + �0���i���$�Z=	L�Kl̅D����w�h��g+��6l�+��Wh�SF��q��*B�i>[�r��-�G�t[BXFA`y�1D�0�j��2��h!CB���j<��@0r���VH�1/6�j��-4�H�X�M
���nl͐��hr���I�V�;	s<ƤnW����c�!SBJd�'���������Z��H�L�ß*2e�����$���%�a��K��b�K&���KflL*�X�X�R������C&���%���&�(N�I�%<iB���烑�@2�ǊFG��=�a��C����P��2)Vdx�L X;"\���V���L��%Cz��S��&G(Ѩ�80QQֽ%����ʙ�-�R�+��c�`�[��@�c1	���`䊉���C�}\���փI04�(�y����I�0 1yߜ��^J'����&�Ħ�i`�!�1T�W�����*�H��r��1���	@"�m�dBxU�Ķ�	XU�FL��^��*B|)�J�$x&aH��c$X��Z�Ν�;w��so�Y���I틟}�����__���0����]o�-�W|��ڻ!2���p�����bY��_�By�*SHmi�;��h�o}��..�U�ny�`s���:�v���~���w^n/�'�~��7]�}��_|zks�jq��xڸt�י�<�6,W2��v:<q��L��G/����-ͬ��:��u�-��lP����x�C��|;����o9��{{�\�Хc-
����AC��Fm���!͇,�yǶ����g��{:0g�����K���mSO
�O'�o��z�<oz����l||:|�w�����V���Ys�2n���ʠ:���G�<��|ʴ</Z���S�魽eY�c٧D�tUN�v����N�R�jr��-$cUZ��f�,-/���KD�G���ki�yu�W�z�Ӌ�;n��<�ꭇf��Jke}�?X><>v�j��雕+K��m�����`��l�Y�\�N�����g{+�G'��|P����/N���9�����W/w瞶�f�3X:ٷ�N�N�Wm�jm��\�m��%�� �m�v�'K]}����YM�뇪+�+�Arݾ���c���i;�;��������?+��Ͳm�7���S/a��^����*��Vs2�Dy�&Ve�T��]�zO�R�E�V���Ic��ĥ��`uc��z�n�h��q���՛�/�{�߹�qm��'Ϸwv��sqP������8�|�����`tc�8�]�֙����*�-�{���Ce.U]�ީʟ���4���:�[�4l��������W���[���/�:�$�4h\��.�,�Ï�g�������wl_ml��5.�í��ك����o��;X��#OnL�.l�:ݮC%i*�)����û*�,T�4 r2!z�X�BK6Fra$�j	`���<��X-�8��"� 1��_qP*�����Vs�~���HQ$���:EH=Y&��Ǐ�;�z���b�����+P��H#&��$>�Z��*�h��� ��Q�L�]F�gb˳�c�����b����^�����;��*�/{�����c�NI�	� �/<��)7W,��B<oMZ~�ͼm�j[q^g�tx5�ԕ�2��eByP�<�6�����g���xvjppv~py��/��k��K�{]]v�?��}��h�}����!�[W�=C���m���~�M�n���0>:�Y�����_m?�-�Bsܕ�a,/�/ :��O�[͕7�_�/x�M/�lپ1j�������g�?��/6�<*��N����ߞ�6�;��=�n_�����>1���fByf���ײ�i�'1j'�RS����B��K�����ò%�kp?E�F<��m�����^�}�9�_�S`�]��Nr�J�S�K6��5C2�y��+�KHՁDfB�l�0�lu�T1TI�JN��2�T�T+�QLBKɑd6R����Nm!�	�����5k�6C�����bmϗ��3Ow01=��$0r���0a8�5���~1Lz^�/>|h��*-���䅡�(SԳ��-����I��}+8$�_���V���GeS�-rk[�n�$6z<s&�=�/^���|&�Th��)GTa���_02��j��Qa�T��b�ǜ�ã�R��W������0�V���;MJ�"0G���\q�s��t��,�ų���Σ���7��fg�P0�A/1��h$`��������n��C�0�km<Zk��5��9��^��g�$Z̚��g9 CI_�%�������'���	�zɰ�Um��/~�sܐ�����&c�+�?k��� �;[z=������?#(N$�?1�G���9Њ��m���"C����M1zl4��s�a+��c�M��d$�J��4Eɖ#�B�"��淙1�a�d����I��PB�a��c�A[��(�u�h��� h�ĩ>��az�x��F�$<a� $BE9sl8%��A�*���bz�K�-Ȑ ��G)OoD��'��@��\�\��FN�	�R��42������$V�Y�"����!��j���D�Q���*� ��1Bx`�KlY��D�F�� �49V�W���Ue�6�-̙~	���+�K��Q��c��,� �N/�f:w�(	a ��_[M6sT1w ��M ȱ��W�IcR��9UbC%H�H 0NmQd(���* R�6�C x�x�Ah�M�����L�j�"`��i�7HE��J�0p���*H�� j-Y�y�	mj�0i� ��f��6�*��kZ2E�I�h���"_i ���.x4�j�]�b��9%y`�j�A�EK���^�P+�]��ЇDd�*zHU4��V�@�!K�3�P'ģ<&�� �P�.� WKpH��-�!u`$�@HEJ����ۦe��Q���X���&*�ӽ�ag��K0d�z2�_H = ~���`hx�ҊL�H2^�b�
�o����*]�yI�c�(N5����� ��zqM�r"3R�H����*=��(p��qf�?<��6+L��[[�dXS�]\��^��̛aH�"�Y� �����5�s:_	�,��_�e��iDUS��LO`�0 	Lh�Q��"	G��j�0�]g��Q�-׫4�Q�F�h]e�Cd-��D#x�&�ėZ��J��,k�1�3�RL4G-e�d ȴW���h��Ą�1b�^
8zB`A��GA����0x�:!M �4'2WIf()��Q1& qMO0%�0�/}�* �p2��O��)%��G&C� 	F6̼@$�UI�j#�
�"Y����<��6��ê��\h %X�LPd.��5!A���K�A� �T�鑢��� �v��P+)&p�t#9ʘ C�˙�)��$J���6 qf��1�F�b��N��m4��!�O0� �� 4r��Z��b		�2����V�Ƈ*z2A��x�I��!A"$Yp�'y	}��$�i]8Jz�ɪR�'�[OU�5'��eV�i�@�:Q��@n�j�h�Iᅑ�#g�ZǦ"Y΋�  �zH2�Ġ���u�!�!��( H�%����pp�
9<Y $�h(%�0��)cNFR�M�<$`d���b.�������2dm��9s��uq�����
9�r�Y��Np�9�n]�v5�G��Ӄ���/Z-��w����Y��>o��ɷ&�[[KW ��M����r�n�GC��j8�a�P����ҝ�����8�"���譭�V�������ۻ�K��������ݕ���v����,4/��^Z_L�!I����]����ٴu59]�V�܋s�<zb���_�;�f���h▸��Sm���=��+k��I��m�l����Iy�_��q�:^�s��hW&��I�Q���+wz��X&�L�uo���һy5/U]w���C��3?��ŵ��>�X���_���y�ur��Ʈ�g5��y1��_ڵ�2��ܒ���%��0��a��������誙��� Ҋ��zj�\���+�V8N��m8��d��W������ٹ���Ա<z�[W��U/�"���\Ї>G���l^�0�R��p�<��m�ݸ}me�m������U�����G�|D��������F������~8�y�1߽������s�R>��:t�����p��ћW�����3��_Dqٷ.�'�����m�*{�jElG�����HR�)���(���xxr9�rÿY6p���G�''�wol�z���v��,�{߷�irvR�S{��w�<������g)T��z��N�*�)KYiDY�ZD#�~�%@��ث�L���G��ЛNO=c�����?�gu;�WۇϞ��c��?��ƍkG�Ý��\�	�˯ ���v�v�/N�f��AU��.z	�{i�v_T[�?�F�{��
�}��Ȯ��J[���j���:�C�y�t{sՖ�Z7-E�5�<z�meɍ��o������w?��\���ܼ�y냵�k�W�]nQ�x���p�!`��^���o7,�`zag���s�>ԙu���	� �� �� G��b�w3R�~��4MU"E��F0ݥ��=���a8��"3!w���e��^e�K/���i.����P������Tw����{r~D��Em\�' ,R�Ҁ�!�x�C��2rZ/P���"�4�/���z13������+�H=?1�K�.�76&>��Z�3�xu(z�    IDAT,L�cU��H/�����K��(�4ń.��-�q�����
i�N�3�$���Ѫ��t6�\^[]\i�9[y�͟��ӯ6�m�\��N.=�i�l�3�:�s�;>��6oxr��ˠ/�0�����e�3l�����-��!
����s�LF�f������|����LKj�S~F�p���[�?���������./�3��!��h�����_~����۸]�y��X����hgr��t \������ת{3�S����Fe���;BL�I9w��Z-�V��Q���^�Q.˷s~N����y9��c�QV;~�r���w��.p��9xgz_F-��[�ˋ��2j�d��N��)�:sI�����D&��	 ����FCNс��ƬSw�9կ�Ҵ���$��0@�(6��`B��hb$�hy���  �*`j��D��hTs'�����1G�  53�rz9�UXB�h�1�
?/��&�j�*�����Z | �u7���%s^�[��Zkl��3A%&VJ0�/A
O���<l�VH�#�rzg&'xw�=z�\�Ѫ�L��S�R���ߣ"[����!��`ƙ� R��?v���<w(`�kc6G��^�w�G�q���Ύ�eЍؒ��e:C��ޛV(�ρa�b&HE�8���9k.��M(�8�&ǃ�@]c��v��Ƶ� 1�+yAŋ�h>|hdQ���EN�0rl�xс4x�F3sC)�cN�Z���'O��n��K%C)NݮE�����@�L�`���b0���䚃=m��2�\��0�]\+�%`�k2%Yl�4d$lE�H�CEӉF���Z)���� ����,6zE9�XӋ$�.�{����'i5J$R��Mc5Y��OTi�Z26r�,������� ��O+h�
��iz 7@ȿ��A�*f�1$@z���QT%��J�UG=�􄧨]��,�*.9�3M-P*�:��@�/BEU��<�%��v$Zqb�!�B�����@Xo@��รg& �TEJ�*y<�"!����4����U���*	mb�ǜZ ��CF�JєS���� �zq�#��$61`0X�9��d	 -!N���h�j�J��je�^�/E/i�c=CNY�AӢ��i��?E��|�u 8sah��J���@+�u/}�
�R�)�jsE^��%�Iz��*�	�R��U��E%�RE�a�'�@F?A���`�g�%�\��2�40��		L�,6�A��ah�cC����>��%���w��o��IH�҄G<�C�W�$=/1�2q&H� ��tT�P�i�O�Ϙ�ט�А�xL'��R�Bl�`��a��R�Qj&%�t&[u�8�%&��/	8�@��M_	��#��V���*<bc.~Q%<}H�)0��xgɊF ^������!�8�GSF��f��!|���b6x0[��U���E����0�%�Y��.��K�0IhUI.	 ���Ö3+�?�� A+l.\�j���	`�A�E.� Z�9�I gj��֬L�c]��=M p��p�=<B�U\`si��� N���<�#g���9ڨOrE-6x}����p�^�X`����H3��~ �
N����0G1AT��Z.ғ<"��ZU~�� `�9���`V�aF�PQ��TK�A�F%T���U� 0��a�^%'!ѽ�,���!,�������!K�j��xT�'�cC�����S�$ y:V�����#��`�?x�c%���.Q ��!���\-�$N��F?�Ti`8� � s�����J�\��K���CH���M؀�TX�]�`b΋b�I-+�%�Z��!Pj����PC�'%Lj)S���\m��\ؼ���zOK0&�����$cJ	C��*VUx�-�(�x$�� �H�$D�$�X$ ʸ��� $�x'�	j	��b@�I	�������wф6�yBJ3+r�0��=��xRI���,=�}� <!$�
���\-.bN&��_-<�GJ�d^��4�/z�^�ON`�zA�19��Q`B6O䵯�ʙ'���Do�E�Ʃ���ZˊhB�9�#d�9i��'a~��]� D��md�	s�b�D�H�F�����-M�wJ�v$%΄G�4!��JC��f:Z 1��p}�g�<y������ooN����;���#R�uG��W�:��n�z
E
��g�Zg���ltuQm'����έ�mW3�{��w����v����U�:��A���!j����6vi�jxAԨݼ�Zm-zY�?��޸Z^Y\]_�w����5���/�߱��:<��`���̡[�248%O��a>�v~�Uˉ����n���۶���1����׶]�%�%U���J����s-��՛����^�ٞ��[:�8bw��rW%���K�={0�\pqоq���O�.ټiv�̜�OW��������p杽��;:����\�7V����3��'c�vL �eͽ�
�ؙ��8�#�T&x���m��v�ϫv���$7��ѹ���p�k���Ո��
o.�z��kw�C=퍭�N���w'��d��9b�6����bge�/J{��j�ֽ�?�a~z2���F���?�����R�3��~wx���?����Wώ.�����?:�9u��̳�����ƖC��,�kò��M]�;w�Yymb��{Ye�/�z��vWG��~�r��<mN�V{^?k�ϕ�]����:�7���{��7:=|�����"���e��뭒�u�M���_@�2�SR!	�(�fW��O��\/V	ىq��`�_�Z蜙��Ë�/v�������óg��5ge�C&�/~������u��.���'�H����o���~���e�ӧO�.�1��薯����w�=~��7�����W�=K�f}����h�����7߸���xW�4���W䈕F�����>�|����?��7壃�#��o9��:�͛˷���o���/��F�G�j�L�C	���J���_�aZ��eE�*0��e^��b��P���4_(S�O�b���K� �L#�i�YQr��p&�*z�>�p�8�q�Y�U��ݐw�˃~:��(D���)�Mvc�1=cU��@a�@�4�!�̈y� ��$V0VCK�,��z/���
au�e�kAn����3ȭ��p��N}ik}u�0�[�s�;�=�'��򔵧�=�i�l��kk�6��zO6���U��[67�m��tv�=׽v'�?��8u�����j��Һ���D��/[Z�������[�n�O������^�1��F���d|}u��ڂ�����i�s6�{!���kN?���g��ǯߔڳ��`��������T�NO<���t������ho���Aז��C��8g��9v��~j��λ�^y��d����~��~�/��ʤ��6������O�V�r-[΃����Y���^c`�-���0��[揗Ï��?�)�ǫ��:s�~ȭ���j�jy�	�S�%�d�Ms�{q5�?�mﷶ�[�N�&���_�dޗ����\��y/�\'�'"T��粯�Y��J(�L$z���X��|c(Y�!�j�����
EIM�z�-%���6��)œ�"J`���J��豑	�K`0eiT%�Km�r��(Ӻ�JU�>�%�x��s~Y�����J�x ח�ii|��?�)%���BwL�]��!��%&��	�E��PQڸ�¨R��c�㓜���»3C�V$���#5�#�k�`�	Ӑ\��X������Gr�.<Tnߔ%�Z�܄���$���.��_o���5��)�d�!`���hp��)P����׵���� &9@N��dl ��t���;M�t�B2A┩ƅ��Z�a�}�������������7~ac�@���ڜ���J<` �PQ��xL�j���+$FD�r��'�h_���VlFPս{�������;���@�	^+0����C&~z�����̻m��(7% 
FT�Zc���0��F ��[Σ�@-��(m�`�J����F����`ѧ'É�-w�SV��/yɬ�=�ȳ�ɘi�q���ѷ�N�*�6��Z��а�5?!������ju*��� �OsX�	���%`��*.��� �B+<Vr��z tT�"�0s�f��zIl�B	<�*�f� �Ҥ	d�,Md�!d[&�i8~~�j&p�H� �I�0�N�T<U�h�`�!�R��a5|F\�Ee�@f%�OIC��3�-�ůJ�r��a�!$x悒; Hz�pb�W�&0���F�jɢ5^%V��9$1Ǡ�!B|ᄗ2x`DCC�#�	%KS��$f1�c�T%�ןR:�����*�`�F)���D��:����ܲ�x��I�� ��M��Hr�e��	��?Y�
>�h`JU��'=2��d,�+
CU�X�D�i�i!��2�t2!��?�40^pR�S�`hE��^la�痕&��	��&CU�_�{���:SP�~��z�6!ѓ���&���c�HՒӍr'M�	�-@����Z- T����x��!È�dА$&���!��p��	!��&G���̖,�#�/���)D�ֱƝ��^2�)����$% 񐝠�v�/�~Vx�˙��L�@Jb�QsxO<�8�Q����9BS=z&il���X YQB
I+r�(�!�È$��b�D!�#��%�J�jx4��V�$����Ñ�>�	�qA����E�������E	VSeV�ƣJ[�\OH�1a+V0.R=p��KL�S�� ��с�By"! 3Đ^%sģ�r�#B� �/�t;fT�l��i0 ]!O��o:J2m �@xP �����\������Ϯ��p�*�J"d���Ǹ�f`�uP3�F�F�S�Pu�y�&�)�<�
Ƌn�N�a
U��a$�`��+6����N#6q���f"��ҙ1TD%N%JݨO�NZ��km�?0i����{�iAB�i�*�Fɱ��	�RH�����&��xL_iT ��1�X<:'<��Tm*[�\h<�	 ���U�U�� h�_�\`�3G����$�TA
�8N���c�����l�5�SU،N�Sq~��`i��hu���	�~0ZfZ�A�G�ʜd�+�qaB��(��66��Ϥ��/���,�H����sz�s�."�<i,[���3��U�!�O�'$-M�F�������0a�"�b(�h`���6��\9(�:'͇Oo'lyTI	RǦ�� $�4D���$���4&b�H=�4�̑*�Q�X��_�lL�ͱ�JF0\'f2B$�R� O��W�%7ܢu����Ot�)Z��:��I�H�.ˠ� @ʹ@T��.VdU\@�P^צO�t!��
d=,�Öa�	� 3s)QM��?z�z�A�ZT��j�|���/��/}���?;�=]]�:����իŮ���J�r��^MZ����4�@k��V|xⰡ�q]��.�#�]΅}ߤ,︻��մ<�)y���P�q��]�]z�P�/F�U'ӫ˫N��t7VzK��;Ѓ^�t��~���o>���=�e��[s��v�n��X�/�K�������7�ޫ�6�ы흓�;��X讶[�vM��_���y-�3��2�^��W�A\�6D�r��g��Kn�<���	ڦ��Oot��!��qy�i�nK0�qr�I3f%��#}^M�g��.�'���\Sߴ^�y�6$�_5������������g��O=�7���ӫ����Ӌ���txn�x�^(�t�\^`��v�=�=E?T��n��OQ����β�;*�=���q���B�Q^��N�f�mi{������¸�]��O�������������F-vl8):\���1����v/'��!U�ᰧ�n��c==�k"�g��bg�cO�kq�ݵ����f�w��B�����=����oݼ�qk����J��<6k��`���^�6G>�v�}�d?���Ј2�5_˖��;���;m���9�9���~��Rf����dX�f/_~5��Ow���6>�1�����/�A�Dk�&g�󡀎N����z��`��ǟ1�����bu:���5�5�Zd�1�}r�3�'��(�Ϣ�VU������͉�6˸��O	��Yoֱ��4X�m���>i��_�~���j����O�����e�J���_,��>�x�k�Ӳ����;�N���랥���Ҕw�ܱV܀��9��U���M�����?���>o���@��8���˗������ƲGM�j(N���+�,K��T_�k����ޭ��k͵���b����;Z;q��l|8t\�>�k,}�K��F����W��PQ�ՙ���\�
��iVE]�Z�k�uKQ�,�X�͒`J��&��4���d�0���-��zC.ˣ�VRb#8���Μ�k�	f������������Mrs_R�0F�@N#�ǇS��FZm�B�$ E	��bY%zA9sE<�~&laԺ��XY��!��=��w֖;N%��ğR�Ndsj3nb��-�L�V{��X���z��tY�
����z[�鷄:3�S�s�?���Mc�HG��s��K{�S�J�m���z��?5~����~�������;ã���d�`��	���`�r�}v��,N���n_�L�{�����S�_�����޳�;���������;�^�up�;�-/v��-O�)��`s�}zzx�|w~9��ݸ��G�>|���'���o�R��r��������~��;�O�]���V/��m�.���n����(oy/���Lgyz�-�8����+�+�d�����ٝw��v2*/Ah�����o���g�孭r���g��J_�͸K��x{�BVE)/WwiM&�r��p�������Ex9�(�𔐘Tr�=������RDJ䙷 lq���Z9M�dBFKP�*y�x����0�wy</��j�<VU��� �-�Ė�E�)�\�%H��=�*��9!��X�J���i0[;Ŭ��kG�[Z �U������Q��g�<x`!�Z�̑K�.����5��,;2{`�L�R` ��rB�H%Z�L��4B�On�r��< n��W���V�m^2 H0�$gʬȘ�
�^��u��h��YT��ߺ��Cf��c�O@"0��tw�Ȼ�!� ���z�U�;_r����ú�`	,C/����^�v' ���5�؏F]'<!�wR@E#H. �f�DN7�5�xq�v�����c�&�G�iS�9BȄ�kz��CՊLE'p����&�X!�'(��
��j)�9A��<+zM��.���UC���E�$<�"ϸ@&�a�RB��'@� �a#�Ŧ�@�I<�0,$	���/�Q��r�$C���w���b��@�Lb@�J�`�j��^S�<̡��4���
	w�� �r��x����#��P`r�u+�C���*E�i/�-�<HUf�\��AN���#z-b�$�x���x$�4�&�4D���;e:�RR�g�F%��2��Fl�LR�=sI�*18�7/`F�Vf��)"�ڸFEƩhR�[�Y���:�49<���u0�[<&��Ix$���ZE��]�RJ��P�k�u��U�O<��!�2��K����S�"+B�Sː̐ �2�$2��2�3����K\��%* I-=���Z�*&HW�i�Q�QL�F�w�8�cb�U�U4� r�A��}w��+g1�l�EH�"	@��h1�FH�D�9��H���g�b�.2.*%�����Ċ>0V9����9�ٖ	0%�H���_.�I��R��Vz	'���8��M? ��DτF�IO#��a\� LN/���F�3���R��(�O������J$`j�J���?+Jy��"E�&\��@v�@
#�z��b6�{��� �K.9/LڈR�,�"��Y�"G�ѐ�!�\� ��1!���&��Pj�0*z�]��*�*#�0f��y/A�X`UxI��k&�!TD�&��qJ~	�N��Z� w4Z��Վ���5X�li�3�#���=��^�|�� ���O���T�������P-r��� �]��'H߳�    IDAT1�+��L�#�&��J�ǘ� !AlQ�\
%��;T: �?����Ix�^s�m� H<���AK�u���H�	��u��
�R� O�I�!WD+�aK��e?[�$!��݋��c��>5�/A�1t�G�L��3�g��D�S0I<������^O�Rp�c �+��f��it�U 0��L 	 �q �?H��3���!�c�;��%���3�`��b��3*y��U:_���KD�J�Bc�0�VǌX��#׊bF��d�8zJ=��>�'<9B����OhX��+fN���K~��Π��G?��ߌ�U@�����_��c�����tox rac���DH@ /��.~���QVU0"�K��+1�g�#�4���ϻ�A��爣�@�U�Rr�
�`�����b<H��X�2t&U�ɼnE"�@?��@V�$<&�p�_x9)�˝���cR��k{~�c��xXIN��}e�0LC�����D��6�Py.G�Y���×�V�}��b�)�mFqA�	��B�J�\R+��d/יfag���"�E���D�������⇁��" G� H`�� �ɨx4�ԦJ�nOx"ģR��2��� h`��I��n������wqJJVH� �s���n&����'�8�L���f<�du�]�M>yx�=E/`�*����;�|Art�9;�U4.��h�-7�6�{�e��a�ݳ+��k��7g�.�b}{�qǵ���&�� ����:���֦�5=b�c�v�+K��.!Oz�6ڽ�cՓ!A�L�M.�|�[�{B��-S봃�~��]lY�����,ї���{�m�^���x��v�a�ONFeGS;��%���=��ywce�)�r������o/itl��(J�������2�e��3�nwK�3�W��ϸ3x]�;�������:�q�̯�N����o�������[;�G��:�ܼ���/�|���ͥ�S�L�ڋݺ���.��φ������1,vu���YK�i�������|d7��7�7�]y��:9��8[}�1Ӡ1-�)�Ss�L5��s>�f�׾��r�]n���u���t]N��G6{m;��0��s�]���QY��z�ˉ�4]�nz��t۽�T���ٰ��_�/�W7�g���zg�7��׍^�$j�ӿ��i��`]��A��l^�B0�1���N�f�������r��&��x�YںZ�����&�ڗe�Z^{r2�@�Ҋu�����W��ӵ�ն�<�4��9�����O�ǥ��-U7o�Z��0�m�M�k�zرyrqlWO����#G��҄q0̐2I���U���Q/f)Ue�UK�T�����F���r�����_>����z�љ���󝯿���Ĺ�ѽv�3<��W���ڹ�f�Ԓ��Ջji�nmm����O���㷿��G&�#�:�U+��0'�}���7�}+�?�Щ�ҩ����������jο���߾}s�����'�ՙ�ð��ҦM�%���q��@V�7{��ž#�����Ŀ���Ǒ�w�L�����n)S��:]���b��eJ?�'�T�0��I��Xe� )��́�\��_9�	��CE^�0'T@�pRF_����	�s��I�099���=L�Z�Px5Z��	��f�Z2A� @{ʢPŚ���;2s�drVr���:VCF�����(��9�k����W�:m<���f�rp��ly��B��ƪKt4c�N������R���馑3�ws��6mk��Z����g�����<+�2:n.&�����_���?Xq�Uv=����q�A���ʣ���^y���5<�M���:�_�ڶU��˕S����G�[m;��Ω9�<�
�3'm�m-�ʧ�ov}��_�x���1z4[k7ܵ�?O�����nݽ������7�Uoȉ����Asr<;ٝ��WE�G��fn\������>�٪��ֶj,����4�����>�.kǥ�+O�Z��{��ouX���y���Rr~q4<s渘�ڿ�n���e�1_].�CFr�,�$�F	@���E�#s��1I�^
&r5��P,c��H�/���C�:HJ��c�)���m���r|�'�<���
'�*H2������J�R)k=M��cG	CEx0y-�Jm�>r�l!NӬ�:B �k�������bH2^�u��S�,�´C���x!Q�_�HI�s��9?��FN	~�����i}��L�0���6�^N�'�Z�xl��o����g�J����m�@�~$�[�l�񛖺��E?��8�!�����c�tb�ǟ�{�Y4� ����S~% ������OS��_�5�����ЏU+*N�49����KG�?1�$������CePo� ��Nd�g����/�z�)����I0��J-�����-��PhU}��w�k�ha 23�gƆ[=������ʵ%�O�<!h��" ��o#tM`�W ��]HQ��L0[IQ�A��D��c��F0:\@J	5M P*�a��F�(�K�.��㑹�c�!����\U��h�e+�L��2`�`䚍G|e8��ϟ'f�4bV���b���ax��F#N�X1�>�d��xҟj�a`H�bK�V�^zU�b�w���>�P2O��s��3}�c��\wiMe�M��?/���i$���)`	Rw	C��C�P�b�H @̯���*�D��<�4�u[�*�MmH\���V���^N	&l��'��	 lE29��+a�+�8���@�cŋՆ\��J�yX�	 RB�NH0d��;��$�ht�N@�����dHU	8�U��Z��4���6V�娡I0uU"dI���E.�5!L��3�2@�^��G/�PQZ<#�#9=N�F�rl��8u���V���	��y�G�`���gp)�A�$IU��B�;*��lrJm�! G�)B�H��3�`�d�R"�6����	����;6z.�4��.`�P���4�L�?�|�;NJ906E2�@0�UHB~���rdΉ��-+T��Tg. HIW�f��H�Ow %�4!s�k���q�i��z����t/8���$2�N�4�E[9�32�E�[R.x�a�5dS{��*�:��U+W��"d���8i�C��dЛ<rlR˜-ZU�Ĝ��2L�	��S��<�	C^�t�"s.�EQ �Ԓ��v������;0���/<��J���\k� b˼�Y�v:��/H)핳�j�3�$/Vj�O�҄�����MĬȻ�<��r|Q�`����U&-$A�d��q�,���9�0�B�oj�x`�L��BRk2��9�T�7��P�U�]�w}K@��a��E�/�I-<���	"���8��OB�G�ǐG���.<���5��L/a����D��8�4r�«��L(�BI0��I�%�L�:f$qA/)��K̊[bV�9��J�2��PQ i��3�6LH0�����	�Ł;r�)Tb����#�D���������l�r��܃�"?�ęHhLH����3�SE�<Bz��xT�X@���Lϗb�@��;����t=���_?N)3QQ�%�GՒ���|�*��+���0x�
@35JTA°���
 ��d6R
���G���Ф	Lpb�L�\RD(�"fa@��@���p^c�4��&� �K-C~���fU��8����?e�J�լc�8�*1�� jU�õx��@a ˍ�V���5A��(� �iҜ ��Ԛ�r�)�k�V��1` ��U�4�r^X�e"l!�?0���:_��������` �G���K�J<�Y͊w����)�I�GmS���NH�9F�	�ﶉ �={&0�4��4�4��$ST05xT"�T�uj���	C� �X�5��_�����^�t8޼y��!�NG�5&���m��M��۴1u!m�~vv4y�l�~}�����X���bv�OxNm%��\Z�=���A��5�W�G��[�\�<Zm�s2ގ���������xrk�5]X�uW69���)�qek�?2��}��qgvrqr<ܷ�w������9�\l�G�wp=�8�����������?~y�߿���k�o��?y��`x�p�Y1�v��1�*;���.�ͩ��v��o\O��Xd�\�=u���u�!�����us�\�_M���\?���m��_y���y��|浅�o��/�����������_<{j'��G�[g�'�W;����N%�����p����:�\��������;[�E����jwks�ɽ7� )��֥���!oɿ���]y���̤�o}�]v�ϱY$T�B��,w���Rw{�+���6#l�9��/'��-��|y೜v,��;o.N֧K�gË�х�}�a27&Ss���`se���=~���Ll����;����+��X�,�[W�j��k�6;{��C��s3m��ƍ�c��x��WH��lإ���<zD06�=�����]|�J�2�^|y~x��A��k����o/.,vϲj��������=�;�w.��eu�u�>�y�����������=�h�S+��F���BC�bE)��CY�����U&UR�ej�����ş
\^�u�ž�a���wy�sr�g�}c}���5y���B�����kk��h�՞{�k�K69�(�2��\_���u������ׯ����on޺��������ʺ�{VBwq�J�Vl[-�����y�u���P'�d��溿�p��Bg_s�����m_�LN|ɦ=_,/nl->|x�5�6W}nj�_6�Ӈ~���y������W���Z<��`z�R"KT�J?V�O�ϙ�����@�H �XQ*f�4�>���.�(��Ba�.H4�!i�HV�h*%�ȱub`�ɚ�爵<yb�3"�5�k��?�8,H5�������	��&Qjd� ���@��M(j�ᗓ��X	.y�X�)9��L��Ϧ^�|r���i��h\�٭�WU7e�AͲt�Ӂ�e��S�N��.d�#kwI8�e1�8�]��s��-Q�=n^>i�Ӫy���{�����5h���g�W;�[���4�K���;?_�����?,�\���`�u<�6pO�w�ֶ�� h5.�E��x�w��r}��{���Iǃ9坷N�QG�;<�	މğ䬬����?������{���V�	��g��Y&��X�Z�G������p�ƙ7p��&��W���c�טZ��)@y�l1�r����a��{�؎f��W�Ƹ�D�!��Ύ�'>}z4�::�����;'���-������j���q��d��cj����"�l�����V�T��SH1�+�dɄ6�kC���	�b����9r��HO/���r�"@HX��$H5�Z�2�!d��f`I1~��-&�IH�XdVj�Ҩ
-%<Y�����
&QQr��A|Q*�4E�IE��*�% NE��h�#5r��/I���dx�W������oK��$`'gJ/MuY���SA�/���s�����˹|>�g�� �B`i���7�|�g�{��޽��o��$B!�Rc��ѫ�J�b�	rmdKҷ�~뤅-J�NZ�^��zaՋ�oҝ�D�D3��*R�`��U$��E�i4�?���8jiF'?��N�Uvy���@�|���Y���ƅ����:�;��[=��P����Q��,Ha#$/"����ϟ�
L<��6�4��@�wH# ��|�!��E���=���	*� ax�L��DEfH�ը��{�^m1�T���c�ȪRm`4�@O P%��/=s)�J�2��ګ�#��éH��K�V�[x�1�4^9�`0����$0$���Ƃ �z��F\����%�F^ZU-zx-xbHNg&N&��I|��C�DQ.A��D)f�%s[��ݨ�iE�6�@)��� o��	�9��&E2!0<�� �X���Uf�Z���j�Q�_�x2@� �)� �T+EV� �u���+����%�x!�EVÄ�Ƹd^��+��&<�Zz���#�D��'��$$*���9�F��,�m4�H��o ؒӓQ�E*�j�ZqRJ	�/��ʥ 8�I�U�M`�b�T�)G��o#Cr�H�6�D���W	/�d&�w�=-�����EFCk<=�8���]�_	R^����fc�*b&hi˩��.U�	4LR�GHf�VX�EE�9�k�R�$�t������s���D�r���5:9M�0���dV|9�aVw�ly�����N`+T_�R�ZT�`�Vp��9%��6�s�Jb��F�_Ώ�0��2�H�Qd�Ps%&`��aE\��G�0t�>1���mBE�
F�����[�"y?��Y¦�4`�2$3I00£$p�0j�����C»Z0	^�����i2CUL�H����T�:'�r1�C#���
��\�aVD%�:$�D����#�]�� G�!QEH ����GN� T!cK`Kf˩\W3	�*c�0�؆�U�K�i��>NYQ�̄p2�9!�I���)�ыP�/����2�<��s�gpc�1�rl4�.�Dȯ"/�#�U������0V�)�+&*9�hj]Bs�PT�d)+�'�$2N��-2	�2I�N�"U:��h�y����LC�(3p&1D���Dϋ��Ɗ� ��r�L�L'R�	[�@#r?(a�(Qh}�
�ƔC%�LN0)�<"�O� C�EBN���6�a��?\�ٓd�u&����̈ܳ��������m4��f$�dӓd��P/|d2��H �"Ah��՞U���{d�~~��29�^Ǐ�;�����������@į��T�����,��Q+��ɩ��2���E�6%~�	��Ɵi���� �B*l+f�f���ZH�oߦW��^��F��1��S��#���� �_C�0�gN�*^�`���&~���R��oMB<��&�"�}Tq�\��l�D�Yج���#Tx�Qs�V4�>�� ���%�̶����)l0�喱&0ی��^[<a'��֡���4����?<�	#�x.���?��L���!�`0�8ҕ]�RT�Y�4���4�%d8j�4�"$�|�R�6���/�0d�3��|`%<� � q�)Ŗ�
���TgN)M��!��Q	�IO�:L8R��JW&��A%B���p�m�!��l��N�Rg�~f�҄��<�����.E�|e[�)������c��i���m�b7=����������WW6�\��`���^�����ȳ|7���yn�6=Vh�r68|���G7���3�֮Ƴ��g��Z�u}w[�䬬�Wh�AW�e_�3���@w�)��ܭ-�]ӲH��|ur�qz�W3��{7?�����+�A{���I�.�Wvv?���vn^��we��7���ܽv���>n������Zwm>�ߵֽ��������Qo����[����w�|��>��Ο�:������!vgw{�|}�,����s_K�n��㞰���icU(]�Zŵ�(In�S��5�=o���J������oY������'������V����zk������'\���F��Y4W�?{j���v����?����`4^۾�Y�7^�;�ELQ^z��υ���m��e'�{�MQ��k���^��ڰ��e�8y�������E.�\_lc�+z���s�)�Ery*r���U+�֢����-a�{5�?wg^�h�v|�B|x�_�{�������GϽ ��������˳��������׏>���o�29N�G��+V�Ǿ�3wS���ٓӃ+w���/~z�ʶ�O=�d7�	��r��p>)�͙��ʶ���q\�(+�m�|j�<(7�	4�p��|s���b������w�����_�g�H�&^��Y�,Vʇ�F��.�N���g�3���m޸��a����'�G/�L�vy�A��}���?,x��WȡX]�X�f�=�~j�دișT�#�ʶ�fT��}}L�EY�s�����,M}�v��s����V��|�u��1{���./o:�����Zk��i�sseѺ�]6�2����s��{�}��'�櫯}"�������O���?t$�    IDATt�W N%nP?x���#V=��o���~Q��p�qN�ۻy�歳���=v�y����Iyr�w4ml_*]��m���mt��7���oDֻ�c��Hh~��\B4�|BpP�39IZ�u���#�CE��d�6Ҕ�2%��+i�y����ت��R.�l8�%�?�Ҭ5qJ l��	 zx%��J �%0���	B��4EXkL%$�ˉ�ل�)g{y����kP�Ԉj�Pؖ�6HL��ㄞ��T����lN�ʔ8Q��ղ窆�|	i���ܛ$�o˞�X�\��嫘Km���1K%��l�΃�~"S"q`.?>1c�5_9���i8�8��/���j��
+�_j�{(ۏK<Q�m�;*ث�����rw}s{�<Z^"��Fs}f�ւ��}s1�y�]��?�0����}���|��	�S�M_�4q0y[دW�<	nXb�[O��n�;�Wo5w�����zqT>b�e�l[�oM������|�*djJʪ�yc�cVy²:���
�g�ɲZ{��/��9�Ŏ�����&�g�=�^��6Y^j{c��6���b��6�;�]6���8�����v���Ɇ�ޒIih%��� lkz3�l2�	�ޥ��JI0V�dT�Q���e�J/%<!$�Xx\>D��>z�a� I�a�'��❠Ȭ�&�&=$!u���aF��\L�?�`�Sp�*]0���2y FK�W!�����GvJ�k�cp8R6�c�.l�Ի���B� �a�r�Gy������+Z8�i�8�g�l������̅�k_�N��@Hs�չ?��1&8���K �v��b�0F��o����D�\��Ȗ�c%�`�R�ѓlH�S��hV2FC������"1p-�5R�L���ld�
U�؄j�r� H���Fa�{�e�eHޣt�Ll�a����
�ԶE�a�R�� =@¿�-u��M��$`���-�d��(tق�N"�� РEb���$�2����ү�8s"Z鵭��	�<�����V�
��G��hl���s�����#���E��2��!�� ��E/Bc����P�E�R� ��JVb!�L`�rQ��Uѥ	��1lh"��e�1.�́�CJ-*���L${Y��o�L����'e�!/<bSk�"S`'�.�bHsuĐL	`R��f40��K��p�� 9sl��!���=�y�r���J���e�uJ�d'c�z	jN�1ɜ!+��^/��=A�(d`���p��`�&~��Si6A��)�� �9"'��I|�&d�'�ɪD�:�~2p�"�h*LMK�Q�A$�Ys��9�� aN�!�B�Q�s
�W���Ra*�1&	M� ���y���vdˋ}G�B���k&E	�;]��[��~yA���	�MH
�^/f/+�J��e~zM��ATɼq��#��ք'@�$*�� ɪf� 儠$l�h	j����A޾�;���6�!�.���1�(��%<4��
�ХV���|�<J��� ����|e,�H��%'�ؒ����"xJ` �bS�92><�a������'�H��ư�;3��Ä9$�1[��(U}��C���;p�ʥN��H$'�:4\�+hȚb�#�t		mF��R�l�Y��0	�I <s<�dH1 (b��`�1���"��Dm���`Ph���� 1L��]�|g"��	C 0!�Ȅ-��'62A�kh �\[#2��l+��f��7�`h�]%r!if�`b��4d.��b�˯.�`t�d�>��1���5eC��L�&s��G�P3N5��ъ
� ��ʸ�a8u1$��\ob�'��Sz N�}�>���B1�4�d�@�p�G�9���(5�M��&��H^2�F�
F�w��ǵ�Ī�C��.X�%#a���Y��L�N��T�"`K��ĀF`
!;��{$��Q-6	�
?M�x�A����X���$�ɿQh2y IH�B$�T����yD�\W�l�bh^����Xr�$���R2.]�^��^.�#�B2�C�Kd������Gq����)\&��!�g���J�y%�4��A1�$ֆ�#~3A�7�?$'�w.��K�)Hz|i&3�VS QJflQ1��@�A0d]�̐ѢX�� �C��W��5)�����6I�7�x��=��$IB����"����0ӛ��l5�adZ�B/���!����%L�m�l��+c	~H���[��SQ�9�Lc�G=��U�=��2?#�{��+�4q�W���H�����X#U���1f+SF��49¦���-�^��G-f!q���߆R�ń2& �j2�a }ƥIV`�+��b���d�	f\���@���?s9! `63�<�Ɩ^)ۢ�N�>�O~�����7�o+�����lv�����b����{��6-��o�]:.L�s1�Y�ON�[��������0��{#ism����7��Γ$^2�v��@���Zea�z��W���Y&|�
��@�h˪���Y	�����=����{W����o��oZz~�M����gg�?<�*�������}��+e��1v{|s�,���׻x1�/���3�u>/<T�H��%�w���Yc��s���ƭk�U���-��,��{WW��������n��������5����jX�����K�!SMɵ��d�s\�ά��e��=>�{��� ����+�㳓�ӣ��{7�������ן6���Ε�nL��g�?��t|dѸg��[c��g�[k��ɨ|�b����?}�J�a��#p�7��e�;�Y�b1���.����v�k볅״v�o�mn�қEa���a��D�	��b�kM{����K�3Y��i�5*��\w���X��g��۶�i	pk����߽y㪧tMߓ�7���ͩe�٤18/g
�h-�o����U�w��������wt��??�������^��o����r�w������'u�}f�C�����ds̑��ͫ�/�s��,���K�K�ٗQ���f�͡˕b��[#/Go��>[jZ������ׯ<��Z]�r���5��5j�\ޥ�]]��[���^�9=:=x4�>�����;������?�����?�Ë������/������z9V��g57��g�V�f��K5�DX�]-�$+H�S;PD�h	�sz�!/��&�y{�s�m V�׶/dɪ��g��^a��������׵��|���l|1�x�������~��~���'/���կ~�Z���K���s���^�cLD�`b,Ϟ=s�����?"<{���_�r<�|��w_|�[�^���X��p�;k��[����杵�7��6�;�[��m/q��:��G���i��"L���+y�$�&��t%9��` NJ%MS�ube/Ȑ�K�K�(I2!&����A�
B ���Fo�jғ��ã��i��D�3lN��Q��ϙ3[&9�i�
G�8�IX�Tn�נ�� ����&����iB�3C��L��8�a�!P�����Aeh~Kb���^]����k~4��%կ&�K��*�N����e��)g2;yy��v�N3�2�Jq���dy����<�����/����Ʃc�e���t�1���r���ږ��6�o�"�^��;U5v�/vf��K����:i4�f�~�wC��N}�xblzk�@�]�B�Xesպ�}�{Sw���Q=�Y������d6G�х�F������Þ3�5�2����������&��\�-.5JO`��5q���d;�N�K���IY�u
f�}��
�U��8G>:�.�ǧ��^���o�||4j.ݺ{˫|-W/C([�D^MwQe�k
(3��Fn.���ԧ�2桪"y+]�� �!��"늡�x�KPj��hn������;J��9�$@�<Ɲ���+�04�%i߱OQʉ^EW����ץ`V��* ��.&�`Skj~<4��Y�K@�r� [6�^�&%G��sHI��8Q1ѥi�s�	C���|~T��F��!G����q��w�}'���G}$i��Թf�K�NE���;J�s�f�3��]�*2ϩ&�;�9�-r�p1m��/F`漠��_�Ld	B�����<��Ǌ  �e���������(u6����oݺ�	�/�<z�H6�NV�eXHy�.���p�����x��>����"[�p�59��S^l&������:�)��f���RD��_��$6��%���_����/<�?K�H]:0A���pfQx$��\�O���P��ZMycBI�(�DB/*`��v0 !!���7�� ���'�덆2��M��@X�-�u2��ҌSM%^�2��pȐ��œSv4̥Z�$P0�l�ll8�v�[;+zT�?9�DP�Ķ�2��P-�`�	زu�Y�"]x�A���x����L�0j�u��d�!p��U
����Z<���L$�d �	�	��P�mM ��JN`n����@�U o��	2Y�e~b�Fϝ�A�T��� ak뭙æ�Fa���:�&*
>r�x�F\��f /L�5k�4�a2��zQ��/�B	���f����0f��J��Pj���SH����&d8a�I�(�j�tq���Z]�zi8"S2q�ו��4$<f`&`8Y�#%�-�Jq[~3�HQ���c�F�ɶ&�a�ș�D�[k���X<`P���	��zal �u�!cK�5!+i�(dR�j�K��0���&J������$g�=0�!�@��R���gҢ7�Jo`d�Hb@P��b���p�0��!0L`d�&�0�gOVI/� l!�a
��R 0L�ES� ��g��6a�̋�	0�Ð	w��d����5�X��i��$M�7Th!��B�$��E�����`P�I/9�IK�xJ��G��`�d�l��0�	\ !���	���QP�KO��f�2���ӧ1ԛ���<��`1�
g�z����
�f��tնz�ir�� ܱ%׻����� ����I�@<��4�A�ǐ�ƓsJ$�.`5����ĩ	�I6
1�!#��Z�N�
5��0��Α9�I�U.���)G<�d,d�x��(��O�\�҄P/p� �����U0�FJ�/!}8��0�+0F�A�dF�\`jVHĩ���{�Cf�83@�
�:�'C'}��0H�"fM�l�)#��+扇RS03�|��bR93r��<�1�) 4
wdz1`CNIÄ��a�!�6�� �PS4����(��F�����8+�C�P��_c�D�0�����`ԹP�xX)���F�_3K�� ੸�?~��
#�I�Ö���"I���$��E����� G�
T	F�a��7#A/= %��L�s1(�8��h��YqGɐ +J����K��ސ�ǣ.��Z$��X3y��Ʉ��i����PG!-|v:���yRdthj|ѳeUQ���,�䇒��.$]�`2F�� �!��R�����"HKF����3R]�VçD�]��q1LC�{b³Qr����_����H���L�\0'0�"+�)L4�/5*��I+^�g�U��_oo҅\�B
	��Oa�E`4���+��L6���d�����ݻg���� :�����s)�ե�Fgk�Jm���yCke�����'O_~��k_P��'�������l25�=����-ӥ�k�ڍ�v��L�׈Ά]�X�6���Z3ģp�x\�%9���l�L���f���g+�����z<����=:n���v��ɫ���g'�;[�~�g;w��t,�LZ+.�/�-������Og{{t2�C��M���b����^�q�"s|r�:|����EY#���p0>}��փ֭�붶Q6�*y�=��x��?e�/l�DH��R��Q�æ)�����_�jM=#x�������h����㓵kΪ�3�eoNZ���� ����Ǐ��h�|ǋrX�2C�z�����|������އ>�t�}4.ӵ���S�ޣXַ|[��
�=��/g�͠l���K=}ذ��-�7����V>L�l�/W}e����7��f�r�o�MF�pP��ll��ڝ{<�����n]�>�tH��~�����Rge6X���_������|e�_��1�\����7?���O����}���w����������[����-{A��FY������Չ(�B.�{J�餻U���%���.�\,[�*lY���V�|KҶ��-��h�^�l����BJǓ~��ܾ�����d׶J������\��w���ͽ��[�{ׯ�<~�p|ԳP�]�n܍�_��w����C9����!I������o	,��mA��e#� �4e�Wz�HY�{a��?��j��\���1��}ɶ3�9��S�����k[��7�Q��ӱs��7wǓ�o޻�����/,�?���������'���Ï�u}xv�{w{6��'��>���J�z����b<{�$0w�sPq����/,��-��%��ٿ��O����'�|�t�k�f�*�sss�W�׷���ؘ{�͖�E�^�>:�(_��������J0j��di���m��HS�:��	0��tE�$c�Vg��\�&�g���p£`[٨1�z!���F����H~��dBV6����3~�`a�9�����Y�\���'!&e���2B_<��^���.I^��dB=HMԱ�I���X�&�Y@�	����T�V9,cvm��qČu����^��#����N��#���zyvy�-��ǣ�I�o��y��Iy�]��,?�(��_3x�~��dS]���@�[�����t~<�uOg:s-:~Ҝ/M�|ë�ΛK+�Ս�5+��Vytݹx��Mk���F�zy�@��r*Y��jF�Tx��� ;Õ�j������hU�.z�i��ß?�����]�2�Ї���~�9����|\Xj�_ؓ����r�,s:y��N��o�2�Ĩv1�MQmٗl�Si9�M>^;'�糣�������7m\���R�P�-T�!�� ɜ������,1W� Y��*ǁ�ieU�����T���!DH����\[���do�ɄD��F����I� 0=$fM��D��I�V�l�F/v�ĠIHod����i
2p��2a��f��)z	�6�&[r�a&���>�B���#M���	�F��(������/Ϟ=�`��E�o�\�&~�3.�0L\;���A�ű�	��ː��ܣ�3�؜���s�0�mb'��R�� ��j���<ـ�������e�ݻwu�(0+��w���c�J�?��=���`#B�o��=B�?�'NWo�:Mw/�5F	��(`�����7��bk}��D{���<�ʣ�I��U^T2)N�pD��-�"`0�}�v=�D�h���&��PNL�|�D���f�%E�F�G��K5��C�� ��A�T�F\��mƎ9�!+�F)�z!�.*��|�L i�B�ԚH�3.$�H4ɐ��Z����F#2frJ��0&پ���C�LH�(����^%�gP��3�����/��� �5|M������S�9c!p��.MH�$'0��@e�$�G-�'M!!$�<���[Jr\�LBh"��#�V����B¦��:�I	b�& ��FEY����(��E��	*.��&�5smȄ̼;~�sJ<	���	O�	@�.��Ї�f���V� C���
��="Q�[�^I6 ��%JH�lS�r"7� �)M6���k�� $�҄���!ٶVh�9SN0$�	�^�.H�MJM dV�Ü�dhh�4:D�!�0O� 	@}vI�����9��d��F<�%��IȔjA���M�`JT4�`0$��i4�D�'����3�1(V��`���3FB��[=M�j��YHx�����/�$��K8�#��m�H �:�dѪ��^��j�H�_��]�B�X�4���4�m�j$ ���bh�ز�ă!��X��0�h}��O$�1�r�
>E�/`B�H�%O�I]�V�$�pft�eJ�	��,���]�2���̵ d�Ro��j,�a	X8Y�Y���8������5}H4"4^�t�Nf��0��U    IDAT�]�"O?�z�y=j�
�bI͖.�$J��� é&��FYEZ6�I&+�L��bH�&��mt��	��^�$����,��%�۹H�y8�
��
9�a��ĉ'�3FzH���E�'��T���X�r��و(i�Cd�6�>B��~ES�m��t�� Jz�(5��9��!�ǐL�U�z��2��b��ì��d&��D�M@6��g;�P�)��c�Y��S0IVk�<�Q�X͔Pq�U�i$�l�.���d�8&K5<!Mc�@H���r�O�/�\��Ao�a��3�!EI�^��0��כ&�.$0�ޔ.�@ѫ����'��F�pP�V{[Hz&9����Q�Ā���DHC�7(�&AOb�O�h*oo�^%`T�D�QP�'&��#$Df�C��ш�q��
=�D[ؗ�d�>1�yx0�/|�K�! z&1ˀy�$á	m02��� 4mN5	b�$�jz�J�5C ~�����e�*��`E//a�}�@&�)B��zx`&xt�)�� �K�׈�JlƘ�e���g�'�|��T P)�X��2��#3Gk[ 3�&�1S~�q�V�� �.r�օ�6�  �&��'�1ԕceh8՚Ǝ�	��=�4CE��:b�KT���Q@&�<8z� r5*��������h���n&������'O������k�/=���r��$Cco�=�~u�����o>����Eky�̦w��ݸ�������ݟw��w���+�q��g_��Y��c�\��~�������ڊE%S�z<���%�q�]��"���I������tt��w�1���{ok{���p�������������Ӄ㋻�G'�go����o6G펁�G�����>_Y�Ng�f������̺O�y��Ĺ�y��������dҜuV��t��d�lvt����Ȥ�[��I��1�fzXS��V&ӑŚ��ʲ6���m�Zv���¼�"�ZYQ�-�6��mq�����=;>�n0��W[�����)�#o�y������ǧ���K��_\�$��6Ƨ�'Wn_���rg�*�t���X[^[�4׬ؚXV�,�ڝ�>~���?m�,]���j[�\�v�mb�]u�k8jn'�K��5�Z.Oκ�?���|��mQ�"�$��E˓��I��DY�<5�����w��Z��^��X�t��.4�ܢg�ve�?}��@�3ߥ[jn�n�olm,oZB]����s���/����'�n�`�Y��i�Xv.��/������Rr�ڮ8�̺�Vz9xsxj�y6{1��}�,@].oX^i�������-I�80􇋙��6<��i��N9& \��f1O߼靝o�6v��xs��]_�\���|�zt����ʭ�WW��Z;����M;�����j�˾ɝb�+v��\�[��R"�������)$�B9ǥ��(޹��F^޸�XYB����7V]<9m������W�^z����o��˓Ͻu���k~�w�s����U�.$^[l:?-/�pC��������9W�-���<z����q�i�����*��;�>x��Z����������߿<xs���^_ݾ���-�Xp�^�V�~�0s�tD��:m1��Q��vmӠ��y��o[��$SN��z��J�^M�58yӔU&�@�8O��3T4�aN/�J`j��|9hc����fs53s�H��l��`�����g|2H�H�NM���i�l�GUNii�����Ah�����DFB|k*�e���(2�(�>�ćAr�J`�1w��SR�2R�Y�L�~*s����o~�7������֊;�����jzۋ���c�m^���my���N7R�VO(Z-1AȌؼ��t{��0I>�i�x�z�U��X�lO>&YVW/���%��ö^����9�����#��1Ѳ���/����-��Z���gҘ�ڰe�y���t��2��t�kN���Ϝb|Fsx�I?�����g�}[���V�B�^ ��hF&�����'�������#��(��2fK�Y��~j��qYE�$��������������'���g�ݫ;~}09��X���'�m2���9$��k2A���� �4at�	j`MŔ�@o�`��ʾ]��a��u�Y]h�ɔ�Q�-�B�K!�┌���^Sw	�&�4�r1qD��	�3�=�P�(�
����j<�P��.�#%0Br��Ҥ�Ԭ#q��s�̕=_�����E��K�,�B��y� �Kᅌ�:�͛7]�:�X�t��`6�?���?N��Ǌ#�lb��_^0�<u	Ki��[򠶖F� �e�6�$?{�l�Z-�NN�\��O>3HfE/CQ9�q��X���EU����L��;��گ����d�����R2��6<�qqD#��. Y��_�����׾��ӧ�2�@� ��^��ϯ�w���
�& �M��� ���l&V�U��0�b�x�
�2=,j�-C�ȓ:Cs��J�J6%e���l�71�߿�ߛ��ӫ����p*�M-����+4L(���E��
sҨ�1C�_x��$��5	ZI�n�P�	�=%<d0d�UM�#�B�+��K�ijlǑZ�a�vY9.�
� e��1XI�(����Y��:sXZ��JF��p�9@�-d�J����"��m�dz�es`�
)N1g�!�f�mzQ)����B�$�P%���	 ��WhԚA9���(=���I4�����jCNSҋ��B�J�.��^%H�:�:� ����(3�!kw� 5mN�1�4��4��-����=�b`BN͐ @|hhlÌ� �2�dBo�dB��Vc$�fx�B��d�"x�9 'z�_�����7< x$�		��m�	I-s0�� F�jN��C� <�؛��3�T+��AIr��{�	�F/<0���@/ 5��O"L�a��p�h3j����ʛ[%�	�>Br˖&��@��Ã�iE���6� rX��#�	�̖^��x�(������&����^�FIl�p�	CW8ix	��5N��|�fe,�AN��m\ ��6M�3R���4�A�ͭIV#a%r��E�<���H����8i`b�YTJ�b��O���#a�MOC/&�d���%�
�&9M0`	���@�L�L���x�d������`B�m`j��R�.&x�$���*��Zo01�:؂LM��v��-�ޘ$M%[S��e4�0�<0u�	�"*]���'S�^h���l)��`�b%c�jD��2`� ���	۶@EH���3��P�ap����P��H=LbCŶ���Q�"5[S�	�dI�uAf�4�#]`2��@9�z����a��, �^�� (#�$\Sod �`���A&W��	�̋���ˡLW8�Q�r��џQ� ��AP�*�謸FK�
�wxT�{A�!�K��,��h�!g8����� ���N�SluE��ލ\oJRTg X`]j����fE+]�ƒQ�c�Vl�Ƥ���)�`HԲa�ȠIf5@�d"6MF'B��i�IƜQ��9�(l#3$@�"Ӈ��L�\��Hj�%6�3#�h���eB���x0C�� �<&��9�3�	FNl��C0z����R���-%+M]4�G0!ׅ�LP�9��)iI2ASa�+ 5�w�z_�x�2���_		GdCc%%�hidUo�.�XQ*z��2QPrA�6�$Sz�&1�3@���ƒ"���GK�0ٔl�vf�4�0�+ȹ ئ
��2"ץ��9�d�f��i	 C�H�X��x�5���ȶ��Dbਔ�S��D����\u����U+oh���T��$T\��cOv��!Y���OE���ľM_��ѐ����rwlY�3-��ɛ�/~�ǯ���l�w6>_߼��i}�������뷯~����w��<|�;��}����������O,u}��33k���=�趭�2�m;_�e�[gf}g�b��V��Iyu��tp���o��7W6-.���x�����'�\m�L���W��W�:-_4�~��칻˓�����W�����y�����ų�[���7�|�m0�9;zu��|��acyV��e���l�O��d�D�ә�VY�t^+�#3O���d�t}�A��Y�uYA�A˽��&�>�g�'��:�L[+���F��փ��x4����x48:s�Nguu�.'�_�zy~zn�Z�a%7�"uZ�c�
v.��^;=����%�Œ�f�/O	U_��9�_X��m�nnl�o���S~�0�<]����ަ������Ϊ�)�ӞSv���V��
E���w����,�6�W�R���������Zױ���/�I��?تo��[K�r��2LF]3���Y�<x�{�{��O�����:{cp}x���dm�^k�_)��.����o������r#qu�hy�[���Բ�\�,�>�iw$�:~X���������:eul��.�m��W�ڎel��w�_N�N|��j����^���iG6��U�v�c����]�����Օ��͵7��=�����m7�������g�Ϟ�9�'ڬ9��� �f_9�L����ӫ���jl	)�4hլ,����U�k ��We�oŔ������u]��l.��G�~�z1~��O/zG�ӓ��ŕ��6繣�|��ՑU;o�q����'����5�{�����k|�<;�,{U����w�]�'�]�߹���]u�_Zu
no�ڥ.���o����fg���;�6�+��X��­ݸ�kL�5�W�N��flhN�䒗q�XrU�t%?��L���ʧ<+I>=�M��0����a]�p�d05����.ۂL�� �RNu��
�LBC�A�	����(�H�CB"��/���?��L��˿�K,�˄P�AWל��2&"�w�%0M��!�rR�{0I��3fM<0������?I/J.���}��}'oMu�O�_�X l|ps�Z��۽}��<�iv�V}K�"��؁�վ�䣟$��U��՟#��M+���Q�z��%?�����`,	�Xw��~��$�#���g>��ԙ�O\<�K��ܥ��¼�1���|���A�2_�o.�B��/�����r:�w�*��3�M'`c7L�%-�s����o{&�C�����*\ 2�.��ȟ�>���+ez���Z���Gh@΍�:�6�/W�^��?*Gx?���������b��xtp6s饺�k׮��&�-Ű\�U���6���o
/�Й<z�Z�%������Xqq�+W'aP��ZT�[MX�.ה`j	��[�[zx ]���T¬-9]�Z��9l��X��	�]$N�2����7M���
=e�L��Y��ڰ�J�L8��춉��fK<�$�9��f�m�.�/BV��kG���<[E \�4I����pc�����)��1�婟��N��7���s��-W��ϟ?�x�<�nm� �r1T]{LST.��F��&ZaX#d�d�@2�3|Fu���z�h�7']"�%_<����/ H���	��z��Ɣ6L�R�e�E\��� N�0r 91v ������=}�T<���BOP��H@"	�Ļ�.C�^���7�lǼ~��F�;+��8_��%y��l``+~����%4Yٸ0�T�5�W�J<���������?�d�
%a�R�i�7�LB3*��d"T������l�]�0bPd&��De�Xm ��Պ.�X����,�zY�G`�0L��LH�6J��6h�ն��S�L�r���^V�I@�Ɔ%_	�L/i��.���<��|z%���+�`Hϻ��JF����	������FWh�/6�$q��#B�� GlQ�$�� 9%C#S��.�2��b��YW���.��АCN�,f0V��R~�h��'VL �BA0�:�I�T�G/}4��E��C������Q�¼��Wa�&�^çᅌ��k��ՌFm&�1��2�I��ƅ��pT3g�kB�;
M]l�CVІ��.`B�%Cd��b�Q��.L���e�������&�T4@�/Jr��r"T���L	F�	�
�_!�V�S��R�5<XzՔ5a6d4�}�0.���R!��Q�+a�,̐`s�	^/���h��E��B�pY{�i��Q�ѼJ��A�8�N4���	L���,�lA]E�ܾ�}P�&��m�E�5�D�)H�����&$s���	��Vѕx�!H$4�C+-�41T%~�M`aS,B^∡�0a0���|GЫD��]� �D��$���9-${f�S��-Z2!��K@�j�nM�ԡ2@l
^t�׶el?�� ��6���Wh�0 ��ģI��`,0$Y�&���NzX�
9��V�`yd]�LY;�I��E3<��H!_`j��8��0��k��&~ �8�cC�`@��>c����m���1��
�>xJ4A&J$jl
��)��V�<B�/L��dHJ�L��
���&XUGs�ĆDX�ģ$Q�q�U3�4�:~�(E�&$f]1!dt�hX������^ӄ'pJPG`(zʚ�m �������'�c����(y��iȱ�,
AC�r�c.�c)bc��Hll�=V��0	+2Y�-�.u\0�mf����'�4������8�i F�?�_N�1�b��#D�p�<zTJ.ޢ�	6����ob�����7�pJ��F�@�OIf=�PՔɭx��SxV�;�UH$�2�Q�@�W�F�@v�F�I	Ðw_��Ph�4L00q�f��UXE �s
&#M.����U� D��ŵ^&d �.dJ%�2��2�K�LM���� Q���PS�f�Ï�&Y��l;"�,�
���c���<��� ���
�J� &~u�	�'���I4���T#�'��Ư��	JGΐ�H��S� �F|^pe�b���]"�ψ8e�}�k����b���wz�S��Z��3�:lp�nF��`�I�4�������ݾ�W��8�/N�G��N�/~�I�M�<���ư{r���ߍ�WN;}kz�n�o]�龿�ybl��f������a����>�Ƀ�����v=�U>�{|��]�]]�͗�6:+e���66��eUY�]�L����������5W6ݕ�	�{����.������~����ɋ�ȫ������ach�7��?-�lY���Bߛ�F���l2���SW׼�����Ó'��2?�1��qϥ�''GGH;�uo#u�����Mk�
i{e}�|^W�=��Ė���V���vi���<��q�r�v������d�P�=k��-k�]�{�3�(NG���ז��߻�ł��b����r�ko�L�g�_�^�zB�(����[V�c��ئ+����n��&�o����騱�큣IyBo��\��VW|��|�rs�ӵ��Y�r`�`+��lMʾ���R�e�����ā�߲�WvaKJ���B5����9��5zӁ�2GZ�d暧�0u���ۓQ���+�;KV�Zn�{������7�}�ţ��`��:��ƃ7GG_�p����n������������ׇ=�>�Mۯ�?��?}���_��^��^[�f�����������CZs���\�ۓ�|��89<�8�����NϤ6��pF
�kq�<ֺ��i�|N��W+�V<-�o�����YE���D5{p����ޖ۳ִ������r9�B�><h6�׺�,E�x~ptx���/^</?&Xn��.��o�&��=�Ng�٩�SҪ}����	l�L�7���ʑ0`V9���i�;�����#�cv�6Ӳyf���Ҭ����nk�zͲ�[k�V2��g��́��Z�hz����ˉ%E?5�6�vs|���{�n,w׺띝�={��o��ϟ�Gg��/~����ho����������o�:=�KV�=�6�~m��fy��+4׷��ʺ���	d�t0�ҲRb����6S��m1No�qɀi^ffuLKNrpK��}�g���� Gl���!z��hP�̕��7dx���į:�Ho64ͻB�յ ��A�6�aN:�dJ�\�N�* r��ՙ	��[:�x�ǁ�]k?^i?��8�=瑛��@��t
�    IDAT�&}\"�? �Ԋ�X��%9ӑ&A#��@S�ˡ�9dƦ���/��ei�/L�rd�`��чo^xZ�ݺ5��q��`��`��(e׬�l_@��R!� ԉ��R)���SV�����wu�=��>�.�1���y�^x[��zY�{S',+���@l�v��_�F�����YNL�e�����<�Me��˃�3���:%�NE��ns�u�X�oD付�孼6��vy�Y�̮ji�,�V��Y0Έ�����NE�78̭���=�<�)M�ml������)e)�s�~�R~���9���p~�[�x�����'/�\a���[a��؋l�
������A�{u�� MC�|���ds�V�ܳ��_]⬒�F���AE/����M�L ��P�ҋD�&��d��5kC�vzӕ"s�HJT�+VH��&��}JM`B��Dn��Q�,{��\�ԫN����]5e�_0��rEP+��ܹc���"���%h�ٺDV(�[��Z�$�%/�9 c{�u�̦����䰅��s�� '�'
�E���U����2@�q����-��L��������L/*GIGH�M�yJ�p"�p��݃0�M�� ��x��a")1�W�dQ�dJ�4LN�ɧ$sW����G�&3����H���f;N��5+��	Fe�ǌKhu ��1͏>���Ud��.�`���!��ݻ2ϝ" ��Ջ_�	�8e��_�|�P0rh���k�~���Ab6���a,��db���/��ՄD�4�^��-��ZSr$?s 9�O]g��ԽqZ1����	a��"��d��ِ2Z��Q��zVI�XI�zi�IA��(�����Y�"s��0 h!��4ɡE('��cGˈ4 *lx֥��LxE�)5��+Z�_xJ��`d�(2�p�#T�t��Հ�h�=Vz��c��qQ���-9��i�jl�w0z���O�� 5@ʿ���	�`��a<
	�h�	qIU���'�Q���R�V[I��" '�l�8R���EH�m4�f2X�7�k
#� Qf��A N�`����jV1�n8 ���vD?�^��X			63A/�d�D���Ho���Ȑ8���	�M�������C�P3�)534A�I^��S�i�0'�4� !H�0g ��ɯ.2��dz��GI�	4 �$�4�..��e��c��VƐ2��9���d�L���1�����nrb��u�u&�f&AIHj`qbΌJ���d2�`�z	8��C�7���dB���b��Ec[�kM�\�B � ��q���:?AF�Rl�`�0^���T��d\zE��^Ͱ��4z�B@(Ñ�< ��\ÊI�C%ʤ(���a�<�фJ�l�C��M�z�;+���R�D�fl�O*�(i���4$j���-�A3��y�+�H�,N l"?������LTl`I C.���"� M5}���EVS�&��,0]\�9�梥$��2e�^&A8�X�(��*и�
�KB��'60!�J0 ��m�+�@���+z��J���aRfF!L����S���	�.5X��P� ��00�D�X/�����F�����6&�C�Q�EK�ӄ,��
U���`�3FB��C����`�K�dJ<J���Ed�a4i�����d.B#�L�+%H<ӫQi³��$����#2s��f+zlqm��i�G���_a���	LZޅ*~cE�7a�)՚�&� d���Y�qAP�P�]3��LfX{���8�&u�#�|��<�����BA�����0 Tz�G����Q*�!C���e��2�d�<��d���$�$�	L��� $�Q�RJ�l�g�0��ː��I�� *�A͖S��4�ÓӫĖ2]Ƃ6��&	�&*�jށ�3����T(�u�7�כ��cCC�%Q3�KC�����3O�� �ҫ+l`���FO�.y����!��կ )E��e#�0*�&����K�WH�3�ĬV���fhl��M� �&x�μ`���� 0%M����^�ڌR��a�q�DN���� f�q����Ϟ=sU	,��=??>?;�zm�|ڮ۶L� �v��^g48��5q�iwʗ��.ͻ;���ۻ����7Y�M��.-��#�H�%_��ͦ�_���6��@��EsٍX��Z�Z����+V1G��|i���-�A펫����8��.�2S�ܨ����0���<�9\=����T�����o��߱�5�\̬%w����l�Ͳ�!�l�fyg���3<���^����omZ�]�ܘ�ʒ��X�q{Ŏ��R����2f�A+�bշDl�pҰ�۠\_�*����Ճ�����O�.|�����?���~�6;ݕ-�E�\m��^��N�sO����I�u<�K��Ƃ��r������,Nz����Ϟlo�޾��ޚ�}��zʇ�\��E��ꃏ��e{t��2���Bk�o͂�����I�^{�㗽����M+��设�F�\�Q�L�*a������n�ۨ��|����O�=|��?��޹�����@�W��_<?9|e��c���ȷ?������6������r��^�c5�Ntt�f2�^�>y)�]/���/������0��lZ-�Ts��4�Qgiuyi�xV,������5��M�Q�s� /.̗��fǚ�l8����֗B-qW�����Z����ղ�f��S���Skx1��o~����OT�x��rxfq�ފ�}<�O���}S��TԞh�#�Ca�9 W�,G�(cB��.�����0��).����YV�y	LBUM��L�����H����kέ��]����ӒW����e'�%����|qa��7F=����3d�}dpu}Л<}��Ӈ�|&v<��n�]��~���Y_�~��������wcw��j](v6�vW;H������Y��l:�W!;ڡ��f,mV����'y �,r�^�$�&�%�#�s=dRWyx{9\�B �[��B�P]M� ��f�#���k	 ~�l����T+�MQ1WX��`N�S�9��w&��������_����'|�w���ǡ�\7���Q�RcD!�xM����Ա"�1=�fj����F�Gm`��ix$�(��e^_�x����=�E�����F���c/ϛ̹)-�O��@�~�C�,{��T�pQ� ���:ӨKlcU���r>�9xV�?wO�uMq�_۔5T�2���	��n/����|���zJ�;�I��J�c�xZ� p�h��d��qw@5Ä�g2>);�[����d���J�%���S�TN`ӱY�	�Q�\�a�M�:�,\��Du�r:�%a˟"h�Ov�c�Rhtvr��]N·�G�燽o�'�vg�\e�e��F��դ�0�H�ĊV3� �����(��X	�C]��d�!hb@a��]`�=D�^�Yq �LY|W��(;6zz&��4�F_2V�9uU�eD
=��� �!�p������lw�,�`�MB��5m�\�1�p��!O�7�b���R�9��ktw�����~f)�;�d�	|�;h$�)�G�L���*�Ç]\:Έ���Y��?��`�0��j+.9Mzb�\�;�)���T���JdpU�o���K�� ,N��S24"Lxf�0����+yf� ,#���z���c�9��q*I��C��2&Z�T���8�
R�b�;�8�"�LqE���WHk�H��Z`�B�ӧO��
���H��>s�>y�#C`��pd����aȊS���Z����6��Gȸ��JBlDuR��A�����4^SB��Z��4�l25 ��ɵ�0P�'��I�	,r]�0�p:�}���2cP`zMd�)C�I�8C�D3r� 5�1g�JM�tţ&_x�<Cꪀo�H���0��S��Q�5��q�ŠKɷ��i�����(ԐjQ)`<U��c��T�-w\0)�U	�L�-�8�/^�
SH�Ј9!C��0a�Š� eFA�$��TF��� �I��R�I]�K%B$`ƒ� �����]�hӋ<��u%Q�Y5]E$��D��ޔ`�ũ� ����Q/�)�\�Ѭ	#�K�9 [QE�J�bD�+ 
������	s ��h�'lŲ�F��g�d�O��Ԕ�Q�OW�
���-�%5����]<9l`� �F��{�'�� �_N��֙�!���~���WM�̐L�2|�� ��&2�^V1�@o���2����;m���<���,J�Z.;�P��t}�~SvGwt�K%�e�L� I8`��|����FtuRJ�\��g�v�}v��G�d�dŰ��cK	CS*N<�� @f>���a��Xw)2��ge\���T�ކ�wUrJ�R�"�dz(Z*��%H���S-���gU��3��>Gi��i�(��a��碫�g}��́�U�|6�V�
Fm�%�(�<���6���Xz��5�ȣofZa4������K#w���04R&<j,+��;0�L(+�aN�@J'=[E�4��Kb���\E��2V�fv�(��	��Ө�ќ���� FC���%�R�����B�!�)� 	�k	U�f�b.�e>3P��3ǌ͠p���pF��@����4fB�jU�#�|P�Bf��!~&�4P�VK�fL�R
Ɲ�;Fr� �\bö����2�y�c�B2���/��D-��%x�����z����%���s]���.<z�\R�"b^�Y�H�*N �)�3[m�� �V��R��!��D��<4U}V����s�b��a�e�B��3�!`�h!�'�7p�-�����P�ARb+f�$�ɼH�%�����1�A��H��[0$lk/�����E%�1�!�@�G�H�$�@�*�P����/A�W�g[�/��(����P���mw��	p�>�����!��x\k�Ǜe-�I�	&ߌpR���%E�r~k��:�b�ܕ�T�P�.E"�P�ϵ�Y:ch�:�&#DÜ� ���h#V+�.LEH��Г]ʫ2����}.�,�X���vk�0�RB��H�i���&!�u��rET��#�G�� 	��1 醓_U�*0-��6�H�x �J��c��£���H9�^���H� l#T��rMO�iܱ���hL�`
��b@�詑`<e�(@Hx���hX	���A"a8��!�/�󃚫�8��a�#�6��?\���w�~�r�磅յ��c��������ʦ���<��s�m�zi�z�����޽��usŮ���7n��^x���O��T$۫�n��tq���x!�GGα�����R^�j��k`�N�x?�X� /��OW.6W��/_.��-^{s���ICo��Y���W�����r�+^;���>=��a��XίO/��S����6>�Vםi���i�Ns�@�4�����ة����=�>A�)�'x:=�����r�4Y����r�����_����w�]/��l.�|�̛a?��=��}������������#W�J�A7i�]:!�����y��h��O�f��������GWK�k�F�M1���˅�m�V�[C��?�:޿x��x�������#��=�;9:<]^�8��m���N���C�p�Bw�����<�w���&��ʱ�,ҋ?�x����'k�;�s�׽���t�չU�� ]������~xv���4%��r�l�Ut�n,�9u����ڬ������8��+{�Uk�+�Yz�}{{���1_��6QF�; e3xz��I�*p����޳�����x���&�qRI3�H�y�#$~���j�;w��l��������/����}��C��^���ỻ�ܲ���Bgrz�h�]��Tn���AoD�T5�^0aP�f��{-`T�� hfBJ�h״"�����c�cY�\��i2sU���\��K{��}��ӗg�vV��Awf\_ݲV�_�����u7�
�����?����\�:�u�S�O���ؾi���|������֍������Ѣ���ږ)b�5��j���zk���O�Αk�$rϤ)��f��|�di����0!�ؒ��c��K��C<1��l9�Q�m)!��D�V����2A+I0rJ��*�	L# U��3���R-+�uC��`���M� R� �so
6&V<���ڧ���=h��Ѧ�U>] +2�	�V��D3_�#����k�qq3A�Amx�F���	6J��*Ef�(C'ؐ;?;|���3�����������΂��3Ǆ5������.^v��Hz���"���/<9���|�ri�G��m�M��"q�s�3����)��qI^;�Ƌ]���X�|:�Y��w��Y\[���5�݆���+Ū���VYծ��8Lj�xQ�����>lx������q�� =��<>�P��a��������3�+h��1�{�-��<�XǇ/�βZ���aw����鳓�O^|���ӋE�>����)!B�����U�h����t[U��$�� &%+��0�*V	�qaˣ�$�ɰY'�l� `��$�l�a��+2�DN�L)B2/�YId�R��o�D�e�U^�g.��K�r��S�]_��s�G�Zf��CQ��M��L���v8Qgk��3�LN0,C�<V��K��I�f䶬�,�ic��*�ل�_�C0����-=Jr���SUx�̶�`£]M�v��Z�P��B��_�Z.0J��T0r2*�c"�����W uT�l���"Tţ�U_I ́a��Ky��c
�!FC�l1�Pu���w�	F� ��˅�.<������E��C���?����$����Vb�� �h�8+$�c�A̺�ۗ_~Ʌ�c�cd�$c��l�̇~�]ru����֬�D�4�Zv[���j��~�;�pʵn�����<��W��tm�{>�#�y �͈�#$0�
aK�(�3��e�
��"$C��j_x1K�`XMdca�XEU���4����1���JQ3��b,hXI ��?�\C xQ�^��>A�L�xto���V1��Mm0^(%�r0 ���Hq��Z�YSxx����X�L�3O)��r&�d�M���2M9��3�dH��#l���#�r�<��a�`R��I(Y�ώ���¿�L���L, z�� bHS0d����h�i�	r����V'�	j	r4�g�Z�
�e�R�G3`L��v�����V$���◬z�LS��Rf+}"Z�H|�Ld����)���KUzU��h�y��
�-!���DH��R�&c�3>��Nx�V��#��KxY�VE�I\_����C V�8U,�T۠����\�Ix���R&0r��9 ��H`C��%rN1��(�II���$�+�
R�D�U��X��( ����MM�v��3Z�H�*A���*� �&�D�6BU���6��ATŏD��$�"�-�4�ţ���s �G3��b")攜r��#�	f�:E[@B©D�@���IH�y~U��8M¨�L�c(gB2e�f��!fJ<�Z�!�b��.N �����^�E�	���0�뷘߮-ȂA+ ��C��K	O�h`⟻H-�$ ̐|��'H�Q��� ���N`�8X&r.� �[E}X`����X�LH�̐R�����U����Ʀ�&�&~�s�&$�	sѪ�8�^Q�-5�B��#G�
 �:��- B��2������&~0+<	 �q�H#A�S�q�S[2aٸ�@.XQ0M %/���q*��/yH��p��F�)#�N����*��otVx �|��3I�Fj�&���<��y�ϼZ�#�7�5�� l�fG4�f�6<�Ĭ��$�b��@Sm�j�&�K�UI���<=êZ|�J4��9ͯ�Ġ�{�D �HU�����._�_m�(�$U�攭��#Vd<��'��.�C�*6H�Z7{�G-p�������b�b���kTz�.R@O#ŏ
@R�J�x�R}���/yTr1���L�U����LC��У���c�`n{�h�G�a�jY$\?XJy�YU�٢R+OiF�V���j�U39���&�]Q��VqnLUa�|�    IDATF�����Ŧ8����E���J�բ����"���g��L�kM�a�J�u �����W�P�/ �"��C#x��ECϞ����m|xL}t���s����?�����wϿ������y��[۾q�ޡǣ~���sQ}g���*��ܽ��'��[&���K��k�'~:��'�|���N��;[�ݻeW��o����$�J�?�ٴG�c��b��ۆ�*�4��A���0NTzb챮ѕ錢C/L�S��iq��y|X�cON�
g���s��{/�q�����+�����Y>�Wk�v���F������lK��`쟼|q�ի�\�j�Z[G@�{��������x���㽍�]O˗>Zٺqsqm˝����έ޽k������Iጝ%`(���;ck���o='�\߸������|�哟��s���ں0�>:������~�YXܴ㸹��ѾG��+�����_�\�8��h��읝k:NG�����4�lx$���MOu�m/T���jw�~����Z�c6�O���85ކ�A?�W�n�o�/\���N7�� ���ٲ�8s��������6�^��x�n�ڻ5w�F�ҥ����ʼ�\:;:�S�����;�n	���Jn�4�ԅWF|}t�O�2��[���Rբ���]R����H0zv���[���ӟ��߹ss}w��������gϝ?y����n��~���q!/�gn�����-�P՚ :P�.��щ�%�eB�(�'�S�"�O��*[ݨ
�4�Ӑr�x�V���=v<��L�}��Y���~K�������|��pq��+�`[��w��{ׅ��������f������r{m���������^�l-r��沝�9��9>�^O�Lk�xĪoj�?�'�{�h����N��]��œ���-_��T��ץ��B-C̭�j	�ݘ�3	�r.
�����"N<�6%�;��"T���#0*��UVLhz�
\̳-+ .2;�ʧ �񚯞���<J.Rq��ٚ�c,�fO�aU�2��RF(8�`唚*�r��Z&l�M{�DѬ�S7�C�'�W?��r��~ea����ʮ�ip�'������y��s�q�oX����N��OTL-{���;Z2��w�b>�8Z}��{l-��H���~9�K�����3�k�V%w�P���ݕ&`����Z1������g&�����ǣ��2����~�\�+�5�јG���j�S�j�UW������qL��&��%�Bc�w���(��� \�>UΎ�������3�O8~���O//���ϸu����Qs��7+��>�Fm��t�E7��A��yٽ��y�D8��X��^.��NW8`�T5�cN`��#9Y�@i�*ʣ��*b �H3GB(�� ��NoI��CR��`�4�x��z���e�e�E�=@~�)ӫҽ�Z�,�@�/��\�EIQ�E�;a��m�V��`S��q.U�Q��b@�3 ��19b�D��᫯�����<ف�o~�<�� P}���6������.*<���Td��'���L���m���|Y�8b"x�&$���f~�����Cx<`桽C$��~��G��rmgN>�k��tE'M����.��i�樥gkX�*�^%ШBH&@<-�9Щ��k�+0����[*���駟ژ���/����Ń\�!��\�2d��ïc(Z�_�x�1�5�����b`�zс"�
��Y���l¨?�Z$T��c��n�G���v�E�i'E%H��*���G��W��ׇ����D$��/�G�xqF�����qj]�/mT��i
[�� % ��8�|�KEŊ/lh	`�U�RKO���`�s��! A����@x�?�D�Әk2�Z�*�g����*��C���	d��dˊF.�����gĊ�BU`1���fE�,�Jl�%�S�+��ڐo���j#�����
'd$����	rU9�$��K� ���R���K�b��^��9"ȋ@1��s0ю>z���	Vi�d>#a�a<���j� �e �rM�o�Ӌ��Fʼ�(b�+6�5�b�a3MZ���a�E��A-��]�R��p�0�R��Q'�`C��F�Hy��X�����̖� ly�KZImE9��:yQ,N^T�|T�8���)yD^m!q4L�5@3A�E�5M=��~��J��w�\��6p���?�3��j~	2�d���-+gG���f�m�XA"�G9�s2<�Z�a��yQ�#�5S�3Rf�`���O-dl@.$U��c�a���b�Y��MN)ix	��.�V���`����PJ\?�8�W�*�4j��H��H��G�����Po�K4�
�0b+l$��٪���RQ>7�-��lUI��"��
�>A��`	!�ZJ��V4r2f �:�K��a�L�	HA����W=@��Tq1�����d�V�E	I��!=/�җ�A�K��Q���U��'�8~9�䨀�4�:m�A�0A#�gB��/Q��;+&Rl�$J9eKY�-ʙ� <��0�`�	�^$�j�~L1/	F$r9+H�s���Yx!�髪V�u��!c��u�ERTlYM4�] [7�-��j`9���2G���B�7jim� �w�.<<4�	�l�!J�H�j�b����E�8k��DI�e^3� *z	 G�J�(Z!T�h��Kj�RK�ǐ,G/Q����@�KJFX��=F���%� �1H����iBR$�b�*� �΄��L3{W�3CT���b�"��g%$6�xbCe	�H��`�8i��4`������0`�� ���
U���8�~�����%�Z��\��WK�<�'�����$�ƯV<�3O�x(�H�j#+%N��d�"�$�Z$Ѿ-У�!!rT����P�Ө����F�L�-BrzU4�y$�/<r����R���ƒ56�O@�}��d%ZE�A�5~�*R[�L/_��
��0 ���UI�#�7�e+0� �<�ȁ�媘gr	�R�Z䛾�$ȭ� �p�<L�@�F��=�������hΟ�z�y������=��w?������k7�~���݋�ݭg/�Y�[��ڸ<9{��OϞ;�v�O&m_�n�,�±�t|�L����݃���Ǉ'Gg�G�_<y�w�����������O_,.m,/٠�۔�����k�ttݕ7�90�=�����Ʈko�����t�x��g�Ӌ7�Ҕ�۶��ۉi���.���Yl+k��p�z{u������2��v�?on���C��^:�9�ؽt��W�/�Err�y�ӡk&�"����G�G�	����ի�������ڀX���^�8��Xs����O�_z�ʁg����$�K�y�o�u����������M�gv<n]������<^_X:p���K����#���|z�1�$��������#��i\^�o�o��W5DO:,����{�}��K��`�1%۷�1u��8]�(���+k�;�^�;ކ�ۺS���sNk�����ŋ5��8��qّ�bwq}v<6�Ϯ��>;&��~}���\]=�r<�������%�'�3}8N^z�䂟̼t�s�B���^_����z�e�qˏLN/��Ntm;Qr�!+˗/^���o�X]9�q���O�/��o>1{~q2^��4ܾ�7�� ��a���h&MW�A![�}4H��
9�N�3ɬF��G��\.!�Z3�lu�\� I��gŬ���Y�;�܎Y�x�^kj��������g�D]5��f������g��X�ƅ����FEZ��;>_����76a.VN\cվ�ĵ���=����EhIs����u-��Szi8���`4�<IK���4\UV�dJU�x�	��� ��$O��ۜ��;[q��U�`c�u�� 9)��6��B	�#�* `�05����*�6u1 +RFB��A����������Iiq�(\N�V�DDQ3����1R�qIE�{�Ð&�"Cl����1����8�2+���x���!��QT���Sq?;�hbaq���\\�z�5��t����bg�Q��/XH���N!���oU��d� ���ڊ�|�3ܗ�'k�r�r�U|���;�ZG������	�4K��oj��CG@�=C7j6��R9��π�F��ٵ4���h�4�\N��ݳΈ�P�Z� �Cm5�,�$VU'�7>���gG��߀��y\��q!5}���ne�EbB���'^�;�C�V�K{B�ώ�}�y�~����/��=;[���k�p6�Z'ZkbJz�15t��Ɛ��<FW���Ue��ؽ�A�j��f�1̄�b��H��R͝.��Eӵ
���#��6�i�P�!y��h�4���F�N���
�-9���P�pZ�a�b��H�0��zF�%�\�%9%����SBb�+�R��WT�Vm�4`���J�Xc�!R`��#�Z�EG�+�Ca�r���F�/�K���Z	���7�|���6����7Ў�����G#��'w��"K�`���Qp��]����ܒe��	r�05G�m^0[�w���k!aV�P�D��E"tǬELS����B�f#�����F��Ɯ;���ga#�{48	j
طU�x$q� @y�A��\���!����?��?b9~9�8mOQ�X�1#�m��֠�h 0�%x�*0�6��}(ԙh�B#ȶq��?ZQ�������*�x�i��'kI���w ~Ua���6��c �!�,��ZA�Q���K9E^��?�R��$H��Rd.�� 0�f���
#�4vj[L,)2�#&��R���4(��y$ �L�p���`5GE��!S-����S<�PM�Ɣ�ܢ��	��(�Y.Q��r'�ib�K��P䊪���r �J�F�D�? [�P��E��M�]3�YeTj3Q�Ez���U���7h0$X�U�W�l�FCOS�9}��0dQ��u�j�9�<+�����%�b#�d��h\�NQ�H+ɼXi���r�S����4sRU�SεsC�Jd�;��4� �\(ij,X�	�@�ZCȦ�<�j$Cr��\��$�:��e���*Z0��G`$ʂG��FNY��AQ2�]���\[�b�Q )��}�P�x!�!�)���RÊ��^ EȰ&Ć?M�y	6y�JS�,�!L
��`�W	?�&�1��c�#�ڹ�:J�%����?y�[�+F���ISHr��W�p�U`�褉
,*dJ9Y�$2+��"=B��()j���L�D`Ud9YUA��%%s�%9�x�P
 �x�L ����02���+���M(0	����N�^�0�x�.��c2��U���V0��E<d����El��a0M��H0���;��J!�0򪸈Y^�O P%�A�v�;wA}2��#!m�	e�iO�R��Q0:� @�#H�)���#Z�1�}6Q +}�u#�#0�d�z�/�&��%s �L��D�<�z=1(���(�K<�39�����2�"�:$�����c���(��N�#��y0��!!sT�&fތe�)�.+��Qa�}E)~H+B�&<=e�r�1�L���_y�г p&4�~��(�� ���R�'�) .j5 �b��A�8c�LH�� ��M�r z1�i�*� /�£�/�[t1C�X 02pݢWkrFU $�Z$�VC�bC2+yBU��H���dĀ�ae1�E^00F'�z�ݵ�i��bB[�8�P�ë҇�j)�<�"�۵�)�P�J���0WT57�G-��~.� �hƮ^-C�
�,`�t�4�����j�jEҧ|��r��zq��,~-�� �R+�2�`E`�9N&�Y+
	X�F�k#@E�.q�=��%������FW�4`X+��<'k �r�h�i��0�gE̐r�Bj� i�u/<�x��L ��]U�P�)	�ImJ�)w�%τ	�R���+�}UH��7a&4 �_�gNC_�h�*z���Bk eM�' ��� �:��֐F����5u�s�ɯ�4~�1�7C����4�O�b_\ݼ���G��Ö�+�k��W�~u�ٷӓ��t�y�l��w���w�.����mx������������/�:_^�\[�O��N�~~��a��^=?=�����/������<��e��&z��9�7��-Ho4aq�[C�;2^��ě֓�s_���xƽ<΢��1gm�Zu�!|�sm�g�Ci�m�p��߫�@��dO���:����g6�>c�Ű�N��w�u�7>���ᧃ�{�>x����ݻw�v�V�;���T8=��p$�уo>��"��i��j��������ӿ�O������{?>��K���߲���ѣ����g/_�-;>g��p�'��������5��.I�͋K�[ɏ�lc����5�Oi��V�=��/-;�H���$?B9����Z˔�y�}��{c�o��E� ���q�qF�[c�T�ɕG�Kf͝�W�]ܷ#�p�m�����.�ga����ǂ8a?�$-�5��͵{�^3鍓�����2?���޸�@w����[�.��q����U�齭joO��>�KN����l�:;823�<بy�����u����fl��_����cg=זWNǏ��8���׎/b�v�r��?=�櫧7��{��d�_�����?ܵdt��K��z硫�u�z�DKGGOW4Y����u'i��An�t�F[$�LȔbS+NnA SD5:zZ��(�w�O7J���a��͇r��}6�{���L]��7��	V���O�6>�lr��$�������e�m/]{�ove��r��L;B7}KG`]��T<}d`���g�|�U0���<<�\ij)�4�X�����!K-��-����9�aT�
9�\��h$lME��c1���>#T)��#1Fr)���@J�"����ᘞ�(B�[��E��+V���FS�[�G4�i+�8]��W�����O���H�@�g� �Ȓ�;6�sЄ�$�$�9z��O9'��nd���魼�ٺl�j�^�Ҹ	hD�f/�ig��̮����ӳ�'?�����wW?۹��a��ۈ��Y�V1�����x��E��؄VeH�J�6�6��[��#d<>�F���_D�A��Jt7.����YYǏm2�χ�X��|NO��P�/�op�
�zf� ��9��<��8�:w�p�I:.-�A��C,�.i��3�cӒ�z�52��:H�_ئf�1)Di<����{�_������׍���p���c�'�G�<:��_>[�:�����x0�B]3�hW�q]4]��!&�'a�ӛ���,Š��X�H�� �f 6�r�8V�yWE#<ł4��)1$�� �mKVC&�A��-�"6Ţ��
-|� �4��̔8%�i���ҧp���"��Q�̼�Ӑ[S���ŉ��0H��؀��ݯ�Fe}�t�k�iN��Z��"ᗉ�����B���%#λ��Wm�E��?���o���,;����S��l\M��P9���;�(�b$~���v��UUż}J�a3�l��e��w-�<z�#N�bh�-ٍ��ytK�Gⴰ2����V$�k��9J�N�@��y}��-��@$�%������Z�J�;w�qZ��t4X|�qA�;Cah�x=z$�FY?ۚ�"�hs�׫�ă_�P�C���_j�4��t�"N�CC�P��b`�*G����`�1?~�^�(�R���/q�W`\+�o>��j�b�Wk�ܰ~��xĠ�@
I����`��k�Z	���@�DQ���	CE9r��,��a��9sU�h`T!��-��1�		�U���JZe+B�0�l�
FfX�4�J�%�$m!c@B�����AQ��[��j6���Y�\|����&h9V|T��	%�lLx!��m��OYl����� ��r��2�r��"���+f�D1��r$!F
�2��1#ל�����p&4D[`U1�"�`j�2�$/�p�E8+陇�cPe2�/Bzm���	%YN�! ���`�ܕ�e	�T���@-�)Tm2�ϑJ@    IDATd$ V�>�3�1=@� ��Y��l��\���Y�e.w���P�L˪�e՜Ð�2�+J�pT	DB�J�R���e�uT3��J���b�A�AB�:U4����l��dkb�D[wY�-ڿ��oE�ӧu	L���E����F���R�p���0�a���2� X�s�j5e���E<\cH�$�èU,~J��D@>�������&0g���ɂWd�z����
 ,~E>w�"��y�/B�9`T�����Q.2�(��h��O�R�ɗ�z#C9/�"!�(���k�|����� ��K��S�V
 �~�(�Z�Ɣy�l��>t�"�/N���DC?E7�N�0��	\�8� �&�֩�9$���U��C�J�3��=6)<ZT�+�"c��0�@J�j��a(�R��b����4���fLHBJ�8ax�Α�q#:�alh!�%d�9NݨHY��3 �M�QG\ ��R�֚��1$B3�����k����̜`z�gԇs�T�ȑ�K��I������b�
 [��ϜR�wJE$��r&țr FD���4y�QU��l b`.G!%X90���S�(Fq���Z�����f�Dms�\0�T+�A�DB+ ZE�0��� %Ū*2T����Ŗ��chQ�Wd��L���a�X K�^m/��j)�Bj,�%��X�3o�rJ�JY��ls��9~���%�@������C?�D[�W�����ih�`���#���Tu�e��WԊP+���Z(�p�X��LT�RQ"�Ԯ`��?e�7�� ѢB�K�s
�Y>�V59Y~1�V��cSE@���MTSh�Hj/����0�Tqa�T�-�ju�"a0Ex��H���ϗ?/r=@��i$��=�?@U��J!�]�4�0� D"�K�K����-A�_x�`V�"!�D�#$��jPO�orz�"g��sHONl����91����{g=� )@ֿf�����<������+'+����o�:�s�����m��{G�;~�skke��=~���֝�?�lysgq����6�ϷW/�
������+���~x����ώO.�����N\�r'V�O��6�>bpF۝��f�WJё=�G���t��m��?_fE�0��n3%�gPp��6��x��#�F�����_��_���9���9sv|���+?������czO�����}���������]��>�.����ZWc�����~8<<�v8���b��Sw���ݍ�խ^@������ΦsF6����?|1���'�I��\أ!~�t���?����U����ǟ~x��;^3k�i��ݻ�s�j����{�J�������흭��G7������Po��-�	+jS~}e�&��Н\��]���^\�����{��q�h��V��~�t��챝�t, >}���oF����Õ֍3��-�����u�<�x��Z�koGrnX������%�V��7�<=>�:��l��F���~�G	�Q>?]|���������������§���}�:�k^^�i��o�|�������ݣ�G{|��G��������$Ѣ����g/\D���ٕeIGhf�V1h�h˴J3�ZU�ӴTE6d���3���zx�� �W�VA-�h��'��Զ�[�0�_j�=�'�m:��i��k��	�u��u�s�¼��2ч�[ �]]L[6�մ1�<��B�qoe_�hFlf�8�Q#fI�L.~E��ɵn8ysKC3��_3��L�uZ�V H�j�T�q�1"����Ԋ�O&s�*H��Y�UE�s<�)�`��P�[���aqN/��I�Cx`�����Z�����Q�"�-J�n#��a��	��N�4}h��4��ȶpY=+��b�K�*zr9CT4H��V%ћ|�d������H�8^��y�tl{�<<=x�é�ji}{�ra��jᆣ���][���d�Ʈ�=D���6jAiT��Us��Y�q6N�͟Q[���-�h�Ɏ��!G��*ƌDn��P�#�1�1Y�V�ܑ籿�;펎3����il�N�Dǭ�^O�X��b�|��ua�@�/�6u(�ժEc�ө���C�ϼ�:6n��=���j�:�p�N6wu�����S��y~z�����O?��?���7/Wt�_�^����fj�t�k� u��i��O=Lc(�2a�?c�[��]0M���c��L�&4�F���ih^_��]�MK�i %&4�)H��Ȗ�ZT+���k!�hg[Qȋ�!l8)�H ��@�<�rQU9l��X/hf�p��Rj! �|�tfq���@rQ�!c��]*s���aCK�F0�x���A	B=`�]g��ള�Ђ#w���H���
s|��wH���G)�/~�ˑ�}�2t�)lO.�9[sj���QHj�`��Ѧ 0+O7��y�͐�R�b��/EHϜ�S{�8�����ƺ�R`j�0�B��#i��Z�V�L�~c(W+	O�}�*$�����R�Bl�S�Aꍿ���� ���a��Nj�@��}EÅ���k�f��)��,^�Z��s�J+x�L��>�)<slZ!!d"i������Ŧ7��&�Ч��ɼ c�����R�`/V6�T�E���8���=f�(2)�V�h����(ʵ"�A7�j9�j!bP�Cv� �wz�V�[��UT2��}���S%<�0�H���*Z��5X�$�N���5l�`r<h�y�W;GB�@��Lx��Hf�-[&��'�F0����	5!��j%!��"ÚV��3sU�D?�2��U]q�f��6<Y^[P�䒪4��P��⫪�r�zVr��3�j+b�#CIq�K�=|=��<|�[6�\3�g1 ��9"�L./�lGS�*	�8	<L�œ2|��0	@�D�J4L�l�0\Ĭ�a��K��*�*T���%a|]��p�YuUf�/�^�!��QD+�3�b3���C�HhJ�gE�"�l�y$Hj���g"�����!�˩߲e&Grzq�%$����sUs�����)s,�>�u&@Z�%�Ṿ&�vC��|�
��%:���RҤ��mz�e�r�- ◀%��`���7��dH_�m��f���u�\[�?l��%T��ēFN�����	��)�	��(�YQ�s��!UپM� I& R3rU�͛�?BE�"A���(�%p�hE㊓0Pׁs�(�E����+派�	�GUQ����!a��(b �+���W,�<��z���e�H0��B"��;0�*&�����V�UŜ&�L�H�H�" �r���ܶ��oI1�"�d�� �0)`l�*��i���#��P�J�<�4���H2L T ����HR-L���=s��c��	Y��h$���0#�i�j]̪�=0=<��l��;�8)-�Nd#fE�}��F����M�ӊ-rx�\�4y0�;<`�0�Ns�oa�Jq�x�����2�"�h��h��=��.-S5��! �/ ����F51�iP�X�'d�\�LH���[�d 2<�`��P��^q�C2�bMȣ"=~�9v�-=��	Ü����e���*�B<`z[Q�*FB����FP�jF@���bl�|�ZnO�uxa�Ex���3=�
 ���%C�p�(~�U�&%<d�"���P � >�
��&@~)i������sJ?3d.�R9٧�� �˷K`�"���S6s梼��7�`�1�ϑSJ@��䴮.�0�r��T�	 �����/	�s'0im	 �j&t�2aK#/9Y��@��ƺ*ym��^� ɾ�"������� ���/�0�Q�h*�J ������}[ ��k�024���&�����6V�OTѳ�'�$�;p�#0�Q�*��>��#��<�P4�<j���~�ѽͫ�??��ѷO����/��ί^�\��޼{��������G�'{+�W+���+v��,���ޏ?9�wcˆ�W[6
�z��?�x����K��._�_�4�����N̷5'H����<-?vj�(��G��fP+����++�bq��K�� �
&�:���1�ڨOt�DX�X�X�C�K+~op�Q���������nݜvv����LgN��{�/O�u�dz^/l=xx���x��]/M47N�����{���懗�{W�;��=�X���觻�����+�����it~}h7����޻cS��شAN�|�^zY���g﮿�s��G�|�/�ol�{o�Ys�d����ҶUo#\Z�䳻Nԝ��9w�wɎ�wo�ony�}zq�@�7��a�k7n���Tyt��î.�6�\_>���5�.�W�7M���1*�x�O\^]��:y�ﶍ��N����W6����1(��9:�z����LuxJ>�v��7�}���q<������S���8�꽸VS���gz��-L�e^(`�͛=������ˤvB���J^[������ok~G��\]�I�{w����8>3ju�a������_��ɗ�>�������s�V���-LҮ�Ǽw����j��{����������2��G����7E�X�,���NߛY���
e`�2��;�잮h�+�	���tU4xb ����i�6@�ML�ԃ��DM��X%��}܌{�V�ima>��eg���+W�Ņ^��įh	ֿk��7���8c����׀�����ư3`c]�����uE�kuUZ
-�(�h�S��(<�>M0��Q!��)tl�%�!�U`�i䢕g��VQBBS�0�3e�_m�	�4���5�H�����.K*^�}N%�R�ʊ������qW�۔����M_S�����}�=Xq�
#��Cm>�y͖@1�	���B2���B�$Jfep�b����G�Z��l�-,��\8�8�UN��?}������x����M�0�g�0�dӖ��W��%q�휥u�_�x�����/�ƺ�$���Xk��Z�����a�:�m!)0��s�ӏ?��9ce[��j��Gh,?6�C�ۜ����R�Kw@�V��|�b/�����@0���㝱$K��{h�!���K������|�.��N�qrԚ��=���E[O!xp�g?�ʟ�?)����1�U���/,�'�������_��Ӌ���5{Ec|�j\�0��i�� �F����L^/a#�7YU�m@��h��R4��G��/dzi�e�P*�u0p<�����3���-`�_T)ah�]��`����4¼0TK9���*� d I��iV�l1��g6GK�P�v�i1� )��*ʷ� ���c(U�����Q���M�SR۵�Dv�����Ǐ��RZg؂YRle�l��*$T�q�2k�wӾ��Bm���Q�9W�.���� �|�����bC�!�G.l��~n����9���O>�������h�M8枆0��h�/��OzHV:Ͽ��"a�V.1gB�3�5���@�H�����/��2���&k Y��2�b�L�j�@���o���U9N��Q騇�bE�*�0I0����f��z����N��!O�_؀�GRK)�
��>ӷ���ZVkz�'r����`4P�oq�Зݥ�t[z�h�P��T̗�Ͼ��R�r�H`ˤ�jT�b�+0(VE��Li\t��Ely�'�N��@�*�Fq-)���ڐ�J\�
���$�ya\ߊ!#+~[�PY)
C�M��/�E�w�l��i��֢��COHF���SVdE�������ssԲ�W���HM'� ~|�xs�����\S`s x��xQ�	����7���z/w��#~\	���''��Eь�!0�K�s{�q9��)�0����6�x$��i � �h���ER0`��MYQ�ߨ\����� �B��6�	54®�4M��@h���I�S<�Q�ϻ\�)�O�+FU؊<��g`�� �4&�"�$�rU&Xoc�d(�	�gLz&0�aYCz^��.�E`�kz��4�]-Br�s �*H���&������)�4���� ��� R�������`~U�qj)�G�gC>S��>g��U��F��"'����0�q�b+fH$R��F�S���IO�k�Q�DN#�CCVK?��� vT���T���8T��V�ɋ\jDL9}?�D?G�,��9LJr�K/09N0	�x�J`0d�0�1�a�4�l�@���CyV�>A]���ȪV�Rd�_2Mʹ�0�̤~����k��6jT�T�
~@��K�
�*��k � �^�a�C�c���9��MN9wY!a�-�U���G	����sh T1����V�Z)�a�j*�z<r0)eV�Ó	lU�Id`ak=�Z����U�umΦy�T�W��v1��@��6C^�qZu�y��3�bFN�	٢TJ�
~Uq��fՅD�XӦ��j0lVl���7�|��8�4��$<��J.<���"�4[�:P�9�"�KL T?��^.YH��r�#��?&���,���
I�*H&r� *�1��D)1�0УB�&�"a�Y<r r=$�3�"fUa���ߜ�yq�9* 9d�iT)6�\�[h>��s_C�,��;�x����������4�b�8�
�z��ғN���F>�Jɐ��(o�`��A�}m��W��h��U~x�R������z�6�W-<�L��� %�xjcTx����@O.����U�;�z�H�3��:B ��䊪����⡟�k)X&ţ@�PR[C�&f �d�Ζ_z�U2��󞋙G+HT|��*9�A$0�l���itbˣ\���=�H�̍#eN�UT�A��Ԋ�k?�Z���fqP��9��%/	0� b���BOC��ab�V0��#2��
fV�"<Lȣ�/C=fiœS�D�Jʻ��mZFU��0�U�����������W��?����]zL�;������n�z��7J+�µWם�:�&T[L��ǧg��׻�V,��'kN�l-��ŗKg'?|���ml{c���r��%<��U�$=?=9yy�Ɩ�����<��"����5�~��Q;^K����N�n%�=�ЖI���5Gy�����Lx�Nf���k�Oԙ����/������x%��ƀN'��C�I4�ih�jo��;���vꖹ���޻������m�\�����[�O�;~����o�#����ӫK�c����س�l�ܡW�Ҙ�P����.NNWn���;���_��S:z�oI�K<�x���g?>[��\�<Y�Z;�.B���cė��o޾嵬�	��������xk���]�P��y���8�c[ջW�m����WG�kWN��g�?}����S��@��֌��T�δ�\q���8��(��+����-��������Ӎ�u[��<���Uv���jI{����G9U��������[��69��5��;{�`��ݝMo�]�p�hC�_�^�.�U=9�\x���ų���嵛��lz�����Ӌ����W?�~����|���/����~]���_�pvzxr~��_�w�ju�ú������~g�>p����7�/)��3��!ݮo]DV]���R�،������@T�ǦC�7�grV�ϣ��w�x�Y�|V`f+`��z�I9�L��Zt�n��>|���L��X�f�d�E�/6�L?&���Ɣ��d�sju��R��3�\�	`
����cfL��֊��h7r=�6p(W%f��A��yB�.4<�p�5�w�|I��K4U�7�ق�![H2�8�J�$�9[9���>�����K���v0�ػ�X��]u*yԾ��+����"����b�*Ԋ��舐�ŭH����d��� MM�b�jyT��?LU�+K��^mI�������7����;'�n�ws՟�X%&�.��p�#�����㼻p�.3p��g×�.Ƈ�8��v�i�������;����5A�(0�'�e�:G��9'�8Q9^ k�_#��65�\�w~%Y7/Xy�n�Q���×?�p���zS�g���q�1�z�̱��9#	f��c��CS�c    IDAT�p�`��s���oJ/O��P�ŕ3���+K�w^<z��������noom�u�`��G���/o�(G�����co�D��H�9�"�0�$0� ز�ajژ'�Nv��0�7CE`2[�du�T�mx}�܍�	��:�(��a�KJE�0��E ��$`���.�j#�I�0��|�SUx ��H���6/q�@����g��: �\
�b�V	�O����c���"<�{P[J6>|��w��̳� ���H�垖Z�0�V�����䒘��4l��p��|'d��Z����WH�rþC�J�i �u�-*B��Ӗ�o�0�VsT!�9��裏�@Tb ��f�$[m�(�H���P��}�FX�"��|��L�Y�
��Ҋ���U��b��a�z�O��O�nX�y��d�B�
�pG`EoDp�%�t=0/|��0�,`}��x ���̵B$%&mN�?���2�c�XѬ�4�#�����i���#���G��@t;�n��]UM0�����8� ��7����i$.�(J���>BU���ș��d݈@Q �X`��#ԓd�i,=*9d�*Rb�c��1 ��T�C��IɜwNңUf(Uы�`g_fB'p\��f|.��`��>62�"x�xǠ�_�Ԫ�QT+	L-�D�5�y����V;Cw��w�]��˭�+�:A`���]n�	MU�-G�#�JW�Ky��R�L��P�LS�x�з0�B$���c )��3�x �/�����ԇx����ZJ�\UȔ��RZ$Ѡ*Y��	�&'�����L��o�@E<���0�%JllUɥ��ɼ��sÐ�4��ȅ�u.^���u] x0U冃�bz�p�ƹ�V���ܺ9� b�c0b@�ڑ�4�Z�8���/yg�\��h�j�EN�OB.�W.BE0G4�)DB��\�]�Qd�(E�y��Vl���!��ɣ|VV��'=6�4ra0�:��!u�0� (K�i(�Ud�s}�H��I/Q�.�&L��XmV�G���~��n��Ѥ�2�܈ę@z�\ �53 %2�� ���g��*+B���!�TU�@�$H"$�ז`r�*[�����4�0�BeN�<I�s�\.H�`P,)�*�i���K &�8i���ˋ_{�J ��3��3�V{90d����DU. k8}rm�T�Q���D��g��ժ(��$�}�g���"[�4�6�R��e.�~3߅��m�*�x
��5�/U���C[ř2!6�����zJ2[���P���Aޜ�8F B*��-ר�瓎@�s�k�f_�<&��ɐ����1�j/��\}NF)l�{�MŢũ��»���_8Κ�D�<v�^G����(H�sH���0s�B�5�PC��ҤT�&��2X�0��Z-ZA(2Q�/z<�u%A1%w E��,<s�jcH���/zT��I-X��Q�~��LR+�#Y�"< �j�Ϭji��a�y�#?_"p]��	<!/�&�y �wlL`�x��%�M�FC$�Ȕ��(T�-r9�$Zz9��"H4\�w5���H-��隢�-"�����b0�g���!~�ƜRQ�<y�F��4pA�7�7�Z] gK ���#0��R� ��!Δ��Hx�d�jk�ܓ��I�gB�Ȭ"$3�,a.)��Ա��(�d�A�X�ң���B0x��k&��9<�2=��J��(f&)�HSS��i&��Z>��[�u���L3�̖�J�/E�*��rʐ��0(�BH&e��� +�)����l�Ely�	�RQ�U5�|�e��k��VK J��G 搔dW��C/�����Q��? �L�}�%76��Ϊ,n���ٽyvr�|����=T^'{:N�.�/�o���^��o�s��:h����׮#9�����Y#E�(���-w{���a�q����7�`x���lW�D�8��8g���O�KT'�dd�ODF�^{����6�pxr�y�����d[z t\�O�Loj�D��{�ti�W�>�b�Sh�z��^�g�����Ь�f��'Ө���ʈ_�e:�$��M�T ���M{]�鿖��0�qr��xк�Fv��4�_�Ӎ���������4�X��c_����%��s�5��M�׬����>�����n<���޺�="d�{	/���m�����e���c6�g���c��B��^Y_�`�/_���O]���J����i�]3�n�|g�O�>���ɫ�������=�u���T�\_���鮳����DG����e���{���z6v���������ۿ��_����K��#p��/�-���]s_u��d�pa������^n���n&��_��D�v����./���]�ֱ���8RL���3Ol�AME��O=_w����p�cw�%�&��y���jk}ÓL��إǁ�����%�]Ͽ���Σݵ흃���/l/�����o��v�Cx������KOi]���1`g��'/|�?7z�����������בu��(��`Wؓ�ܘڴ-�mW;���p�))��Ӑ�]�d��4|Ƕ~s���O{
T&z�b�b(�8ɥ4��H $Z��X	�rk�zՀy5����bF��䛲�E	@OI����Գ�	�&/�Ҧ!�x&<�������Ӕ	!eC�a�Di��!J���eB1�BCR�@�R�����T&���7G�����y800��(����@�F75��W���8Mٰ9;�be�����/Ҧ!kd0���IOȷ�0H��lYi��al�B�h�^6�����8��/uo̞��s;�7k�����W)7
v>���+��k�?;][\����NΦ�������}K�����*�Qz��x�o��9~�Y��Վu:�[�������N�G�ec��XL������o<��˛�=:�����HS��a����f�����ǫh�� ��o��3��=]�s��/���h��A���8�h/�2��v�q}C��c)�M�I�΀O���х������5oQ�F�/�<~��_=����ۻ�g���"_K녃a�j[Q�D�D�)�X�L��mf�µI�� +�K�>�*@3o��@�SvH�Q2Qʓ̅��:��&�A:%VhrH�^�G2�~�dOf*�&��Q2i���%x�Зp�qr'h����<�ʅR=��#�t�K �2�!pz��L�����w/���_d��[VY�r+`��#�ux�Fc��rB)�E��`��'c���	0������_~��30G��������hvN|�Hp�ƽR�{��!w���MW�`0S��X<x �������3 �kxp�o�������ܝ9�O7�\�F��/7���{*\,�!Az�y��mu����J��R/A�$ ��W�$ 9S����;��,U$�8� /sie���W��k�S~���f�A)��	
e��r 4e �`��`��VP�����`��6��c��R������M2��R����`)�o�rPC/y�q77r�oSV+H&[��-�X�|��F�dH�-��	������#�!G�&(S�(Շ#RO�C��sg՛�"����E_�ܑOAF>s�0����rG��)8w-w�`䖒����	�˝�j�D�,�j��'e�L��5��K^zC��iH_��
F�{�	��ޤp��ަ�6%�4x1����M	�+g�S�s�a8�(c�%I=6��%���>=�!9+�@��"KO\T��դ�Kϑ̗`�#�\�2F���O�>憦 V�(ޫ�k3k/�1�慆�{<�nF��y�)�4�2	�_�L�Ǚ;��������4��#�iѹ������`d/0�)���a�[K����<�v|�`U�`ӏ�?mx�W����`ॆ�sr��G(�0��Ĥ*���X%�,h� 0!*�<$��B�B�@3�2<��MDJKV�v|s��MK��Y/Ca�\PY��pII?�.~z��29Vj�����Q��è��PU`f�de�������(0x	�)�T
z�\�����M	��ZeC��e�i� ��V�f1�r,b����L�=<Y2B�Zi��PY4�R��Xsă'�x�v��5J=%*mf6&HBq���a�O>���%���|��'Ք����� ��K�F�
V�i��c��"/�fZ��z��,��� � 2a"�}���VP��B�#$N�	g���,4_z�/=krs,+QX	z�|-���T�ܙ&��>""�F�q�L�!��>�bQʡp1�"9���}��P���'�L�b0M��������G�O���/��tX���R	��½LX۱0��X5&=`JTeR�h�P���8k`ɜ-���r�KO��2}9W(��+)Z��y1���E4$ hf|��B��T`��^	2WU��誉�8���"�U���#[�������a.��[Kf��\Y�q�Q��]Bk�nr�yz�4��� ���4;�d<R���Wo�a���y�qVs�* .�W�?��?�4T%� �J $��L�� �*������CJ�Db&p�6�(0!�sijV�j`�6�۷o�:���Q4��2'���P��B�St����!���D+�dæ�;�Z���#��F;���0~$�BH���p��/�^��Eo�W��L�Vk�3���bz��$!�VΦLgY����D�.�F/7�h5���5���YqN~cv0d�fF�`������$I�����(��0�9n0�zּ�3e�8!5V��$h�i`�S���j��E�Eϋ2<�����w����wF�����!=�5��E�LJ��<;���κY�9[V�CJ*0��4�(���ٟ�r��s�!=�׎����������a����O��������J���Z-�ܣZ[Yc肰K�nM����qUy��^ll�l\8_Y�t������;Υ�^��jO=:%��S�Ӆ *Q��\rs�G�r� ��݁^s䔕�rvdP�V\}���:s�7�>�Wm̔�#`�w�x8�磍*�Wbj�y�S�~���#z�;���)�����ދ�q���|�����g/���a�����ӽ�q��������^=��o��g�O��Nݖ�����V����mck\��Y�w�y<亴���yaus���;��~y���?������'��'���b�����Ǐ����[�q��S������[E]T8�?��}����W�}�۫ㅃK�֞��/^�|���~|c����k�=�ƭ��Wg\���v|E�����ֺ[���p{�����X�U_�8^JN(���vN6v�?{��P�ã��q�q0���$���w�շNn�`�yq�w�:ù������/|��o��D7Zq{���ݝWO���?{p��w/vΖO=�ꏅ߽��ū�vx^�z��Խ����;~{~�ny����w�p�y��҃���_{|���v>�覚���m��旛ņ�������X�7G~[��ݾ"���铑���ؐ��0�E!@t�/��$U�0��`K�0iee���+���E�� �4#i�D���"s���%�6��Q�5��r��(�Y)�K/sJ�\t�@OCO�'�EI� �i
��z#�8vM1{;2&w��E/" NV=_C��Z�9�*��\H8��P�(�G�Gx�x��+�Π>����QW�������H[HiqƋN6(Pk���kL4y���WD ��X�6+�C&S&c�n�1��hQyǜ���"��C��_�*��������������+�֯^p#r���dc<��Qxw�V��������o��~�E��9���7ee��*=��q�g W��b�RY�^����E̱��F�By����Ǔ���p�����5�/.��a��9���9*9���iL��c�/�չ��:�QgJ�F݁�c��{�b��;wp#ӱh�{�s��[,���sW4�=Zp���������=z��r�|i�7�x^��x友�k�vzu��՜2|�*�<�壷�d=���5�w�d�	M����@k�U(	ZV¶����%=̔zmb��h`�d�G%�����l�e���h#	f�f:������c<��$�4z �8�E	�Ō��f	#" �a畆����0�P�@��J�l�}�ݿdu^�J�4����gy�r$����^���$�{!.t�:��޽{N5��W�	�)&%�S.�(9�&�a��
�攎U&p&'�SR�g��_�m��Ľ��9b����02Z+�A���acu#S�mi�aΝ]��!篾��AU>\܉q��&��$����x{kjL�L�++M�u��ӥ8MD�N�%o:d��𫏄�	�t+TJ�|��X��Y &	����n;�|�MVΐ� �Eq%�Ƽ0��*&_^��B�&��P�5�B6p	(��#K�4���ǪgFvK��!���a�ע��X���yZ))ٙ5W]-���Mk8�����J�
ȶ���L�bi0�����#�A�*O)(=N�\���4��i�	J
�Rr�TD;S��� �Z�,���x0�3BS�)���E���d�)�"�-��2�&A���2�?�^�L��7��P���99�^��4��CO��f�D� Ѷ3�B5�v����4�D�G�d��ϋޤ8R���7L/ki����0 ��X�
Qz�4a�h��`$��L4��U�@6Yx�^hY)M-�y.qr�O0��s�k˝F�% V��&B0$��u��:�J8)�6�,�P�y.��iW���ؐU.�d�j�i��C�&%�y�����IQ�y�HbN�%X������4lx`�'�kd�d�J�Kɐ�ЁHtS����)I C;M���G���0Qj�m�4ج��Z 2�4�=%NTdV�I�K���,�ͅFV��4C�L��8�l����3��c��:�ȑ�F�E�V��)�?���k
8: �o�MJ�L9�-�pjK,DCz����	q��&�LzY��$���!Zx}9���4i��
&M&)[q�	5�/��%o(
*0��L��'�!w��-1��7.R*�r�ck�/*�!K8�F�ߡ���;�����䶺���$o�E�$YK�S���I��4 � ��Pq�:��l� W%�"rD�/O&rT���4S%��U�F3#HCqŊ[��@b�7,.�9��V�a�!e }u���*A>��IA������
SV:C��FC��2�Ť5���"N��04�3 3J������m������/�s��GVzMsa�)�L�����z�`S&��K^0ߒ��5C�^��)�td6/ɨG2�ܐ����m�si}z����ʡzb0A�f!.G=$L�V��(�ނm]� b�j
0��K�&
0��� A���l��%CO���LB��Q��BK��4S���Z%��],0J2/J$
K�l��B�?/CH����V�$a�y]d�K� �Ґ�	Q+y z��B���(��E&��ʙ;��s��H$ i��q�%T4����P����yy���\b��ͨY��M��{(�>�QҰ
����5J�Pj1Z�4zɋ.�f�+S)�)/s�X ��7Ǣ0�CN���	RB�'S�i���z���1���=��&g�[�`z&'`���_ʄ����XD��JS���ڬ'GnE
ZVq2�j�9ƙ/|�0���ʍ���yI	�>�i���$$A3����e�WV�^�b
��`�v���{���nj�S�JJ�a6�C�'A�/+}9�/"/�r��=��N?�03gx��2_��B�u�w��Y���W���_c3��&7�HL�9��㝵��å�ݗ�|i�͇S��U���<;
�?���8���#��\}u�nuw��ӗ����w����}�ײ^���˽�>|<~�I�yj��`.5���fh:�2B����W7�/1J��<k$�|ưO� �L�= �C\����F)��8Vq��x��qN2�^��kA��܅g/���?}�������?x���';?��#	��w~��������7�&�K޽�œ�����U9���(��kׯ{t����.p}��g���s�+��~��G��w�>z�����ϟ=}��ӓ���'����tq�ҹ�|���W�-�z�1�WN�h<;9���_l_�ܵ�    IDATygese�d��o~s�7��7}���?������on_�<9�s��Mj_37x|�����+��k�G=�v���Kk�^�v���>�|��-?;�T÷:*��ڪ��y_���|��W��}bџ|��`��i��u�֖�o~p����ųu&mm�¶�+[7/_Z�G�[W7/�׶6}�����;}��(G����7w�}u�d�p׊�������/}��oV7VO��v�	o��ǫRM�o�?rr~����|�����_�,�-\���@��i��f�.��g?�Y�flk
`�	V��!�=c�j0���%�v�xeMVK?cf<�͠G wMQ�ȁ>�I.�9J`Tz�h�8�[��0*C�Ƥ�ېi�-Z��͛��������Z�6|�K�9�T����=ܙ&��5� &���d02������:���[e�Q_���\?�	��U�r��7�I V����#�u�Ji/1Ѹ����: ��kq+���5tSbk�ĕ���O`n��W^\�)��%	C�j�-K�&<����S�12eu!+��W�q��V�qҡП.8	�q����ࣧ.��������]�v���ַ�V���v��[�x���x�\�=�q�p��t�p�����8�u�$ڗ�N��8���ќ�>���Z؍�R�qrڔ�t(�>nm�Ḿ��0��݋ӑ�vZv*�۷OV|I���0�TX�ӭ(�~�x\���[���g=v9bz��-Y7A�c�B��X��Up�O�3lӏ�;�.�,������p=�~�j���;_~�Ͽ~�b������u�����'��F�M�z�Xʖ�]K=�~n�1p�"d
6
2��E�f��OHE�4l���R�|y��V�i�uf�����D4�Ӵ�	�"����kðڣL��0��C� h�so�dV���5��{B�P��#6����a�� ����	2���1Gȗ�{%N<�4��Ml�ud�Ag:��$��i Ew�C��cgKw��u����;[}nt�" <@ÿ(�S�v]�G%+qݬ��$iD��Tn`L�@rQ� SpRl����aMzLb���e%C�q��ԺU	P���KCA������b9������!~����.��>&��x������O~���p�,fm�0_|�w��("����5CM��A�8we�{��{
+n�mA!EG���< +�������☚��W.h-A� �``%�s�:���ɭ�p��5�d۝;w�h���p4��L�4��:��)�5M.je�bi��&I����B75�˾�����'k�;�)�ׯD�u���]M,���Vna c�
gVg��	F�5m`9��k⦬���#��c�gƀ�fHߢ;��dLr:�`V�����#�M·F3�;}~�2�*;�L��	f@�|)5�*>Bʢ�e�'X������_��#$4����	 �(N �/A	 �SU�N�Q&ziԐ��<���c�O���4�u�A��	�Bh�Y���**}^��4�/.X�%�=S�������/Ƕr͑�1������8!�P\B�����ΕO/�f��!�2Lc�p��ck�k�C_z����F>�zM8.�"�!0_B��D��zH&u ȁLPR���ł�=��Y縊�}��12N�Ò�H��,~�=f}�ث�&N%w$)��Ā�)$@�`d�h����\�Lm�J�#�0�*�)a4��	�6'w$"M&�ϝ��f�v~&}���u���B���?������30��0��"s4�$Fi�轝I���Q�NVxrC���!��Bh.�-t��X�c=0}��i��%��@b�dH�Ԋ�{�Ҧ1D��E>��XU� ���6+Y��L�*V����$�bM��&�֤*:A�0�	}B�0��D�g%��0�%1&��BoW0���U�VK��p�N�k:��)�3�f4H�yf_`2=��PD$zͰ��)[/��2�T@�x$I��	�zY�vT�?60�B&	�� ����z�D�i����	��3��
���?�qb�t����d�m��7��hJL,�*��%�^+z�l�̤�ԤDF���@)m��K;6�^�ʐ#y���2i��hJ]zx��S3���s'��K
	 �>_T�̧I�YP��25J�x̢��D�ǜ�U,���1�#���/��aU�$�W@����1=�T1h*`H(a;PA��ȳT�;�e�IXC[��a�-3�]���@ }鱖��"4�d0���#q�H����`X��`%i�S�@�fj(�4��6JQ��55�,�1L�G5�2}�����4� ]�	+�p����;�>6�"��P3,
�<�bojN���j\��,1���`��@�J#�i�xh������|9���&eK����#,[^�d&=+6Q��kYi� |K�೏�v�h��X�y� �k�jH��VDl40e�\��Φy�o[1Ћp�`Z�Ʌ���@a�c>��-G^�qa�$T��5�D9�=Sl�2ZV��T ��,����H�/s=@�4eH�fye�$��5�Q���/��FV�!����Y�A�p�޽����w}�o��oli��dN	i�;@"U�6 YJrp�<?u�f��JCrО�*=��@jJ�pB{a�����57��/��.?���j8j��Ħ'�������LlN�*{Ud��#�S\�Jm�YP;�G<�U�#��*��~�ӫ	N �w��YAX!�w��K��ׁ��sk7�K�J�9������ח��|����������q��������󄽗/������=9�����֕C?{��Z�'ZW�w�#
�VV�^+xzt���ܠ3#3��������{��=}ⱥk7߿��5����jUO^�YW6?�G��w���s�ߓ��������g?�������`�|����?���we����.���7���|w�|�la��|wg���y����v��8�r�w�.�RY¿ua�ol��z�w���<�;p_����Ζח}�������k�'����>�ri��O޿|�oR�9�w�aq������_�|�����͍K�/m�����K����������]y���^�X�r}s���#��.����f�t���)'O�z�:@�
���m��9�ۛ�=9�;y���m?����?y�ضv#�?(�-��?�����߭��K��c����c��	�V��K�~#��!g�妩�EHV&$J�������:�X�7�LbQ�I����Po��b.�0�Q�2G��t �c�8�T��`B6B�$K#M&�#' �	dPn���L�9��K�i��r�P #A��А��jɎB1�3��w r�b5)��z���0�x����6=_��\�Α^�	���4ՙø�o:óѥ%��Z-$��\�WBzD	i���b��K0a��=���(��!	xd�W |i�`��}��Px���My�4���`����󓣝gO/�x~���O�_8X;�Z_pws�m���/8�yQ���AZ~Yyt��2y���L#9?�;}%��i�e�'㧃����-.��C�ȹ��i,�����q�����ՎwȕU�HW����1,�8o�=a꧆ǳ���ހ�!�u��c�c+�i�p�9���j{��B�1Tn�e���ϮK�7������W������6/��$�Y=��&�7&���pLzJ������in#���
9-�X,�V�	��%De؂�8��a��h�z�mKVx���z
�;M&x9�ZogȪ���f.��(	E��		Shi�[��dғ!�aȨ��!��1�L(D����r��d�� ��0ߘ3!!�zͷI���p�����U�m��o�uW�F֛7o4�p�}�]�v����JbF"a�|ntG�w�L��r��iYw#�����eV��t�!Az>��Ρ�),���%�ȁΙY��L���j�2;yJ�#6�q�	�o���P���@u�q�~7�|���/)Iw+Ұ�Rx�F�\�a�HT�2A��E�-/�LM>0�'7g䦠JL&.����e� fR������Մ������	ҋ���M�ڔ���'�����$_��C�-^|�j���/m� 8{��5"���T� �y	��כ��m-���5�o)�I�+PY��`��ˁ�j�YEi��Q�M���V�4\42e%Ekh�*�\`�WB
'QP�빋��T��)D��i�z2���p�c��[S�6Gi��^�ͅcz0Q�EŸ�M>s��$&=M�M�6��9X��G������= GK܂♓d5}H A�ï���Y�YDJ=)��D.8��4�4yA�p10���ژ�m�eNr$�+Ί@ɪa����0 ��[Y�Q-z��F�K#���i>��R72L[�# f����� V�����J�����%G$dي�9����TJ	!�0S��E��T`A)[}Y�kv�M�a���@��쀓�d��
M�9�p���B��|�
�^tx`�Ȭao3DU�b��(�
�{U*[T9 �Zz��0�	�P�h��c�����W�M�|j���	0�ȅ#hY-�!fl� k���h�͂�,��SL��.C^^G���N���P���sة ���ͥ@oW����^�@I(�4h�$_u3��`���F#Ôj��ߒ4L���� ����������9�X�1	)s!��M�p��fD���aS������\�
aػ�yEKP�6r���@b�� ��bf"���&b�`8y����ՑD�R0�����2��Œ� ��cl9��Sr��/
�T��)�ް�qRb��gpH �><3<�|yQ���L[<�U�e%7�v&�KQ��_=�VQ	���Ds�M*_ x^������b� =e�z2eVC�Z��T{�& /C�7��^yR25G�
��-=���u��:2�T�^P�{����ɥ��*�o+wx�rVP&.�>���4V�hL� _C� T���r��@�1p���`�yu i�&��^�iRr���%���	��ge�`���C�~T�<R	%�ƅ�sl� �\ʖ�ư�2$Ǔ��V����غ�,y����H4.����l m�������@`��f�r	�9�޼�ܑC·�H&z�!�
IO	 4�!�?���Y���G�U�����|%,(�l��I���(�ra"�@*�����f�E�.���0!�|�kR�D�] yJL�T� Ҙ�Egœ2M�JŖuf&x� ��}�U�G-�5��E�����$��5`���C��W��l�X�'�H�],`�Fk���74ق΁�H÷�\ ���wֹUp� z�6���|i|����1�i?w��k��bᑏu)�rF�DFc#�|i������^�:J+�5�]oH	��5�&�K�/��/q������J�j�}�'xM�u1�m�faa'Z�P���Y��{�����ӕ�s��n�R@���t�x�O���$C?v����ܵjq��h����)��<�MO)�����q@�ѹ�'"��h.dI�#��i�)Uޟ%k*��`�C�l��lmm*�?~0;���?���a��uw]��X[�|���7���%�����ÑۥKW��sD�ۛG��_�����tf�B^eK^��6��,3e�w�|����#l/��_e2Y����ŏn��ݻ������Ӌ�kϟ={��Vַvƭ����珟���z�st������gm]�䋏����_���oܻ�`{qu���{���_���}x������O�C��O:9𝎻O�\��>�������ʥ�>X�yk��l��wO�.\���Ջ��~�u}m\9���~��򻟽���/o�����o?y�����'��׮n���/������e�����ލ�7޽���y�{u�_��p4][w'ǚLupScy�ʅ��~�흯�߽�����~td�w���pt��n76���Sc{�i���un�S����<�}uk�Own�M�}��/������r5�u<�Z{Yo��kY��.��K�d�v�&�J�f4�=kg�$�rRb���J���M�EEH9��K X.zl04�i3�XYgMT�H0s!�3R����C��2A3�T�^���G3'���s�x4���BS�ՇM9��'7n���Nz� �g/.��ԗ ��/*����)�Lb�G�Gn��&S��EB�����5e�9"���|mK�n[N��AɁ}ܳ$1�;4
�Ld�]# XȄ�ҋ�Q61	��ח4[ʼ�j�At $Y��BJ\����{4 r�CFb�U�����������?�{���}����/]{����;�<�7�+���#�K�g0�S�~��ߞxѻ�hk���V2�iM%F-7-��7���6��B���ڏ\=59���;�BL��1VNϙ.�_���#��2)��G�s�2�7�z ��I�~�Yqc���c��N�J���*ָ�9e%��lz��kw<�N������ٱ3����>޽s�ɣ�g_=;9޸��\�W]��w���O�|W��o<���N�����,4l�&��\�LEh�ch�+%w^��1�iG�m	`	ș��� �VDXA	�1���:�qzi4��9��h˼�?#)����ᛵ32,s�(�ٜ	�3An�J�#�Z��Ύ��e65��b����\y2�M9�`�� � ӼK��a�K���g ��	� �C�f!�#����]��[����z��_��_�����;wL�P�%L���_�E�+�w��?�̙́*.�3�����۶���}����I�����E���C�tʫO2x����Pd<����t���+��4/ٚ)AqP������o��l�ƍ���q����:��uA�N�?���M�4ռY��o~�̬�Y��<�˧�~�"�'Aqbk�T+r�0M��M1w9���|0�2r����f�f�~*Y�8�p~��'�%J���B0g-V�	F}�:�X-P��^P	LV,g<�B��/�b�������� O{@�d0�""4ql�d���T�2UiȜ�޽{�1�R^`u���;/����
��jH��`86$0!�9�p8��'�)(����o`�VV|�,%HQ4z�&P�*`��EL��ID}�`&�ɔ�آ/�W3�)(YCB�0�d�&LɎ7)&=<~�\3)C0�z�4�P	��\,^Qѳr�RF�q���ȑ�c;�>AKI.d��d }$��`A�ĕyx.�\�d�[�i��aixEUC���V$��DY��Pbz�c�OɅP�eE�a޼wb�r�VU�Gh;9hT�`*�D�&V��T%�r�k"F+(�՗�=a�4�R��dG)5�3�	`&)�B瞆�F��'�L.���s����)V)�a��m��1k��\Ce�+e�(���x�C��%�׼�y�ZJɐ�C��dɚ��*���J@�"�CI���(��"ӳ4��s2���"(E��g�a�f�!}l�x���K_���s�,��fF��Kk. ���L���N���kd=/=Zq��L(��
ʋ�4)��ǯ�c1�r^zz<
AY��
Ҕ��·�r��=6CJ���#6CV`@�b�����F>�tp&�Q!� ���lY�)_T�E�c)H {�����AK�	T�4T���c.+"��(�\����; /&�9�m�����ˁ����ɝ��I>��]&f�h4V�0�jR #�T�f��m@I��v�h����P���Ѐ1a��� �ӤWyV)��iA���z�,*��%�	� �#��ud�E�F�Z�YU�PC%gG�dC�8)i����/+�$���o+b���/|T�H�Ro.�Ȣ������͑I�&E�K#tÒ�Ĕy	�� 	�DB�ge�ǩ�7)~�У�{.�p5���#�{��P"j�KI\��	_ '�4hE��&:%�#9�����2᥉��lF(�M��1��,����9e9�Lo�!#̽�8V��� 
D��9�ܙ8b֊�,�͂�pf�B_>bq�S���`�X�YC/��B#���?%Z������� ��p�`��#3猣    IDATk'�a�5q	�&��L��\ 2f2S�ĠQBJ@���H4V2Z2L��%���'�dV�(a�b�[` Q`�Ɇ 4�4h��ሙF>L9�ӓ�th�	�P��+���+x(EA˱9�"\HV�"Dӌ8�Kɤ�$ Qd0 V%�i��a`"��u`�X��S8�L��
�3e�"��1S"1/=_`�(z�P}��c��5�9� n�y���af-g�����
yi�����J\H�zV����DFɷj�����5[z4�d�\0���h^B������k�kj�]BqX��U�#�)��V@v~�k'��ZJpvl@�F�2�����Ð|ݘ���z���+��<�ny6�pU fx�
%ˍI�}j��:[��Έ>�kT&��TU��q�0J��iФ�7/m�\\p*o���.����������z^��ܤ�9T����zg;��:�}��r��̃�G���{:pJjIڮм|�{x<���V�o�eP~��?s�Y����Wu���VB��q��c;������ŏW��w��������O�����h/^�#�9��O����~������?��o]�r�k�|��7�޻�W_~u����y��R/Oݩ=�ta�3�ϟ����O_�?�P�L.^]]�\���Ǘ.l.\�����u��k�]��V7���������GE=`�^������G�v�=��$fuek���{7<x�vami��η�����}�r���_YY������ڹn���Gg���Br����с_)���x����v�ǿ��he���p���=�u���޸Vv����v(?��J����[�>���O��/�I�I��y����*f?؄���.�B���0-���=(�+bH��ZO�4d�4ˬ���b �x(gw@������2/$�T����H�T� �p���$������#S�!`�GH�C�ny1����hl`"2)5���z Br^4bqi�LB���p�����zCq	�c�g%ȟ�,<0� �JH�C�/��=S��2��/�ӫ�9*�f�M�я,��߱S��k��w��}"������#Q�!�C�C-�1
o�b�
�d^#�����YNo�0. A��b��3!0B0z2X.�8�����ʰ��e5�l&���O�jO��c���2�z����﮼��;7n\{��������8��g�[������zj�榇����X�^TB���0..��o������i�ű�=I9Uc�ڡ��eE֛���%���>]_;~jأ��4����eO�xσ�y��tul��<�I�6��ǉ��0�SE>����:���-H�|Nm���q�g|��������ONv� �����Ս�1v}���c��M�_�\��b��N�H��p��͊Oy��u��v����jX�6�F�����GË� @o�!i4BY���Rj`�L`|����5��L�@S B=@�;+yb��4��7%�@s�ds�,(؜0���¡�ї�<�c�g�Uʢ�-@�`8)�K�LcGx�dB�)�H���~*:��.#'%x�8�8������#xJ7���9�0!t����&�=��`:���c�G}�aΦu ��կ�P�h����i���:����M���_}���KL=�P�ǎ�u#�	G32���1k��{��]����:�������+*VGX����a��d�`x��冥f�nCv�JAd�8\z U�|5��+�Y߼y�9���O�Gh�T�X��a��3�U(���TLH�nH[�?��?�c
��`:��V� �����bP:kg�[A̪g���`4��#Pb����PJ�d^�M ��#�!���&�����'�۷o[qeo�aP��N戇0����-j��:������C*=A#�k��&�ސ��\�j�(���#�am!��9:Xl�PC;�֭[^� ,^H��bU(����D`Ў*./G/�)� iA*>�fZ 0f�@6;==��j�B�3I��P/(/�W=��E�ԊLhv�fđ�܅��	@ϗ,��*{r3Ԋl�H�;/A��
^\.z.��`���'赐\4. ��		Z���p����͛x<�hK	̶�Z��z.|�G��sT��R��Đ ���T�h��"��}�����c�^2C����d��\9�2{�X,�`�6YVz=6$�9J���g���a��a�b�_&� W��Y1P&��C��6`�`�&
X=$�9�r(\J=%r���+���[G0�Z� ��q����8BCV2%���R�i �m��\(ˁ>/�4 |grqi��疉�V&z�B�&����c9 $�hL�4,Ù� 	`�L�ʑ&�Ls��0��f���#�\�Å�3��`QtC<z��(�`���\�j�ʍ{�&��'�E�)L���$ H�^&R�`���_ּ����h�rP7�dQ"��9�?�E���Ӫ�@Rj*F�! k0I�JO�L�!*.�WvI4J0$zlz�V�2�į9�C��$g2<zJC��¼M���%V����%pH䔐��� ����pZ5)���	C$3��$��)	x"�
!x�]D.	�@����bc%{�I�]_P}�z$%L��sQg�4m�.�r�Ʌ����LZ�cK��-�F�N�I�d�0%MShwqi#���@6d�Y�D'�c�*��4����4�h�J�#(�����R?�R�%w`��hpjR���4�h��B0TL=k��H��U���p `�K�or��������ңm�1� ���4eC0eq0�|�7G֨ ��-e������c&H�\�͔F�%�5Z�"[JH�}i�b���Y����0��R��oȑ�R�Lý��cҀ�gN�m}���k��|�1H,��^�x���Ug���B�Bʄ��2����!7;���k�k�*`�f����,��}0�Q��!�X��K ����50��5fr` Q	�f`x�9D� s<�)	y1Őc֘18��XM*ِ�9Bb��_/C&�����Y��3��H�S�Ϟ��|�V�\��\���b��AXY�� ���_)�.���ټ��f0���jS�4|a�h}��M�b���\'sq�֭[�+u]�] [\��i��c��*8�P�C� 0�(���{}.d/�����f��%�jx�Q��X��L'(@#�y
��߯�`ZD��9�C��	�zz�	P�s/1��՗ *&���V4���-дg�=���������]�f��2=|�������tz�߷.n����o9���&D�WV�b��jǾ���3����7+"y	��s����/�1I�N���!E����8��ث6�G}x�ι�<}���˥����?~�up��'_��Ó��g�v��}�t��`g�h���'_|���w������W_y�ᣧ�=z�<v_>�ɱ/nrksճC��C_�8.������ŗ�/��n�oyO��~p{��r�����׮�����O1�[3wuݜ8�?|����G��o����#|�;��v�o?��׷�޾kӮ._99xxq�G'~�sc�ʶ�NX9><?:���/Ɨ0��?���=���3��=�:��|��knݬ�e}��Փ�y����e�i��ݪXX>�d������<:=:�]�,�����Ts����`��\�]k��L��FoQڍmۏ�\?��pb&kv߆&����W�P3�{^Ƀn��G�C�JIF���f^h�4&^V`A�h^�R��0;f2l.&H3߼bh�9Z����&�ٝ�LX�TC��|5&.��h�NfX$L�o���G�i�,e�3'S�dTL͝ Č�<09�r�'́�C=�w�"��VJ�i�ާl��ܹ��T�?�]�tD���i
���N���hU���ܚ�^~����P���9�F�Ӊk�ʡ��X�l��3Y����"�����+m���E3�Z<?�s�9�;t �]������ō��퍥��G�{�vX8]u��ڎ���˔����mL�9�t`�hc"�k�7,��l�3�ed=nwNɛ�G-��ڷ�K�!��Z)R2�<l�q���Ӫ���ZO�����W�v�o�V���&2�7�=�7�V�M8���ɉ���㩿���ӗ�b��#��^<z��W��}�x���������USp�Û˱[��==�z~<�Z�4�K{�Z;eWp�*�>n)�kY��X�i��5R}s�Ж`��ѣ�0PZk�I�G�'H�D����
���߮�!f{# A8��T��`
���f��(�&s�$�E�5����<��#ʟL�G2�JA�s�Q��)B���A�Xs/DQ���� �i�i��],J�><YYȕB���|����7�H��%NH$�w�m��nb99k�錙Չ��۷����������?li�p�5� ���>�N�9P�̜u�H/�ܪ�;�N�0x���]g�����4+�,�{�r0q���L�t*lj��:��޹s��% Кra5����Q1.r6�N�i�z�M=st)�JO&�龃�Ў�H�[H����y!1�*�&�n��("���Rg�_|�~wy!��R����ɟ��В*��2/���H�`jV�!i�4ؐ��8%�2x0X9�P ���Q�,��6�)��<)����x �����J��N� �,di�&��8���"��L\4��� HpR�T^ӤA(O����U#KI���Pj��Đ`v����Wީ5�;@���
!�&�=A����GP^V^,q�4�\4�)�K��̥�`X9��cg��2��7Mz�K��:�<��Zt)7�$ɋ{=0wz� ��fA(IV���a�/*zÔ�}�*~A�'�gr� ���Bh(�P���)Q$0OA���1kɔ�r��!_V��7}[���i�ę��!�b���4q���d<�(��e��&����\t�	���D � p��諏�S��yii�]���)�aȔx��7+/C���!�!1�U2�^c�J�x8J8<�R����'�K������fb}��dVz%����s���N���"3�hMA�Ы�L�`�9��#��1r�4$T%��Z	�����
����.39.h焅NI`����޴�s�F��R_)x�� (ez��s�ߐ��<�"_zJ�9V�����<MPjx�gʚ�~�	���4��Ͻa��e�!}MPB3j�� `����;}&Ѹ������V��b���iK[�4�	a�k�]U�X?'�3��� а�K���(���w��%��ܰ�0�| �Ӌ�F�d��/.�<A.�&g鑫����kG�4ťϑ@�
�(d�UI"��3����b�>3C��i��L��f	��[nr�4Lz��F���[C��c�S�T�Ц�aM��a�_�)�|,����Z��>��X)��
#CrCz�XL��9�f���ޠ/Mr!�;}�r��A�*��� ��dM���MLK�'wH�0eE��Q�v8kH�s0T49�5.zl&�/*� ���O� )V�R��^of zld0z��)�!52|�1�tb. J U�Il���OtN ��ʙ���ʑRyi� �@`%�d����az���RE�a>��1TC�ƫ4�yU�D�A>���F�� ��X�+�0z��'�pd9�0Y�aޞ)M�QV��(��87C&��L��	X� Zl�2!�K����� >�� �h��P�k���dˤ�4^
O������qR��(H�8��#қ�3R�%��BT�H^d&`�dJ��M�����>���(��G�5*r9p1�h��C1���C����~8]j���L��&P�@}�U"�h!�!Y�{�i�ǚ�qVH�>��S�������dV+(:	X)�hՄL���j�
 ��)�}%��4w��u1D^~��pr4�����6��r$ �8�5�|��dF#s0����o��x�q��)o^�eXh}�L�^�뺓�(�IY �J�����}0���hцO_/����a��UFP�Y8+��%�u��"��&1��D��|����_b�҇)�N�Kŗ��4 ���Ә��z�������b�a\�he��y��v׵k�|��-�.�����7/��}2w�W���~����=�~woǬ?��C���xd>z��������^�������66_��7�V�Vl�CW���w^����6��?�s����g.�΍������񓟾*vmi٣���<���_=}������١�=�۞Ӭ_�z�Q_�����ۿ���Ư����7/nl�z��ԗOω�gk����+:O�P��񾇟�1~on����q#��l�4���#�s����
�i�'���<�����?���o��}4�R&߱��A����>�X�;ppM�L���!=�X�7�	i�ɒR��H��50�Li��!�a$�m6�|�ccM�8J`0��ɱ����9ʇ����S��P�"���9���L�<<!�lbe�G�9A�^���f�A6e��(z-/<aʍ�Ɗ'eiGH���`�|iȐ�bS��,<f$8��G32������^�^�%C��r.8�˼�B{Qw���7�XG'V�o�ua�+"�D$�c���
F(� ܘbp�K32}s�E�eP��%�|���`fҋΤq\L3a<��r1���Fy	�'��Uw"ݕ���������������w�y���K[��V�W7����6��ڳ���x��c���x�y�N���c�K�g(MB�{P�Dݘw�&��"s�\�1���,������ҁԯyz;R)SXvs�ėĎ/�]<wOԊ�#�� �G���Ϋ'�ώƖw4����{7��Uy����}��_���xq��e���}�qD������p�hZ+^ai�G2��&4Ta���. f�gKnQ�#�Ƌ�!��\���dxz��c�h)i�`Hbc�`�L\L����D�B���zQ�E��Z�!�ټ�GPJ.i�i �S����g���ʤGN�7ĉY#�)���!�֙"�9(�)�#�s7l"�HdB:0�&�^cB�-�!�ˇ�l�8�8S�;�����������NAܣr�p��}ln���P�0�ߠ"s���0;u�3l�L �v�RZ�+�*"Ǧc�ԝ?w���Hrl��s�>��V}��I�	���{~�˙�c+*V�N�|p�!ZG[��`�kj����W��d�U�i�Υ*ɶ,o76�%ls�\�C��pI�#:"���ؖlK���K�ê�~�|K��΀��_~�9�\s�5��*`x�UR��S�����kD����~��Vz�*�k��?����dt�^���XR�KJح	�>鉺{���0
P!.���E��MU��şj������G±y l���ʶ���ҙ�e��1�n� PiP�t������Q��}.�ҩ��oxHF5��h��-/�֐�Ma��ڜ��F��Q,¨�8y)�x����KQ /]_��%d��St�k�Mel�+���#CȈ�"6 E
c;E���%jEQj�Ċ�֨N
#Le�U%��\\�G�V [�e��
3�ف1S��U�f$*a�-E� ;b�w�0x�+ܱ� u/$��R�7�^�bu�R�0t�ڗ��L�P�'�� vG�3#d�4��H*?<����J�nj�`���g����q��@v)�m��Y$�H�lreKg�4�Q�̛R��1����H��Z���3��/\T@Fz%��R/3m%�j�m��`��g�9@.S�Q3W��!]"���3E`F^e�CF�/;#�`�i%ͼ��d+Q0x�h�NA�� �B�jt�Pl��њ��	�X�IM��sA����h����T��,A�QB�C!5b
Y:��g����H*�b�rz�9��/����*�-Qv�r卐ΫH��ybjs���Q,�N%� P^��H��10ւ�2��]j��,ye�v�D�Zc�M!g1sb�!���u���T#)AH7���32�!�6�c�6a٫GGtF��XgT����D�e4��0Ό�aر%��1S���XT^Huҍ\l�_�)�@��7@l��Q�D��B�[� ��d��.�xtF �G��RT��F���B��-$�bS��P�&�Av"j    IDAT)�b�\֫'�L�b����bM+�[��kL�z�a+����S7�V%]T{@VI�ٚ)*.�]F�7�	`����ʹ(����j��eaY/�x���Ĕ]` %ZƘ�h�#�;��N��j	�E#x�b�� h�Ũ��S���\/�+��Y����,�Ƥ������IT�[S��C�vc�/!�첈����H��P3] ;@����Ea�����T����W /pxzY`Xp��RO^Q� F)�&�Y"��^�#�61�fԅ��l���1�%�\F0##��tJ�Ě����JI��z�-��,�%��MIu(�8���e�� �_�/ƪ����+E��W9<;o�������ő,��E�b�Ű+l:���������n��^� t��(#~��K/F:�lʹ�`Lt�K���>1:��4�(v�3�g�.�U� �@R��l���d�xY(M-��aA+<����N���L-�:�.�K>�w$3>x��G]F��X��)�I��a����v0��������]�u�0:c�(Q`ȉ)@zJ��������g�NQ�Q,E������ъ%؄FNa��f䵤�ĺ�����  ٍ�?X��Y���Rv<m������]�A����Ԏ��v�(�'��cl�U�#~vz�
��ۋ�7UXFv��u���$w��'fz��-G�����)�_�:R-*ˢ�j�����H��h}r�·����K~ZV�������}h�~��7z���k��m6~&q�0�Q��:���k������L;n���;�o�����?�������?����=;>��{}/��ï�>�������|��||���_��P�S��㮖ggkG�O|W�C	߀�۴�8·~��Rx�q�4��9��Ď���т��������֎�j��O�:9���8;�tm�ճP�<�f����?q��#AyKIc�C�����xJ���H��o�����GXT�t !�г�d�E�Y���M,�}t�PL�1�R�4��?���g�f$46�dF�a�	�ds���>��=ɵD�u��E*���/���fr���kn�B�}~����8��y����9�s�[,鍐:y����~|���Lڿ�V$�W�������4�+�TuiP+0d�^�U3e��$��'�o^�VLO����GWc�YI��s$['��[k�8�N!�P]e�\7���/��:Z�h���!i�N>�E8X����/d\b�6��G�%�&M%a��1����5č7ćm�S��,kF��03�������B,＄w�]ۇ�f�+���^/�xLf�x��G������ɬ~������W�l�jկ�0��l�jǙ���G�7�_�g�����lH���=~�T�v˧��z�9>��;��4�w��<����<
D_�������g���?g��w���4����ó��F���t��5�������G���oo^��57��%n_��N�F��ׯ'��Z��������sqV~��g��F��.�pzUy�D�N��߉��~�e�t�hD�U}�]�
R�3V�C��9��"I�F'z�i؇�w�ha��
�S� f��qb6B��sH�s�`[G �����\��)&���R��Iйm�ts�bXsZOF��[��.����LANn<��S�����dfi< º4}(*X�v��Mu�Q*�l�8���.|#���~�Q�O��w$�;^JӺq�پ,������Tl���6�}�� �U���D��1�0f�U�����]�a�[lH��4n�$�~$G�	Ip��}sMn�)Θgr�1�*���b�/� ��x���C�N��DS­��S,&���ם�X�1B�&�-���?���ߙW�E��+�,Һ��µ��H~�RL6�C�����d�.���<@��6��ش�{�2��h��e���L����3o�.���*��̐VZ�HN�����'�`.s����cQ�J 2E�w��z�\�`A]��p�C�]w�o�Xm-����d~��z���������䒬���wH�-�P�+x��*��2 �!ـǭĹ��7�Z;M�#�0��܍��Ag��b����J����[����%*�#��v���gAe:�6_� 9�Dsb�e	�7��4Dy����4ƨ�͕�
��j��9�yZ�A^����9̗[/�lx�f*��G�93��_Y��[KE��)��Q֞�4]x�L�����>W �^
g�p<�=�'�Ș���a����&��
��>-Ѳ��>9�VGy�W"QO;���M�����-�k��Ϫ�oL�����u��X��;�@Њ��:2<�̌�,뒑X�pLF.��DF�ꛂ�2�4�M���B�Kk&b��#��B�{��k8y�DB17��<)��W;^�1��S�Z�Ĵ��:���w��װ�)i�_���7e���C���uq�օ�ıb�Ќ2M8��ɢґbi5��w�Sޱ�`tJ�rWߐ����$X,[K�(�j
tN%a-�'6������+@��kf��D�����e��x�2}���;3��.���i14�+��P�~*�{�sYc2Yؼ�0u�B�Q[+W66���yk�@�{P��2e���B�#�W^�^���B��۝K=0��c
�D����Y�3]f!���ēkh�̩}O��k��g�dg*
S��Ĵ����)4����R��7+�l�8-{|/έ��������-	���Nq(��J4S&����k��#ֹ�%��z�!9�B�٘#��f釦��͹�?���H4f_�rQ�%��.�� 5�u4e��J�YЀ�KKb���I���\��G�#��E����>���_$�zc�<h!t�.ڥ����B����r����
��Sx]�͵uu4̓\��c��#���i^�oM�'g6��q�(��GY��?(�el]�x��~��N����T�Z���o��h@��(J�{2���L,G(���!�Ơz��K����[|N��۰�~�I��Og�Nv�����I�Q���m�����<�R��.}�t�R@JL``&٬3M�q&�B��?�K(t��M]�X��<О�����G�uq>ƾb��o|�$
-�H����8{�6-���"����r~$'#>8�6f$k����P�VB[��BTe�F ��9ҋ���]%_�'?*�	+�ZO=��(��v�X�Z��zK����*����̙j�s7�7���Fyu;�9�i�.ɦ^kOv�z��@j��(/uX���~���'�:���}{��&�
�{�]�X���B�$�[g��$��^�|I=VS��}��*�kӠ�!f��wj�;�/��j{we�l�c�����������;�W�U�Gg_}�}Z�5�:���!�J��i}3o Y%G�֜�(�,�sFq�Fq�m����jɧ��)M����A/q钾ݸu���1Q�¬��M��A���ҧ#��-N������zR!fdWrؖҶ*�>A�|(��� ?�������4�gP�J�Cc{m{�����K���Yn%ֵuNBA�`�p�G6�	�b�/��Z��}!6��6D ��E�0I��=����g:nj	y�%=����#�{=��P�Hm�B��a������+be�^R�^&0)J�݋�����'o�J�qw;���C�J�pSh��@�p��z.��'��q��|ћ2u�l�ۘ CA�>�g*L.��s>g2Q.�{ {��^���G�������y�Vl�)����|C��>�m�!���Q�&�D�kJ��irM�P)d�b��5�y@k.aG���.]	���f����	��.��[��'#��ꥻ�~��%-��_����sb5[U��n���q�H��_]wy�㙾�ǔぼ?:ͷ�c�3�kr��'^��)��{���g.���纗�df۵�o�[ԏN�t��߶�ޮI*.�|u] D*:q�vi�Pdl�T}�q��Nt�]�(A;��-�=��}�G���ZU	x����~�Б�S���f���/?����>�VP��͟fB���I_�{����0Zo���,M�� ��T/���w,�?h��U��)���2��0jٜ+ `N֊��������H!�_�cפpG��K��6���&NR3¥�����$��Z��o���Y|r�Yn����B�[ ����m�1�5%�{��9k/ጆ*!�ܙ�d�� ������&s�Xw�����6��W�>#H����V��`K���x�w9���@�RI���ܡ���!?���#o�́�ʭ<$��k�4���Jb�U֠r���b.��Р�H� �.i6����hC�lj��c��[#�<5�K�X����[jH��9t��yr6F4d�]c�!w`�2�Q^h_#]�,jZ18��ܖ�����Z:vߥ�ާ��z����)�Mw���l��;�_X�d���^9|lIOd"ҋ�}�F��`9�<h����Y�߸-�ɒ�������^�����{8�-�u[�C!)0.����d��%� ���XE�z��)��d�}-c����N�2S\)�%���$�@޵�u�������/e�7ݺYE3�\A�߂���P��7?M%�B֒]9lɛN����yiר��\��d��R=����������h���B���#e�F�z8?�*Qjx��b �R��_��ۨ�|R��0�D���j�n��/y਽�Ϡ��9*���* sTܚ#�gQ9�BA������%S��hi5b�N+I�Ԋ:�QZ��n�3����r���Q�h��˭��z�1�#�����R�:(9��X��� �wӞA}�ys��S��I]����{���I���� v�8}[n��s�Ϸ9'Үe=�ky�H�Φ}O��=o3	��.ƴ�9|�6~#�����&���I��$+-&���`�2��7�"i~b��^�`���L��6���.3��e�r���L�P��G������7
�w��X�X}��D��@b/�?�SA����$�%rSJ5z�υ��d6��(��0�����P�v'�0R̈́e�-s���z1���.�i����\�˼�����K�_� =�0�-S+���$�06tYD{r�3�;$c��Yz�%��q3*�>ޭ[^�h�V����'�c߳CJ�&/h1B;\�ƍ\�#��Iش���8��yb�za�T�W��E��%i&��H*�x�[d��Y2�Eλ�n)����cµ�5_�E���S���Գf��˦��
ٿdE�_\4�'���q*�)��eo��Ę#���C�R9��`�1c2F���mV?�; �?AbT���դ!a��j�F��[X�"��Y�s��pG!-=�c�>|c��G7���Ǻ:�ܶ�G���(��D[�Fm�J�$�J�xfT�Ψ�c�CO���t�dg�/���j�)�tv<�0�/��6�E>�x�׾�k���xm]f�^��+98	���~��P��n�� U���8g�"K-�i�ΈGU0M��V:��͂+�5M�ߢ�8�LÞ��+�����d-��-���&��u#��B_��e����9�<�d���r�L����3bk{g)��^h^0�	��������[�'���-��F�jS��ֱX������4�W{�����d������֛�[e&��9u+��S4�g���Qh!�(8����>ƛ���d�c����5mu,6�܅���D� Z�>?/}���n��H�4#n l�ѷ��b!���Vc�f���6�FȒU���1=O�����؊��	[[�.�Ex(~8բ�7e�RF����e���v�߽�����BXJ<hYh����8?��m_1AE)�Z�����P�ޭoO����b,�閳������=۩���4�wm���δ��i�1��6�Md�����ŷO�z�f��.�u���LM���� �<A$�]h�*QȮym����Y��D髹�3v/W��揷�_���;\�M��������I�pez�ƱG��_��iA��A��҈�"o����~��o!��`5>��ܬʴ��ߊ[���$����<������N4�I�`K�a߈lŷX�Y{4��B`�������jk��7�y�Ns7��_AXe��13���2ٜ��/&�9���P����ANI�`���~�E��L�Ԟ��w}4�~�s5�y��2%�<�Hx�I^YP?H� �^j��"z��FP�Q�{�R�U�y��H2���s����$�5���;:G��?�0�����j
3(�A/MiϹ^f4X{����?oش�����J~��^��;?����]Yp]��?5��/mα7��E	� ފY���*n[;����T��'&_9��d���O��2�B�D@$I�zkc��o=b� �~S9}����n�W��wX��J���ՃIXu׊��i����߶ܫ��}4�og$�n<���{G����[��oy�m��d�]���Q���L�O���_Ј���u"��u��d�(����b.�m��\��t1�%W����8�Q�D���T���
KW�.���vw�F�=��F�חI��]7Ͼ~�^��~%��w����o�KC���/vF0����r�,J��.B����d�{"����rsX��I���2���l��4I[����4�Y=�L��)��� �l�}Cs@���FW��CK�ʆ3B' ��^*0�AD�/W���%�c����r�$:Xoh;]�%������H!��ޣ/�Dۻ�lO�P#f֨w�:eɹ�@+)���F�wM<��ٌ	��O*�y�2�d����I�������AilS��J���v}C�;P{� �ˌų
+��쨧����)Zjd+��}q���hu6:
�3Vn�����C �E+��9(������}Ҡh��w>8��܌�?g��RQ��ty��n俒18���z͍&�_�Ř�d ���Ϗ�����ҍ��ۙ������euH��_��|�w�&�{� 	��.\����-l|��3E��_I蹁$�]�4`}vPz��~��|Ҭ�n�P4& ,����x�ܦ�!�e������Dv-�v�$��8��	���,��.�'a4՛C{� `)�TL�� ��^s�Q.��������A�댘!Ԍl�xǿ������v�3w2�b�8��gI�2��t�G-��r�
,�����k΅��nA݁��y
�\��?R�!1'�f�\�l;G�2=Op(�qQMR���L�)|�P)��͎s�)�Su�Z.~��哼B�Y�J�Tђ���F��k}�^zy�o���>�תuc�îuwF��=���1Lֱ;/�U��m�t|�V@Fe)�i%�uDG3āN4�0��BA�Y�!�\H�i!} �{Y�=�� ���׿C�M�7~��T�i�N9T������@MU��5�_c��NQ�)�5r��MB���� ���ϫ�H�	RCiϢ����o���p���$������s�b��	R�ZF�5aX
~�%��6Y\ֆ�azw\�I��G�����i��}H1饔z%i���R-�f��=<�M���g����Z��>#[�����#ܪ �jH��0���Ah�RH�{?k2�4���	:�^+a?����)|-]�`6LIfV\��.�iy���2>�ե<� �w��"���ԟ��;8����P ��Y�<��a(�k��מ1Bơ�h���Z�����y%�	�ĭ�����!�k��!r����M�X��2��IK\4B+�
�&�g���G�8��0�
���	���A��x�x��ƌ�齱Ls�c�Hj��D~�r���[��
Ði
^�y+��}_��`
;N��ds.2ҥ4���0�B�Dؒ�p�������"B��9+��	�ps�
�98�~�4._P��@ߗ���"L�n��4L���� Ķ8h&0��7PP�+�+,}���%%͊ ke⼕�Gax�ڜ��8s�{=�~Sz�����`cN�Bh�4IL��2��۩���{ƹ��AFAz柊mm�D����@w\��]�y(ƶ}����pgߋ��UpHP��TH5���hwHp��kS��4Ѻ-_��/�
�ub Հ`��s��?m�p��.���g��B6��/��Ŕ�P�]���fR���)�j�T;&ѩ���3Y��⒃Wքr���>>����)���!E"p	ClǃYj�Cψ�a&F�R���2����G� �]�(m�O:���2�	+���v�ӷ0�8!ȃ\ǧ�-l ��ق:'�4� !�� aù=� z���%�>��I���.��z��RA���i�{Ӥ�LӁr�`
������;���_�.p��� e���� A�$V*vCE" ������ȃP����䛯-EN���c�*��\;��~��$)<%��ӈ���ʀm��4�'u�y�W��`�����Ϯ����+sFpD݀4���:L�@f�	c'~���J�7ɣž�<tԇ*r��|�l���_�ƫ��?�$���R2�A�vO!ˀ��ٴ�;�n�kY�}������_�Ҋ{�I	Gj��w���`����J�mLu��"�G޹��kJ/Q�v׃_����=�j�S�`�f�%�����I��)m��F���B�U+��t}��x��2�h�u��I�m��粜8����k�w��_=����i�"�S�?�5���4�̎��g��W��{fºя�"��d40�2�ɪ�P�
U (��F�|Q	��� ��B�����?�ǜ/�����A��i4�EAP&
��>>'@�u�����Q�1f�F�~jS5���Pr��\8F@�Í��·UT��� ;�nI#�qҐ�&q�K���ԋJ�w��!����xߟ��Y���go���ѧ{��e>B4%dFK�SD�\dĎm�	e����u�/X�AU:����`3c�	�q� ��v�IK ���N���!&�/G����V��>�����T{����؏O��W#`���]�!߿�.����~|�]�y���x㓧i��Ν'����C��Ҽ�䪂���U����J����r,�N?Q{Z�/G���O쎢��j�|��^���݀$ݪ"ځ�D���'m��,K��dE��.�����l��������t�h�ٻg�����{ۋ�� �Y���{'���I�ʻV���u�B6����E�Ʀ��� ��(���G��}����%ԓ����������6T!���A��/���_�-�͆Sj��,I�>��W�k!���}��X��_{7]����	0F8+Ť���SG�Ҭ���rLYR}訽2R�\6��P}�|��ҁ�S�1U$*_�9��+��0E�E�8����(3x}�|����m�Q2H�i}Z��O�纸�*�f�����_/3�5~e���b�,̌G�1����ͶM\�U��#�=�g���������p�����@tt��6�$��s�����~|�`��~���)�ȕ��kǡu6)waNM�����(��W���U���uy�j�u��/&=M�.���ݏ�E���%���~���B`Cj%����+�������1Ԛ��M��O��c)����m�2�\n�ޞ�g��%���h���ŉ�e�&Xr/�.�i����5y�!�>��){mC,��w�u �5���֭�sdY#�u�4���:P�.lb�'��4��Y���w��'f����f�g�/7�Uʅ�Y�w�m<+ﶿ�����V�-Ϲ��0`ج��+X̸���	���ո�^e�}�3�tQ)B �4l�����̝T}�<]��B>�s��ʀh�}ICL��+n��6��6oh��w<(�f;w¡bƜJRz�	v�<C�-?"�b�H��`�������F!P͕���Q��1@
�I1�.�!�W��y�m���L�
m�2�`����i����}�N��ηb��~xl��hr����%B����H�J;��:�=zŤ�;9�}B?+�-?�5!`�\����iu5f���N���M"�#���c�ݾ��e ��c-�&t�d8��"� ����V������'�fR�Ǹt�}7һEH#�_g���,�k�`r}�ْA�&9��?��D���x�9�q�l�pt"���xfD�Pz�2�E��[2%�v����Σ%��n�xІ�.<6�#��
gd˽.#�W0����7V|����c��CP=�:��Қ��7_�����3���!�����@��Y�4+#[ْ�s��0���	�[`��p�D�B��/��[�i���r���rvA�j�o�G�6�������&��|&U�"Ř��8��~�a4����Zkh�Pa�Zk>�e�D�a�)K��n�w��G,{?�al`�����Pʱ��Y�dp�/�SH���;u��'���P�叒�ZV]�01̥��toB*<z��3\
��N�zj�\�f�!'���7���苳z^hc��*K�;ܳ�ݡ
s�p� �2H7|j�&���\4��c/�W�B�=D"��G�e�Z�E�Px�=��'���KM��b>���P��7[4pL�HE�?�d��) zd��ɠ~�d�5����71�
4��8X5l�+e����4�IV'B{�rM�O�8DM��,1E���:��օv�Q%(�t6��`�8N�@�aN�^��y=���B���	���9Y�:GA*qR�>�C�f��W�]�3��6���?��-�/����y����8���ȕk;1f�tރ6�(c�܁)��� u,�qbx�2,�,}
�J�cxWG�#��(i����x5�|��<���1��-Qx?Rɢ�Rҭ�+��b �p��#��&%�����|�:W�-�cx��tQX��C�WeMQ��5�J�ܵ2ƌ,$3�2����e�;2�yޖ!�a�r���2=)���[菶ߜ�nwY2���m��B�D=_g~��%�m2�U`�O���e�&E�A�2
d��!u<�(F�[|3�	���I�J����U�"ٌ+-_�bLz�Bs��4)]v����l�M�&=2���~Nr�{�䠮7-��)�#��H۩s�J�9��24y�Tg
y�Q~'��e\'�=o:5�(ieh�U;:�d�;�'���ʳVr~�ީ�T��RG��ȯs�#{Ӎ��4����~=t�j[m�t<�x��yE�RII�ӷY���O�ӠǾʶ�D��_������+gߺ�^���)~��0�<0�TL�~�b��0��c(���o�����⍶��?{�Ț3���/��|:���A��(,�i�����$��"���H.�5b�߭S�9@�����9RV����_?��M��'����Y�Q,�����-e	���M����;*'@Ҽ���	�W@��b��D@݅��nN�T��B�,��=.@���sa���;x���hlޗf��xB�,�w�nN,��w{@��[�^�Q4R5��Zh��S5x����Smz���̘v������4`�:�nn���9Qx��h���v>���y�^)8�I�Q]}!�g�%^�N؄�d\���7��R�cm���.��Wz7r(�/�ۍЗ����i��/�'5�M��袝���n����KK�[�^[�?����3SZ쿘�q|A���h����
ӎ{Nh�����O$����%��;�6O�R�r���3��M_��-3���w>:�����#��xܴ��
��}���N�ݏ$.���g?]�����=��޳q���Me��Iw*���,Do��:ӻ�Ŀ>j�oH�o���Z>ֈ�F.���u'�&� w^'�Y9*�p�ku��,�I��{H�4(���hY�u�~���X��Ywsj;�h��Y�53�s�T��9_ʦ�25������ 	�0�!��nb��E��bx�	�q�֖��6�&xD�c^R��-ޔ�+^Q�`�r�����1��q4�h_}o�ݨ�v�W
�,.(zf""� ��A�S4k�dKw�h;J�=��9�����'���,RЗ�<]���ov�`� ̪�eD
4����9��7��U4��c%�eAv����N�K����T�dyǦ��r>�$T[.���9��6�ت��A�Lj��ٞ�ԁ�1���Uaa����ε��gL��z=�H0OXߌU�8g���=��Q��bC�����]��j˞F�����ASC��E�m�&�A���/�*FZE\��M]M9\�ӿ�� 蠢�WD�=��W�EjX��U��b�U�J�n&��A���L�z> ��z�\��8��c#ar�#��w��h���P�k2�����oGȏ�\˸��U�
����Q�e⬙�颎���웆<�@�	��
k��[���rC�QE����陦H�E\~k��o��g2>_���W����wզ/x�E@7����U�/b"���es)��a~�e<�*���� ְ+#��f����t$����C�C')�����DØ�u��N�b�����R)$������/�%L��qF�z��˓��r�֚�KPθ�e+�S=j#'c�����X��3Qj&��Ɨ�+�����j�����0H|�f>���B���*�2j�5tNp��6���`��Hl�ͧ
���:��BR<���9~�/u����,�W��0o����k���J�y���4vcx� ;"+�"n��A��":��Ѿ�mYE0�׏��̥-
_��+R�ϱ��P\��
���0�}�]JO~i0?�%[���+Y]�̷�����Q]�N[�>��ḓ��EdpJ���>�2��m]4��,��i�)i�H^�0cM��`֓�c6�!��g(ЄdE�b���p���0�������P�����hB�[��4���{���VC�]X�^ �0Y��s���mTa�T�@�p�[���g��JQ���|��-]�j��W�D�ڄ��KX�5N�)�E�ϣ/�_��w�[)
���nB��)Žu�ٮ�E�
��hTUt�*�%2<�=�R.˯С< ��^(~�BLK9��HL-����-k��������}�"��[U�JM������*�dC*
(�V��ʩ� �KE������К�9�}p��o ��j��~M�I�:d�3Hʌ���pnf���ŵ�t�+�y}�s�����f� h���+:r�E$���0	��v ��c�5��K�� ��9@"0Y�@%U@�<v�X'X�i����jJLC��>���6�� ���Yc����$P� Y';��;����B�wp`٭>I��ɗ��+�[;�M>�R�"�o8`Z��>@b��4�h���zl�"+��~��>ƽ)WS��R�	b� �jֺ��3#�͖;��R��bT��P=X�\Y��r���F#Q�륱���;D��FIdZ��(׷{@ G�������9N��ڐ���{)���~$�|Y|�o��R8poI�����ɻ7�|_�x?=兇l�H��Ӝ�8�Ć|n}9����{��χ�V2*n[+!�n
�c6*%ƃX<o���^����;��-8�-g:�j��}���`��!?zʯXv����OsIis�_�� , ���|}��)#�����L�&VhI~b��K�<�Ù��}ޙ�;�K4���Z��#�Հ���x��Fn �/B�FiP�l��'5�|8�2i �,��F}�����tn�
����v>�Y:�gȷ�b�.9~hk�5�=����������q�@�7~�7��o4�Y�[���{e�������oA~�O⭮y[���=��>72���ô���Iٮ�@�]D�Q?�+��QEdۏ3N�vH����ͣ���nӥ>~�ª�\N�Z�v�{��mu�����QE���׶��H�	�R�;�8:z����_�38��f�|�|c,�KE��TP�\�\��q�Y~�9 �N6�b�g�m>��u>��!+�р<���{u-"��EM�n�BF3!I�Ml%(7Ũ�X��V`3[#	�TrD�f6Q�<;� "�
�x���2����� u����,a��,�V�TV�qOGk�P�5���˳�n�.+��M>x���lI�]�3��p��kn;~T���ߗ�9�uڭ�_��� ����:��l��!��=� \��D��Ϭjf+�&V����>!�9���J�>�]5R�FE�����IN�Iϥ���H[�H�K���@��E�f�o~�U�w��������/;����Wz�;��~(ܺұ����w������OO���?ef�r���cw|�8�B_sx�����b#���;M��g�t=\3ٲ�!od��u����x�ؑ�8z�=��c�P4�Zj[��S�b����YU����/�%�T;s:WƋ���T��Vfk~-U[UY}������Qj�(�XZM�~(��!�u.[4�_��=6�x���8l�Ѕ�fE��r�fH�D�7� f��Ukv<�IP�߳U-d�*]P�Ԥ�m\�|���fK��S��.B�8���`$�ڒV��2�8G���/�3c�
'}P�Kׄ���0{{�	��ǝ�o���ё�{[R���Wb�7,�^2%=�y��R��A_�N���f��RMt��*��[�q��B�̽�������~Ja�b,S�,����L#h�F.)d�/?����v�cШb�眬Ұ�/����������w�Y��'���X�����#Z�/��딪&TU�2g�\,�c�N8P#,\��`Ͷ���*FZ_���֟ͻ
RMe����<��;L������v��a����:�l?XԿ��aS|lm���T��J^���ʡ>MbPO��ρ����2 �Q��G���%���A��eH��xx>���=\�*�OT�]Xi����I%�
e�I%��4j�l��!��͂�%I�J���	ǐ�#���H�p7�ܹ`P������~[hb>ܘt�j�s��:`'� g/���A��r�ܥ�Un��/����n_"�w�n�j���&ը�2���g�q]���9��_&�ࣻg���g:h6�N�'e
�����)��ף	]7�hT�T]��k�5� ��T��}�K��K�w� ~����=�M���,\W���}�n>��5��܉ǻ�푺h���4�����2�|8�I���v8�ě� ��*�d��E}H��}B�����ֈ��K5JA*�ZmѶdt>����m�L�؃�r��t;���UP��S���\\_�.'�����!��)���f�%�1=iK(n��}i?�2Ɍ�m8�3
����~�w���Go���h��<Úk��%'�7�х:L��߭�;_2���R��ԢK+Y�y\U
��dj>įL^R�+Y��	躞J���Q����B6�Ke޿qO����K�5O"��PG5�j�)�D�[�y�*;n+���d�Ӿ/,�PF:=�$!�,�DA��v1Ua{�����42.+�u��9n)�0(�����'+�Q�c���T��q�L��J��Si�a�ⶬ�;	�WLAOL:T{�"<R��n4QPT6���ǑXh쓞%^0�E$���@i��"赗0� �L:zJ0��B��`5��/\��E�y�̐�$��jr��o�G�W���D�`���d�{(�E�H�_�r�Ҙ�-/��Ofҍ#:0�&���-E�`���F\�w��Lqe�m���6��L��`p��cpB$Ge���y�2�������K���8{|�Ο��m� �	ylj`m�SJ�B,�Qq��p�S���1�ϱ��'3S�������Q��D�o1+�-o�
�_��Y&h�ޖ�F�G��pa%��4�HM!F:�p�ʯ�Ru�!��=뾺S/z?o�����z�7R�dg����d눌Nn�J.!�jNM{�,SWcn��Z��DQ�� d.i��	�d����&���t��K�J���o���9�?@�XI���*��d1���E�2D /^�CF�Xhp{��*��t�U2b���9TR�~���������ՂL	O�)6�Ki����r��[�0�5LD ��M0��
bc"���M�?���P�o�ӳ�Ŏ��kB�­���Vڇl�����A�Sȷ�����~�¦'<渖��V���F���]M4S�0�T�Kۥw�T���`x���6 ��p�wWV�g����i�R@��P=z����R9Ѻt��w��:�r'zP�z��
�1	V57�=1Sι4�t��ne[v([���϶�R '�Ѻ���)(bX�<g�
�ʇ��5�}*�F��^�����d�;|}Nh����@��Z���������=�F���mN}���(��i�L4����s���[��Ze+���q����������|8<��Ѻ��������ʻ�(��/�[�7B�;C�]<R��g�UW��X�;���F�� ��ɟ2��KO��y<	�����v������4���@ݺ������Y��鍿__��n;]�)�]l�j{��Q`��bp�ʭwXT��!�#��ڧ�o��˹�:u�{��.�v��cjG2HY��H��д?[5s�2D�V0�\�2v)��2ecxX�_��Af������e�܂�����wƴg�\Eh(Ƹ?�
��-���3��*��m7��|o���Ű���#��� ��S4@r׃$��E�t3(K�j���[��B8�F �+��|�<���A� ez�χ��)���;o埌:�d��;\3�.���X/Ɖ-��Ok�½`�_kYs.�������p@����`J���ۇ3\!�&�ܢ%;m��\�jP"i9��')%˗�����VK��_g���Px�[�������;�G��3�V�N�����������;;�r�¿��ۮ�2���%�ŏ6y�~�<�V@G�N��4��.?J��g���M���X�Z��0P(��>?p��ꓓ��n�s�+7�.�$�*��9+U�h�C�rI�ˮԒ����C�o�Ɂnsq[�ЛfIIv+�ކz�'z�N�ݩ�����@ؠs	h�S���Q+������l'�b#p��a�0�D���/"F݊��]"�X<,0G�Ѱ|�;���:����l��$p1F1�8Y�0��0��hoQ��^˓����|�o�j�oF	_y�����K]�9)�,{�Ps�vf��-3�_��Ep[}�x��T�0`���+�)���ۋ�4��������,���k��TՋ�$X	'�D���P<rv��}�T�;z�A��ͭ�O�S��:B�V_*oLӽ�]��tW���)�*�ϑ�X��c^,�0+�{p���B�M��������p�/>cb�X�(2���H.%��k�u.3��[�����:��"��~��eLn���Tʭ��U�}~����x����8�s<��N���{yN�=�m��Q4DYø,:���8i&")r|�W�3]�t�Z
��"^��:_]cn�yN�Tas�Y��๿�A2)F�� �-��0\f|[ͦH.�CJ�Aޖ���~��(����J(q����k�X>��0�=�%�_�M�[��� ��	+�R,{���J6���8(	a$0p��J%�CQx�	���,�w�>�x-�	��CS��5��첽�j�с��yz�N�z��g�:�c�@����yE1	:(i ����� ��(7÷�p]���iɶ'�&DA�jQ|+�G�sr���������;���q�E�m3b�C�9�R=�/�z�敄v�*�L*S"�J����-ϥU�]!�C���-e�LR����:��K��YFš�af�#I��įEQ��7<C��ݑ$U�����^��P�z��kX\n�2���25����3�Uf��!�)_�Nl�	����-#5h;e��.5�%g��ރ_\�_m˶u!���g?W��}C���ω�7��3-.$	 ����(h�� OJ�$�����\\��f�ێ���|�	1d��4�®g�*0RT^c'��h���)4)kk!�LB������Y0�n�-����97����q��9�-�Y�A㖴%v,_#��Dӵq��[7��o=�mg�'�$Þ!���=tKf(J�^a��LS]d�(l�K�����l7(/K�&��7�t6<G�����G|.�&�
�Tr|��\@��/�J�&�3ʽ�MY"�V!e!���
�e����c���@@uRYȡ�sK����v��C��405l����pn���B��ш~ �<��#w�#׉�ܑTt9@���hC�ԭ��>�a�L@���Ht�OM��ױ*�	�Hu�m���_��+:ͱ%7gYP_񢁕4����1�\Ny��L��t�G�jŸ�R3&�	��^0l���c�T����8��y���2��-��i�ex;?�o0i���yg:�1q������0���� ���Z6(_��+�1>�:�q	��z	_;��z~B��/�W.c���'$=�#W��;��.+��Gϓ�����Ы���ͩ���� �͍V�!.������6nP�����#\�p���%a%G�]�L��׽F��Y
�ө%5�cZ	��V�c����0��M�EU[BF�����1[J���
�yJO����U��]k� �1 Mր:e�5�w��>�Qľ9�q"oN�?�TDS�0��vR��(V��3��:�M���7���/�H��`e�yc�[p����^��QK�h)1I��'�%q��]3��������_B/�d�����G盫xc3
K|��;�υ�b?�v�Ty (��[R�a����1��<��/���~�%�A���sd(h�|�ԈqP���'@rdP_nqe�9�Xm����^�a�~o�?f�I�����64X�4�%:�$�YU<穴��Xg�]�x0�f
yQY���K�;i�r ��5B؈��6����؜��Q��������.�:'��V�&�ʯ��F�d[���f7�t;#_��>�M�*��|���lHI[�(6�?��֦`����!��j�;,8��dE��q����խ+=-wJ���[_D�<+x�hո��[�z�曙�o�_}q��ɻ�:8�{�͛��߬Ä�E�{��+��������~�Q�C�߫�}_V�ψ���B�):kF�Z�h�=�z��h{��Ѯ��VD��А�z����Â����d����|:�
���q8���}?^��a�U�"u���*���9ifOx��17vzy1�i�keGq��mM�{X`�B!Іl���h�����p]T,��O��lt�f��Ѐ/�"lt2�f&[���<.��s2,�dЅ,L�&#5�*�B��Ԗ�Ph��K��hzȰ
;�{�&�B-Y)���4��Ƒ��ԯ��\O�-�r*_g�Q� �DT�b^�x6yD�b����}.Ҽ��$���߻nr"uf����r \��]�[�f��~$eG݅��~{5�(�W���o��.�+%��^�ۦ��1��8�d=m�ވҵÚ�?�k�\E'�0�px�����ۉ@�~���G���s�eR�i�s���]*e�Ծ�	�����(޿�Ӽ�7��DY)���+JTZß����N���c�ӏz�N�'�<�,�-��}}����	�m�8��FbG�g���6ZYo�7_���D��b��'q��6�9�N��[���Rb�n��A�:.ߨ3s-�������,R�ٓ.cx��k�m�K��
�NwQ�s��są��Hx%ˆ7 M��r�	���Z	�����G&1 t3U����T������8���L�֭;�. �%�&mR2̸�I������o"v{>]����+�/=�,�>#�����Au}5�0�a�1�#~;	a�0Tt��d~5�=F�y�Wo�	�#��dK��j�Q>״N=�`h���Q��^\�$�ԝ^�d����9�}�M�|ceq��
ӽQ����S�/������B���;�� M���íC�p����D.-h�e]��� ���,Qɾa��1:���R��OxPȜ�'KI��9����O}/e,�TU-����3֭�S4�#s`�N��e�������t��SX&�4l�?Z�r��V/�����
j�ٻl�(�>V�DB��R�����ֲi�*f��UJ�ig	��*䪸����l�b�À;jg3���ͱh=�(��3�M�do��K����aL��~[��:�!<�9,SW���?�uS|
6h��ӯ������5�9�B��O�b��ԔEu��.�5)+��d)+
��ٞ��o�dW�΅�>�(_
��1S3�����q��56����g�����aM*h������-�xa܊J׭���=�u�9�Һ����}�[jv4r�ė���z7s��$�ϴ�����55��2�S�' �62!#7�]�c��O?4.Y9}(�E�ݸۓ*q�6��5��b�f@�R��FK�Lf���Abu�!+#��R�NGC<g����*��MPxH��}��
�4w�,����B�,�5�2K�i3<t��ʵ���"7^��,��kb��nj�+h�g�@�YTz��:��zu˥:q��T!���I;�rIr4KH�Nv�o���!K�0�������DٵE�}�D=�$
�R�s(��_X�м�x�ױ�-��ǙA�"c����j�шz���Ӹ�g��R
G:M]pC�z���&,n�|\�"}[أ4��'����"ۇ�~�H�W3�zz>I�)�ai�1&�Q4��z6XM�Fr�ZWl���s\>���l~�6�E��6�+�>�TѶ��^�+�K��\��K�ie��m�O_�"��A��%Ky��4�����T�����;�כ+A�s��s����]��N�,peHS�x-t�k��KF�2��U�U�)I����L��y�T���1�E��v��:(�5���T�߬�Y�e�e���{7b�*��iD��	 8S:O��J �{�q}6��<=�Ӽ�27�FD��\�������i@d$�lL�P.��p��^�<ԨǁUQ)��8@�1�'�R�AWoY��w;��\p���Z� �f�j��ڤh�U�H�z{?�ek\���+>!� {��}� �%�C+K��Q̓��&�e�
�<���O�sQ���0����	�?8�C��^I歭"#.�s�����f	�X(���0�]X|���h�!�S�
@���)���x�u��~���B�I)�����qҊ�-[4���Yp���Q�]9���4���ox�_n��[�$�#`�:���w�� dY���p8l�]+,�I�8>�'�O�:�C�J��hB{)6�N����vvv�~�#�?�P���b��zMN�[��V��*���yQ%V�$�n?1��n�ЗF���F;�[I+Qv��Ț�;ҁ�e)�l����� C�QQ�<�b�9Gȕ���L�.�)��g4��yZ�T�C�E������!����ݲk�w887Ԃ{��(2��<�����eڛ�~8��n߿��;�rT�GCܣ��Ůq�C�Z*|���@ /4�ft�|���h�}#�	��_�!��x:>5��Rn��h)�nm��gz�m.��w��L� Ч�q�;8&r�+u����0'x����C�����������K?�K���p+���v�^ʦ�ý��W����~z�F#2�|�cy�R�þ;�G�Ʀ�gW���N��Gg���o�Y76�p���;Q�➣�Ko:�
n��������ϧ�=�>Ov��v�مO����>z�t���ط��Xr�S��B�ҍ7ŷ7����YG�J
!'r�#_���`����#
Q��$"w`�¯�A���Po��{����ٹ�|�=�_�E��pV3O�X<�3)д$��Rǡ��i׿Ab"ێ��u�A�4�?o��)]��O2!U�����dƻH��`"V�J�=+����[�R��
�&�`���
/t�>U<2�c �HA�^g�H��gv$Bҿ�*,WP�ԗ�o:��[?������V�[�Э�(4n?)W��E~�)��h�%�F^SHx�	�uHZ�#*�UW��Lk�g��He��@�~��d䂈L�N �#e�7>��E?��h�%}-�;d�q&>H���9>���V��ϯ�[�����S�g��o���tn�����4M��c����?-:�b�C
��%��Y���y���ӿ���#�b�VhZ�az�ݿ5a��iu�u�֬���&դ�S��[i�}�_���`:B@���#��)��U�s�����o �!��*��-�����͖uc8EL�c�A�n[3�/�P�&.�-VėҠ����?�9�C��ɯs���zg�}�@}�y;� 'q�JKÆ���؎��n#ީ/Q��y��O\(if���z����a�=�7��ĸ�Ҟr\�#h�]bK�վ�(�s�w�vjO,i�P&�Y��K���÷|���9�M�b��B��!_�O�q�������>�v��T`랙O�T���Oy�bS{I����IEݫ]��dK��囈��}6\`���δx��fP��	m�w��r�/��
�����]g�V�H��Q�H��6��iђ&�L���t'�,-@� <([�N)�>��0���w.�F��r�-|c���(�`�j\	�f�4Gm濝��ߒ�!y����(P�����+��N�xZp��`b�,)����Z`�Fpw���dww���0QY��3�b
۱�]�Z�� ��n&��30�hz��؝P}.Gp��ږ� �Ru٦���]�hԮgX)Z[����|�rE���N�K2箉��5��-h�.���jU���o={�5��dMC��X��''{�1fZ���M�r�Ṻ3��NnV��'�-1܍���#�/-u1Ov��rAK��zĮ���S9�N�`��;�a�!�R>��e�N9E��ݪ���v��-B�ij�FF.��;F��l+�N�Z�S�%'�>�5	Ԃ���|�D{� d�\�L��T	l��f�S��1����Ȇ�S9�z�@jK^�`�`�F�����g�ꡥ`����5�A떪
U�p�� /�yØ�1=�:kD2ʻ>���N��R=~����)��1�D���הTc �Yb�![�ޥ�t�O(�'7�oŔ�[�<}՞yC��^�R�w��ٿ��38{j(g���ϱ� �0T���a�mq)K��7�BIBy?ܶ۲%Pr�k�;�\nML?уB?�s6j�Q�̡���� s:�R�|�>S5�F
��'j�V��X�X��o�����{�N��gDQy�KT3Nb�����>!�π�'�]/�V}6�(`}\�^�K��^b�'�ϵe.�5�әHt� ��lq;��Q�T�	(�O��/IV�/.-��x�c�=�mAӟ�6,>oXㅆ=fU3�OԻ���\�����}���G7���d�+�q`��%�I@�۸�h-@��J���q8{�5F�d{Zk�!+�$�\��k�}���F���l�Zoe�wM�����ËQj��|������)����4%��*z]���Ɲ��N��2�����s�U��5	f3�Q1vLDOS�V����Mp�#[�ηᡲ2tu0EsU����Q� ��!庭�lڶ44�h����w�/�o�1���4 ­�.�7�'4����E�&�L���VⶁP�=���PE/&X���i�X6@ր��#�י$W2���Et�t�p�J�U�_}�	�~Vl�1�*�U����.�H���R��aH�_���t�©�+������0�c�j�0x\\�k#��n�(���ˮ�m���^�6{��捋]�U��i�����q�hB��*���b�g���F�����f��|g4D��V��}G���~�kk}i8�1��]��A4륽P-"i!�/I�\�b]�=�2��B���G�>��A�=m"��S��P� �,�XP��B��nț��G����)t5 ��J����#
�P9ߝ()���ѕ��Q�d�	�$��)��ܝ�f��[��}����YMD4j��<�������ۺ�A�E�!��}�_<�}�J�f��֟?�~7;�l�Y�Ď�Rk#�Y��o�˸��[������`g-:��5���gP�ީ��A��i�0�ꟉP������7�w7+���s������y��; ��fw(�9�}���ؒ�:z���|q�I�sy痒�[�������n�6���T8r��FQ�c��?�b2��g�:jV0��'I�CJl��Q��h��QQ����os�0(�X���(Cl'��X4A���%	N��~Y���/s%�v��69q����at@f�?s����8��Y_MwU����xEDl�V�7f�E6,����.I�Z6�>\`��T���Ƅ�ܥ�����f+kR�`�|����Qr��%P�F^�iW��&'5Wr�c2���� ���\}�3��|�.!�jN,&��=�;�M̄�s`.;?�'�-�8%J�r���Tތ\��G#���)��}�!�ancê�%�ְ�v�R��68���<��i6p�0w/9!�V9�e�L��f7I�'���˞{��/��ھ?w{~$4;���o����[�X���k�s�9s��M�}O�z�h�����[A���)o������ɜҴM��?Vz@d �
�䋟amMnk�q��1<�;g�p8pVW�`!X ��{&{'z�������n�6\�@C���YYi��%���u��?�n�FZ�x���v�}��Cp�gq=��`.;�v��M��'xūR��nqFlEYH�ٰ��fv�L��R�� ���W�?��M��e�s��MK�Y�R�gs[>��m���|ɼ�����)��٣�g�%QD���o�R�pWm�v�S�r��>W�G�P�I��.��:���ɻ��$�J#�eTP ��Z!��R:s��p��e���ٝ����gwZ� tP�G𔍝}������k93l#ņ���wo���������4�|�W����Ћ,W�<3��/!}���<�?�,�g�U�
X�nǽ���@���QO�I�1J��{��>��[[��'n ��>�Qy�	s��/x�zZ!�����KwB%��.m|�̘\�)���M[�;�����l$c�5��M�F��xjh%�I�{4��X~�L�.>�U�~L�V���1��I���Br0�����#̡��bΕ�ˮ<����Y)i���7������5]�/Q(�����W��d���_�.�1q�Q��eL��-�Z�E�/�{���3��D�K���+r���x[
������H���b�� �������l�h��j��|9�2f���a��B0sݵ��3�d[c��_��ĩ
�������[�F�!	����]�u	WC�������%<�o��^6����RO�\�P+GC��9��:��0<� ��-��m뉻<�f�mx���ܴ�B���]ן\�&ZH�iZb�W�G�@�k��=��GN�МP���%�qO�;��U��6��(�B>b=�y��2�&Z���y��'s����6R r�,K��J��t�7_�8 ��[g�[�臰�����Mvl�嶷W����	i�pU��|.T����Ms0��c:��PP��%{K�*�����b�ߨM�����I�ZR'R�!}s������Ӛz#��9�(����^�
9t���=�,�F������w���m47m�()3��� Ԧ�ҫ��9=�����\J�����H��=jJ��筹6
��E���z�`GJ{]	���Ⲻ��G�S���(�}���f����І��p�*G_�4m'�$�e���Q��tt��u�R�oJ	��J'��}�"�j���i���K1��ۄu�E��"9� �CTRJ �aQPb�\a��Xʴ�}�Ɋ�˶r�y�Y�m_͆�Γe9�,���t�T���8��AרO(=^$(��~��5�P��dO�jK!_i��x�mc7��v`M���Ivy�<S�OXk�7S����/@���9mw��`I����X�_Θ���ѻ&l����6� �$r.�!Z�#u��Y�!tAB!%:�إ5��c�����JZ��~��/b��U�f-X�r0�!m��2J�_��N2x];�Z�VP��[n�`�ۯ/Ҋ.Av�*���.�%���n	H�ʴ5��͂��q��n�w�\*��fWDm��x�qv�M�|�F^w���T��O�R�;�/�RUWU/f��<YV��j�b@�pצg���tT����uE��t�{�#���xd;J
��jvV̉�}�8 8���	q�J҈8&���އv7'dƨR��#U�Y֨����{�&�_TH��3��	������l�渝�@�D�?#k3K���R�#D�H�P�87�x�پ\����a	���0"t��w���s�R �Od�I\������߶(a�L0�A�E�Q3��'�����4���[�k@9��Zw����hkI���0_��=�d� �Iy�'�Y��;��sW�T�D�_1��ȱ���j����ÝE?�ip���a���u��C�qv����3_~��+x[#9����_�g���<8�ؽ�w�x%����ԣ��������>ٹ^T׷]�r��/z;(	�a�*��m�5�Mw������[�Dwh����t�C(F�����)�M�^{�SAk�i�ʣ��-�3'��è�?����a���GA��ֱ,�Z>�)��.	������ɞ$we~�PW��?PVĠfsp�P���K��0A��(�瀴��e�J.��=-D$ә���	{�b�[[�>��Ȇ*`��Vy�Q�_ɏ�����oNɼ,Z¨P��v$�{\�N$C�\B�8�y텾ܪR�.wPs���6���8�
ª��������o�k���T␒�z���>���JeLs� k���r�������wƩ#֚}����\��zI�7�2A��/�.�tv<��v��PK�*(t��d����6�� ���𧻓�C������۸hwg!�ȋ�s��0a�Ʉq�z��J's��Λ<�&����2�!)jhKuu�A'�C�M�`vH=���n0�'��g��Fz��������Cy�-Q]!x'�AX9{�Д8~m�xZ\@'i�
lA.�����W��~R�g�*��ܰ�+�y��%���X�	f�}�L��bIՅ0�∊Pe�BtJw[毒�K��ڔ�����?C����~�:�,�~I���"�yz�c��F,��|���0dwu>+!{��/s"�a��T�X�Mxs+(��,D��A�Q��ʷ��>6B����l��2H�!T�e�E񾱺0�b
I��{#K�#���S�����.ݰ׍K�(���'�xrT����/W_�K����_BX}�'��Q2��w����U��Y�O?�8wgo-�\��I�?�0>
9�a{/`a�*�XWQE��w0��r��ͰK��쾼�(U��5�V+���������s۶dNL�q����j��y��ev����j��}l������g��Z��bCx-�e��2�C�r���x=�lYs��=')���j <��"�;w�K�����Ҡȸ����n��Fx"��Ҧc?��8Ҙ��?W�T.{`=꺖/���+���`��Wuu�� �J��\�Ԭ�����ɹ��ރ�����<p����3^m��<\YjF�x�X�?ݞ��4Wә��ii�x9O�1�^)/��o5b6WZZ��wC�;<*�S/��m��IXrY��w-�B*ޏ�����7ݓʮ=gЎatU�e�_�>�]պW���-����u��M>�@��3�E;�J����K��Y�$5��q��nL���M�!8N�"���aP��#L�F�1�4�Ǉ�	G;��g~+$AKih�W�Q����	�_�ꐌ��n	��A�+��l��SX[�B�Q��L w�4!`���O�D��=m�v� �`��m��| |>p�݄�ߒ3R�0$Tк�d#D���b~��?3�ͪj��?!�&%�Z-\K�=l�ZY)�	Ʒ��m���%�Qt2Ɠ�kEd5>��DD�H���l�񏣼r2'�]}n���N��&+V;��.��v��GV[���O����a2�y"?l
�ӛ�j5WԄ[[.�S��>@e��B���^��#s,��	Ib��-��,~7l�܇>r�7��zmI�܋�Q���g�Sc��*�*���TB_�V�=f��q	E�UF�$���ʼ�!��7�;*�+{zrO��ZG��\𔛴�2�1k�M����}_�4Ls�����e�*�a-X��:R�\|C�M�8�;�]�sV��`�pf�js����Kq��;;��_*Ռ���7TN.Y(� ����v_�S :�2��$`&���Cs����Ʌ�����k��r�e�M�f�g"��ڀl���ͺ�$n!@챓L��"�株Q���Jm6.}c~������H��,̌��+�&�u�m��,�P$ ���r*A�[^X�֗��9e'!Ͷ!�h�#Z���L��E��v�:��zߖK�a�ԊM���� #*]P������p6�s�w���c��U����U�ؘC��H�*�Z`��� v��TA�|8��ULr�olB�k�[i[�x�M�p՚� �Ϭ�SC0�뼴�@�߇��vLER�Z��neut�>g�{'?����b�IX��:2}J4-L�.j�]����z
�zC�Z�p�5�+�!0�Bn>�}��0��v��%�#�RߞXol�@��rk�v�ٛ^_�Y1���mq�[97&��	M�����8�LW����21F���e��PFU	� @b��X����R�����j��/7]�X�16N�L��m��h;�x�Y�t���,}�Ŝ1Jx���]`ݲ�2EdR����8Y+�����x�<E���\�����Nf
�X81�uTS����qP��P��A�*vV��T��F^s�g�#�ers #��!���W����'��� ����Q�t��̇G(�ܒ
>��]�O�<�dAkO�W�����8�w)J�')�����Z��7�u����ϕ7=�����n9߾�yx��z�ַ�[�CW��7�5p�����u�Q��Ո/�ڎ��w)�(~�(���E���8��T���jZv95�Y�1M�_����ro��Ҍ�oq���e)�Nw�?ۍ[�N:�Q`�v#lSx��Y`}|FС�-�	��\�S8����K}�T���.A��;A]B�E��Rn��
�;R�C1m^r�.y�#��4�hG�kT�6����K��}bGbf*��0����w�p�KUs��~���4����2+���0���0`�n�(��F���)���gW��$�������J��*�s);[��.(�ѫ E�X٣ʄ�+&X�ٓmC�߳�+� ރ�s�~/d���Р�@W.8k�VGj=�dg(���;N���WR��)�O�^����8�2%�����G2��ǏJ5�2�j��63b��������A'��x4�]t���{���q���l�;a�9+�^tbg�;�1]RW;��E��7u�3���,f9�|J=F�ԍ�L�Hĝ�)17�O�+�ZfO3&I�1	� �����q�,Y�L��MT^�Ƞ��Yk�����ӷ�]��_�G	o�R����.v�3�U�����sV�lS��uƹL���K1/����a�1m�}c�	u�kˎ7�[����'�xa E��祇XD&��o��_E �̳��8��t;u^"�X�����l�p���X��xD����o�)�������RBE0�"Th^��L��czｯi��$�m��u���~)r�h�։b�[�����V��?Y@"�Q�l���N
$��KT�ԁ~�u��_�H���Jz$h:��1����7�_����/� �a�o��O�&Z���|Λ���E��=x�y{��}M�:�w9؁\������+��#,}��x�������Ò9��^� ^7�X#x����\���cso�6 ޜ�.�_����t��"#�E�ʋq[W�Cn�Ie{a����)�9�����!:�vu�������=���h�tmP,M%s��-�A������?�D�_X�nD��/=����T%�e���X�2��&�[�/�#�yv�ޝ�~���z��e�b������Z�g8�lc��?�4�����UI^S�,9�0��m���{]"~N��3���b�\�9�}.���:��)16Dцn�^#��eY#X�z���BS�֜�X|���o�z���.{��, {&�<�m��)�r�I��(��D�����p���x��e�SZ_���R6��Њ]��u�D��� �ܜJ�2m�#���\_�
^�1�f��[�vܨG
�]J�[Ė}&2,d�3@�f���R$���>�n.�4\�p�rYn�y>A%��˛�vşſ��NWS�D͵������/U4�[m�߿�mA�(.�hڮ�elқY5g�U���N��ċ�
�ȘM��F�4W��5[���P
hS�o�,�jJ�1��ʇ>�:���3Y�.� �$���=��>5�@� ��(����u�e.xǉ���ɰq�����^ ԯ��~�ї_�"������ZϘ��H�q]w��rI�Y�VN�AoT|Lvq�����b�/��N
k���a�3�r6O��R,�� -��QV����;p�����qe߿�8Y;:�+�:�(XYT�4���y�ۼ'RQ#�\��f^ "��������-g������c�=�jۚWhUL#o�!�3���o[Q��Q��N��99'��Y6�n�<,P���e�Y�ɞ�q;����e�<�wȹ�|��QP�a��BZ����:�ԮR[�k�h�[*w��0��֍���
�X@�|uMW��)q6�*�5�� ��r�B����E!���������xnZ��.��$����B�(�V*��b~��P��I	����m�@���/\��	�~���U� SA(S�QU�yz_����.Q�����&�M˔(D�?������
���r,�`M=C�#���4Z6�-�VxZJ������UX��!B�W��V�w��,�lc+�")҈~4"n��Fv Y��x��Xb������
;T�Ar�YZ�l�&P%�i���fDꏎ ߮U����f�f�����'H	zx�Ӥg�%˖��VW�B�'�O��2��I������ף)1�~��� �5����Щlr��p����o��᝼h�]��lY�G���M5u �j̯y��v7���ۙ�>����Em�H�?�JTr����Y���&U�<6�g�T�Bn�����.:'��lCɧ�#�� �L�:��׾-2�>�@α�wu7H������(O��d<�v0
�y[��l��u��H;n�&\S,�ͺ��z�u��1���ʹ���<���g�޴/����ͣ���nN�5��0ܲMMk��T�*���ߞ$m���dsﻛ,v�ӊ���&r��ː�!�x��m�p�RS���
E��a�C�ԅ1?�,�H�+��E��I�^��͞&���$p*�*���y6K<��T�f�%�
|�i�>�sb���EU(�����CO�F��ۊ��E"���K_���z�1\qaq��ӣ�_�ٽ���i�%{۴���VĄh�u�򩫺]���	^�=u浝��̅X~;"yc299�ㄅ|���S��y��;p�+	AB
�A^}vt��E=ar�#hj�)���uU���ø�P��KP�����.43��Z��;+���H!��{�/��ox-�p���o&�ZP��Ç���\�y7A���+���yi,p�88�]�G��|��C
�V����_��2{�S ��%ˉv�l8����ۻf*���Hb��ƪߊ�nO��)1A�#��Oye��t�M@;m�א�� m��:����5Vx��ު�#�WPyk��pM����h����������߹��xH����\i'�˽8v�%���A�Y�rg�9I/F�_�{�øC|�i�"�FblӴ�����!ig�y7��+�ϱ�tE�p��i��fЀ>F���/���S;:1��Į')��l|)�s(�d����{�Qʨ5�֖{W�x��_[�7m,ڤ����Y'�g�5PB�����2����Wg�� d�
l:1Y�Z7���>V=�Y�\xe�Q-�] �y$�(�̷�?�(�)��`�L�`M�٬A9)�F'�F��C[)�����|�2�_1;�H�-�:�E\(���T{�!�K� Zf�����;��)���@[�E���8̔ "�
Wӯ�I0ą��]#��l�d!�4��ݥi��n�Y�-��S��N7��-��~*�<k���9�.��V����tB{j�{��w�a�;�(��C�������"���7�_���2�H㔗L��}�i�\����\�t����S�D�^J�<��v�=���d}��\�/��w;u�_��#A?�/d�,����[��Z��$�.dH~Ih��H[���Y ���Y�K����^|�8�V�>l�=�V���i�u���w��e<�tc�P�Xi8��R@N+��v��5�ZN|�mE �3Ԧ�S�*z��������L�L� �b6�`�U ���W��hs#2��m`=�L
B�_Z4��T}����}��Ωa��\��O�����$�Qa 	wJ���M��i��+�����ɠg񳗦�f��qv�!�Wn������������3�}Yw�+ŀ�3	��ƕ�e�K]��P3����sAIq�LnE�~�>t��8t����:���L��S��	�YGx����(��#/�s��2p�vq��:x��$��w������j�10$]x`��[d�p�u�		�j*ڱ��)��U�o��N�iDl�^f��/��sC�}�Q�V�#�����W�Y���y�����u�S�-���ʏ��z�B{����9�:puI)'4g:�:�Hv�ޛl�N8R?��-\A�ܜ��.��T`gD���`�ˌR|,��.�H�����릵�v����4�H�_�Oa�~��ȧg��KH�%k��c#�
أ+�꟣�p�������)
H���Ͼ/�5���o�g���		�i�r�� ��L��}�H��ր��iᵣ������?l�D y�z�A���F겆�Ow(-�|u��*�8fv!����s��ʈ�aF�:�^z� 
�@�� �9�g�T�����XJ��7��!(�U�vs2�[/��kͪ
d��x���g���q�_���>��ჱV�1o_��:t���%[�M��?F*�Iv�F޵4�*����@�tG|��W�n��e�Y��n������R�����kND�/"�#���H��qU^����k��)��c�b�	��9�0��|�I���G#�>û���	�n��e���\���K�g��c@�Xm���FЅ��������VT<W�L�T�%��j���`��-4��-��b!�S�;�ڼ�[��(�I��	���*����Zk)�iF��ɭ�X�#��=�ݐC��b�^&����*]��d��/��n!Vo�V�N֗���!��q��s����-߁%�z�w��"�IH��m�����Ђ��\���t�AM(_!����*]���!RB�Ыz�"U�� �BGz��H�ҥK���DE��{���;�g�yf��̞=��L�C�?9;��R�j
�T��0�f)�$���s�-�:��rے���|��O¨t=���AO#%��a&>�wKP���)�c�!�W3w���Z���W��CR�Ю $��G�Qב/L\ c04��(I��Ϗ�?��Q:M���Yo��\b�I�fXd�y��K������U;-djViP)`�̜A�4�f�kv*H��YrZ���*�տfJ, �����OHfӽ�Y���b��
t݂��?nf����-kę��E�K$3{�˴\�u����:	ˌ�RV;P�/��|��+�h����1v�H�[K������� }������f� ���t�;*�-Q#�3qjxT
�8nāO��L�W�$�Ŀ���,���dN�/ ?M��B����LV��������o	֦�\�����軮�A����p�y�a�{� H�D��{������
���4��$����������Xb�� ��	A�#�F��\$�т��i5�!gMFiӽ��G�W�kL��;��?5���}����=�k$Vmd�Kgx�ӣ˯|���v�$�,8^˱yB"ɔ����p�g+���?��a/�����}��bY������嶧�S�����g��Nݗ����?V't��)꺕�7� �fװ�b��k�C$,��$O�ŸV��T�W�+�g&]�Ra���N�B�(��6�9�ms�\�qқ�"b_�5�9K��M���$أ�ڽ�ہvBۄ��
��6��c�O(�������Ĝ6�������	�ׇ��"�� xEh�	�a���3�(�v�i��ց�]��Ey�J��_��WH�#K�%'�m"+d���%�V�g�ܰ}�O�?�J���3����z��N��SK{�P�%��d�JLEBz;�'���+J+�� &L0+�G�&6�7���'@�?a�^�21a���r��L[�WE�4Xz���L~^A��A�������(m.@�;H=<�8p�Fm@�P�� ͱ����ѮO�^�_2�&���۪߈�D��z��z�2�mtl���:<.%$�B]��v�3K��j&�)g2)5>�K��Oj�O2ۍT�i�wP�0�����G����M}˼s��Ŋ��	$Og�A����d(�cpd����N.��q��|۔AR������j\#u�޲ATq��`�uK�9����ͬԕV[����[r����n{��{����0��{��=����Ҿ��Uj_���7�~�i�iܑ�4����_��'���ڊp}Z�T6BD�齍����hϚT��$|����:��{j��lU�$q�������d%��ׯ��������X��2D�|b�얰�@��zjC1B�Z�s��hM�<�:�4�@%�o[��Y���H ��ȱ�x/۽����Eݨ���7�<�xM�S��3��g��$�@�")�'��YNK�r�<��3-e~��A^���<x%(�ĶϿ��MQ.���f��GI7��Y$/K�[[q��G?Xز���,��}1�s��
h}I�(0�ag˗�Tu+���%��I=�b�A/���[rn�h�����2'�_��!�@���O����"!7r�z̖e� ��m��߳��EC�c@�F�.~�w�+�l����fd���73��|��_�ƞtxv9m��Zà�3X)�V��<��OΧ0�Z
��ݒ�8"v�)�)�xT	�����e��t�Ja��S����A�e���a|,n#޼�e�`rb�������8`I�8R�0�⫒�����4ɴ�F:���D�.'2u�d�>����ca���4Ҫh���M���h*#}WՄ�D��pE�{������M��i#m
,�Q��M�>Bk`���bO��Z��N�h�(�ݖ��C9�j��E6�$!gA������ą�Xz���9`�"������ai�Jg�3�	�R}L���0�	��Vq�Ӧ�K��;�>�=ḯ����c�K�z�A���bVZ��@j2tM���I����OSiQ��p7��	�f����ؠD���\)��"=���ؤ����P_L/#�M0t���b~�"ck#,gQ��uk2
eo�X���pZD��1�vf<�'F/�1��qbw����E8�e�����|0-A���.+�m�ž�D���<h4�AC��n����D��[����U���Ɣ���붣e��Z��o�m@�P(��Ϸ��л��a1���K� ��5Έ;l��/.Xc}Pg�b���P�Y�E��Ui��nF���6�6���܁�J�.ߜ�yKޞmm�L�a�/��͐�j��ɴ1��bU|q�Y�y�z�t��z�p
�5�#�h�H�%��}�d���&��Y�_	�7z�s��� ��B���
@�����y��N7,����&��];�T���bd�PL����$H�� (�P�X�04��ZF�?<�$�MR���sHK��ÌS�.�_���[z�p)�`]�n���T,������O��{V�����*T���a���ܙ=��4=�kZ��/"�n�w��|�w����oj���L�m�na�[&W��L��)��O��	���ky��jnߦL���5���"�	'*;z0&�@�m�'H9����36Mz�GE; f��鎦<4}���4��j��T���rA����p�P���l�nJM-X`DU�0�̊��l�dzI�є
�"�d�Q7$p7�� ؈�"��8�N�e�m�c�#T&�Z��L�.�'A�Vd��y77١�Bi�,����#����G��Ufe,e������\���S6���Z���k�`�.��''�#v73��&;�����b+�d�w>� @��=K���S�#2�M+��������̤iA%�/��Oz�m#(f)�(S�B����	���ŷ��:����7�x�&'��"RnI;��!��O/���g8��,�h��F,LBFUwL�^����V�q�:ŁnaU����X��\M%��^J��"@O����*2�Χ+ЏI��0_}+a��+qh��_k�b���?�:�Ӵ����
���Lt5`-#~f����\)��̚�^�=�r��ﱿ�9�[_K�1��>�N���'#�����U4�.1�$��}�7��|��6b�<��0PW���
YΒ]H��ǂ+�A�ļ�c��{�po4ZI��� ��@�[�w8�Ӿ3(�
�E�\k(�dTw!�����Ơi䷖��~K'xR�_��y��r*C�G����ߗ��(N�b�������I��#��Բ<���c2:b�*�^GV��e��B�k{]��C�X!��Y������{���b�7cU\�Vm=�h;Z��C�h/��{���[5/(�4��a:���%��E��	sh�+�k%����d�����&0��eW�Kk"�T��upQ�$�Ơ}��n�(��.����v��K.���{r ������^P�-�0m�n���?�����/rp6nu6�ᚐ��ŸI��w���h�`���N��&�y���~��F�|Zuy��ϞQ|�?H�"�
���X;�������n��S}�]��u�!/�"�A/�Zf0!����t~@ϔ��L�ZX��v�f�qF~�}Z�Jp��a�H�9�c;��ڴ�âd¬�L�����c\
�1&x�@{��4����% �j�sQ#� ǖp�8���L�T��ݔ����/��9����tp�r�GAG��p�:�=X��y*Ӳ���|����z�˥�J�Cj�r�މ��C��^ 6�؂�4�t��4�;O��(��T�\�q%PF��Q�itJ�{�E��}�1A��R��ǋ�:�RL�X��b3lϒ}���䋸;C�P9��F��ԭ���JjQk
0�_Y��o"B�h�'�D���Q�_C�ٯ��N������6�.�f�#�%w��R#!�bb��R��y^�
#���

d}M�gJ0Īܳ�݃�,� E{h��OxQ��Fh�D*����]'������}">�U6��d�H� 9!%�� �ַ�jއ�)����t�A���c]{���V��|������C�z{�!�����j�C��y��4k]�ݛ�P=g�S�ӟ,(�Z&�c-a�vtN�D�8ja��`�Y9v�����]W��6}�m���UIl �J���u���=�xJ����R>i�gi�\�mサ�*`~tݓ��z�UlЀ;Z�7ZيrO��v?��gN-�7Y�Z�+ڴ�#�t��Z��i%<�!h+h�w,H��W�3L�^J�ǚXE��~$���W����.$L���ݰ �iS�RL�B� 5��$�Ȃ���H�B��`���%���Q��.G����~�Q�37�Xꦲb���4t�3�+o�b�E���3c14F~���^]����n@�5ff�|��ೈxcHtd{�؉Ὃ��W~p%�(��Mb�� ���X��l�����cE�'n������=a��4vn�L�y�ɿ�@iG��[�4t�H�ҫ���n��Ko�$ݸ�r�
IG0=yY����t�����;�v/e	iN�8���?��v"YG]���Y���mw<1�Q������SX��������z1���<��Ky�8s>A�1�Um�= )䈷Ҷ�Aj*�ӡw
�03��"��p���6�n�{��bVeW��_��J۳���ۧik��!ڥ�p�`A�Ò�%�B��pS�ڒ%����x�_��#Y�������/�Z��K�ڹ��rÙq�c���b�p�z����9�&/�a��t-i'�=y�����Y�k'3��B����?\Ȏ1�Ks��V&r�_��DA݁���2��$��o�mz-�
>�1����__��\ޭ�>A/��3��~ZY�&�X�Gan�����1q��=�)�Z����əMqv��q6_�/�+.��G�1Z��0� �\�q���;3��^�2RPS�"�$BN��z�|C��5�0����(^����ooIj�b�럀gIҫ�J 2N�W\�m?�'[C{mjr�(rW���ut�b�z�b։;DV#��e+��n�8��@w�M�"!Tġ��f�Fqs:9]&M�Q��al�3<^��/���'+��#7Y�G'���3�} �l*"4)� �$V���������&i�0���|��79�N�؋��g���R�P22U&�.�k��6̓g<���n�S鑰����w�a�<@V��bf���x�,w��7��1���'A��d,��z�Z����o*�<h��F ����=E��Օ17�}�����B������M��.�(� �a_�$!�ܫ5�h�M�r�j���3e/Lc�F1=��o#w�e7´9�� �gf�ϡs�R.t��⚌��i�j�,�p�=f[�(hz��|�����+����f1ދ_��k�� )-�\�H/�Ѡh����g}���Ջ_`
e놓8ɄBA��kڪ�$M#�� �z+�N��r��5��_��w�z�;�1j+ԅ��uFII�g��UT�7 � �e�l�t2c$�z���Ϲ&��Dq ��ᱛ��|5���hh�=�`-l�����f0�L�=�/";��:���&������du����o8�EXH���rh��C
����v}�OѲ`.T�߂�w�M<HN*�$O%�6c'��M��f��2��Oq8.V����LWu/s�Dm��{g+�vX�7F5���ؑh��;���"=�b�.��ZnU_�tGo���[�͇���w��MO��r#���|~1+��XP��+[iZoH z+�q�pm��F'��VZ��,�$n��lj�F��0(!�������E�
�ꜧ���L�C��f�`�3A�?x:xP���ך�N'�����=jl�s��g"�,]�I�֗;�d\ɴA�4�}mVl@�'X�-8!����wpFN+�� aS���'���3������w�R���A�P۠��r��tϩ*DP�f�r���E:�q���+�8�)Vv�Sh41�g~P�Y��YY��4���WΩ�w3��M� �����%<TZ�a�����5S����'���O���(���C.v�)��!T��|&6
�hR�A{?<��Q����o��l�(|�P�Ϫ{�-г�z��M�������Hg�ަTM���|��v_�A���^OΊ�ӭ���Υ�����*����/��|���ԇKN>x����貭�4YUb_Jj��
�����_����D��n>,�m�	�o���S��17�������$�wnqL��;���7�	BlJ׫`����+��b�è_(zA(_)(���s��}O�{V��\ZV �8���������R���p-Ӫ�&1Et;;k�d�,���&�$�:tӸj(�C��|sS����L�ԳRS�C�#V6� i�Y)ș���B&)\ ��ݼmI=�MCZd�KI��yF�I�X>�1���KV���8$T��I@�,�*AU���i'|�����Af�(�Gz7�a�XEk��;qTI�Lp����y� wi@�,'�ܶ
3���<��9���y�!���eG��:�����"��J��JFU-�>�*��_��`+�+u�e�� ���{��-7�S&�B;�Z��?
T ��^�>乸�_�����59I�	�Rv�z)to注�*��Z,�%R�t;�4Ss��������ܻ��������=���<w�(&ќ��ix]=�k/���.`��N�F"E�W
]߱�yP��=�骣;�&�b߲k���"������~r
G��Iy �z6K�z7Q��2V�a����3��'�o�:�����=hˡ�ɧ�I=��/F��&�A��e"}8X��9_�n>�3�}�ͰdA�v�=G�Y�=?���'���[$/����=��N��R*������i`�q�F'�#�@Q�m�*"�$/	R�<�XR,����HDW�'a�m;xG��M�Y���N�2@�7-2���)l����B�<'���r�����؆4�����i�	_Y!r��X�F<J�O93����nƣ�e��͘��̡�>"� x�fak���hl!�Bq�L
�̢F����S�sOf�Vj&��%�֚ G�;M�Ŋ��7��>����2�C�fս1��$a�fj�[�O{�v9S*#���X3DV";�pY�f���<���s\�m}^!�ȽFN"Bc�W���'V;f�$���m��12-;K�J*�yY�}(�i�r����Ne�o\U���W�p�ᘺ$�� �x� �P*���
)�=��x?����>� ƍ��CUT`���ԳV"�X�E��H%�����}N�.S>E��X6�sF�x�y}c�Hz�(ߟ�a�58 ��0<pSK��>v4�^S��m��i�Y�~�x�T>+����#�n��S! ���>�/
LU����v dl`�z@��������\ϟ�K��M�3�n��`�ʱk+oU�C��;��>�@H�p��M�J!�>Z642+�DةR.6�2�v�wմ�:W��Du��CPj�'�����9�r�I��[� ���;Ɏ.��,����߲�J�X���Y+�*�a�\�DŸ�5�������)�bR烹&�_|<d��e������^되sm�U�q7y�Ǭ��g�*�<Qf'�g�� k�3dC��ŭ�b��� �-Z���v��X2Q�#a�ר���SW�[�����	�?��LqdF^6-l�om�@_C�/�. oU�Y@��):.�·x������6�m�j{S�k�$Q"lWc
��_IeD�ps��zѡ�1�$(+7���+�QO����Ȭ�n��ST�]���#���ڜ�e)W����fB�{�,�ʖ���r!Ơ\#����[��Prbnm_t��9q=1�J�ډ�P ���ֶ�m��2�<;~��T��k&�㐕�YpV�8Sa���W�P��T��4q$t��e�Q!����§�g�y��\�d	�΁/��f[�K��I�������9���Yl?}%ha0�D�P�M?��O�1A����q!mD��*^���˓�Pys}f��uV7�qb��3�S�w�"@u��꟰�M�ٝ|]�Q�O̧k�CL
�ZѮ黧��Q;QxC��D97�;��pPR�lr���M�Q�~�R&n���0W�2��O*��?PQp� ׋�$<�Y)Nx\�;�*i5��5b�fö�\�>���% ����h��ի}�?zb�J���2*���j飣�){�w�Y���agEes;��O�ؐ�A�����E��*./5�!1&���A��Y2�:���2Z�-"�B�jmE,4@zֲ�[��nuH�[p�i��8�����[k�Q�N�T���W⚭�|sjr@����O������a3L[�"����^��]ѻ6]�f��A�6=�q��'��g[��?��Y!�-��������m|���m��QYP�*�R_��"���j��ܒB����5�Z�r���Q����+��or�q�}a��_�/�NN�˞1)sRXe"�����)r���&O��ӳ0��Y'Φ�8�<��=�y~���R�)�5�j{z��Y>��'��vB)���P�5E��@l)TE��b�.$p��/��7r,a�|���zry:hz�j����m7oJ��h�i������`9�ww7�;RN~�0�m��;Zk?�n'S�Nc����'t�j����yR����vj�`R��Qc�%��7H4Z�&d��y���sc0��Y���7F���s"�ALk�֘�ax��m�k��O��v(�M��4�Mm~��"�L��AP�5��@�Kc�4�vc�P?�J ����{��^z�� (�}��q���%U=�����o[_����.�����lty,1�4?����d:�,��R끡��^>B���r�'�;��h"R_�q�L,z9#�Yְ�V֨]�\2N�hӠ���7&o�Q؜�Y�^�XT�ϼe�'U��J7m�h�r1�?Ϳ��;W�Xz��Q�IX��QW)�[��EdM�y�Z�U3Ub\�5��3�b�qX��9D��wWn�C�7�����N$q����j K5�ղ�s �7�?Ҵ����á�������G�K�*��dW��d!�}�������ˀg����m0�,�-��ݙN��)o�S(g��Y�o�n}N�C|o1z)�-��/Ĥ��As���$K:����|]����*d`�s�d�[���3-�$X�c��?���~��2-�����������m��������a�cFzC�d��nHPBC���g^�{��a�o��V��a�<�iMǠ��ȊaT�O�={bf���dy�N/J���o����|V���YN���ˤ{No��hNm�f���~�_��ĉ4Z���z��f�����u��ɪ�w"��T�UJ�V��rW+&���K����-��)$��x� �X��4yB��vB������7ݥϾM����s �.)��t���e(�1�p#�!�s`�L�c�[v� 5g�Sf$�B�ȳ�g���K�3$����F|�7��-�hh؇$k+�VU�nG� $w��l�[��SK���[��҈�<b&l���[�y�!.�4"� �ǫJ�@}��>�%��o���w_�ޮ����l?��P�|��~ѯ�$�~њZl�$V�36i=�B}�������O�_��Sĳ ح�m�����L��kD�l0S��<�"�>
x��A�sgr�.������G�Wǃ*1��jC>��	X��cG�־4R�q��4�]H��l"Y��8�#�t�r�|�{�zw�ؙr����-�P���jS`ĝ&�f�=�L%�-P����z6r���}��6�6tm����ZL��+�G'�~`��Y�s�x�e��r��<͍7�t22�kz����Ѫ{%7]ݨ�Φ�?�＜���m����q=�vb���T J��Z
��a�R'_��+�a{뜞�u�
�@�]�G��Yx�v���ÂO��H�Jp�t+2�n@��Ӿ����3�s�ʙE��B�n�$wF�Tos��>[��koLFo�)�5eb���5�Fm�)���Uَi�����@�%9��h��0F������q�W�jK�q��Y��#z�W~�1f������ZB�a�~{�P��M|3�R�9�
s7;��y��02F�5�0|*>��(��>[�g�V���kĸu|;�����6,�$'�t��0H���BbیFN!y�3B�1C[N)��%�*���ߍ��fh����m�?sz���ID��-��1��~���1,�]]0��j�e�y����<����U�䱶"�,XB��e���p2�������%��qg��/c�Jl�j@���K#��|���TV5}��N�`" u���HN��/�_e�C[f�&Ŋ���&"�8�P]C�r��'%�;9B�;�.����i{���^�-���-��@��Öπ��@���V"xѬ^������6�/�^���VM�iS&T���TdЌ2�k�tSM4�S�j�[�Ө*]O�LF!�32�IԂ�)^��7��'�_�=��U��X	U���zr�x0��rm�"���ҿs��eOF;j6�.�&ߘoj�>���	��S�V��o��?����}e6��y�Qݺ�kkꍡ��j���cO��%v>�}�ο6-A����h�|�|��%q���t�v�"��4�ߗ�i���?��-��(m�F=r��Տ�˒Mc��ts�M�hq1(�s�%Mʠ�J�����w-���̘s^�f�8�a�b�����1A?����b�k�T1���r������"Lm�o܁d*DK}�^�����ʜy'�/�M�F��~���Y�eK/��Vth��80�< F���W��G��X��F�E�X��"�z_͙;��˵> ��<�� ,H(:�z�=+S�{[�Qw�,��;��!0����Y�����aW�ȌPp��6���A�-������4޲�o�.�Qn�>d)�u��̉R�i����X�3'�C������Z����O�1=|��{�n�'�o�&�JT�1R�����5n��a)o�����9��M-�cB�Mi�ĺ�)֝�D��0�(D�6��Q����npӮiu�a�mf@A��D!���,,��:N>Q�l9�����70�	ǈX(�j�&�a�f�]��>D�w��������Y�;�X��	Xpy�wW���]���k�^�y�y�s�*�^���|��N�T��/���U���<d�}> 􂉗�Ҍǆ=W��R��6P_�^ΐ���G�̙/�;o�l�@�B��kuL}���V�������mW3<�x�SSR�������D�[f�h���_��sGSƾ�-���꫌�F��.c9�>ƍ���Y|ƕb�X�'�Ñ��zo�\��4��~!�7秴8�uj����>��:�Aݱ�P�&���r:d�t���~�3 ��ċ9�n�O�q�����6��y_e�2
�,�j�r��a�����ћ���, A����5�/�h� 1m�Z��h��W��a���
��Ah��Co/�6XYq;�Յu�����no���+.-)7����rL��><�o��c�X���[���('/�
%��ܢ��-m^�P�H�V|TϹ��͡~%�W�&��_M�ŝ�%F�y�-&ad/T��3��4YK�&��eݢrI��j(��;��������&�޳��E>P�v��}�|5#6��F�4h~F��ѳ,4�'"��{���j�?3f�?d��3 |��ż^]1%�5��kJ�;ŹK�N��WCM�D�*�s_�㤋0��D_����\�e�����1焚�#�<q���*�ה4��c
�p�ibs�|[m)���)^�E׆!��@�)(�]�g�F,���n��T��,���<�M.a���O��� V3�!p�
�����}����nB/�d�!t�qb���!���g0%4���/֔m+-����Z΀G�W���O�cj��a���ۗw�|�-�k����L�,�DzS!��;ޥ�Ԝ�XZ�r��&���x����Ku*0�\x����pA;ʉ򅮤�|��6f�ͅw�Z�r�����1 �\(
���-��o#��4���l���DF����<�W����x����/������s�3^���}̻TÆ��"���;a��g�	�n�S��JWaT�~������||k(9"򤞞�LJL_�R�똘��*8y�_էP���`� A7uy1E��:�;��c���h"���YӞi�y�o��dj *��!��<����(Y �Y��C�Q��zb"�NF�@���^{�A���G���i(w�'+)y��~5�Ҁ��D��jx�9m�b�A}�Ca��u�3���*���#���j-�F��(*f!�� �]7�9p�
���&��ۗO�Bd� "��������t�V>C�>܏�`ۺ��:eNDi'�7����x�f�Ĝ[� Cg�lP��N����-�n�Z�����y���P�w@ ⵜf������F�{것��g����鍻�nq��$<� �b�*�{��"���G��!�?Ϛ��I'�&(kݘe k`Vm�;�r�1H���5���‱�^�����C��Bc8��9��W��ط|�HPbeAe�u웟n�n!6�t�t�!�rs�ai6f�f�����7w����JՒ�����a�	5<3%$����`��b�=V�'��9�),bNdWC�MaSPU�r�.�Q$��w,���N����,�v�E��g._�F{:e���g����ˑ�|�A5`�C��V��p�mgte��<�}}�]�\ӏ�N$���J
~��|���1�^��0tݴ���u��WsO��Z�X�ԙW{^�|T��K_�k:�8��"l4�o�'eW,؝JA�I�O9�,�L�	>��hр(��Z��������}��Z�X�w���3?j���&�X?�G��7��t@շɛ�.���̟��d��e��GY�;��-K��r�(W[���g�m�,��}oکz��+J�Qʁ���<ޮ���G�}u�k�Ohw�\��5��",1{\���U�����=�#�d��1&�288x�QXR����L�㓝o>�/8�<��T��	Ry�%)'�/\U���\��$�f�p�8�9���;�s���?ѯj����&����Y:W>��E�>�d.�A��rM��d�ȯ�#���ev�(�PU4�;_�f��\*��A��7��<�������'��ó0m��auo])FR[nc��铪�ڥ�,q'������mA����I�3�m�\ۧ�����~k%ۂ��a���L�꒽���$;���3q��1��(�,�~&���d*�?!Ŝi����`�c��)�q���"3�΁j����8��W��
�i,��`<�Et�y>�c����ή�2�k�{y���+�gm�̟�T�E�ͼz�cH7~�0�L�HA�^��;Ef>�t9_���$�$o���WF�2���m�2��f|&�UY^�
P���}����e�g�U�6�
���&�WU�f�d��'�nb/%=)`�?��e�?E|��oc�{�4�5��
�^<��rK���i"�@b^����/�ۃI�PYI�ZU���{t�>�o[L]l��k�����O��hr�����V�}���� ���s汳���{^�Ģ�����~k�]�M[���:����4I�q��<�<����K$CjlJ?5xA�.��׏����v�}�)���v8t�W½�|�[�+�]�6a�%�a�:�@aq��u��YB_�b��evRR��ݍ�����71S��mk1�x MiO�a$�<��7�1���m,`X�'Um5��,�0ݼ�����<\�cM��DC�?�2�U1���� D�]��N]��9~��ǅ�u����R�j&0�MC!$K.�A�#�ׯ�	������ދ�PCDJC�A�Q�}��9������W��)��/V�I������Q�!e�Bh�Aƒt�m\�*4�Y5ۤ����Nj�Xd)�<���UG4Q��=�l�*����uQ��U��M1)��03� �\����-s�i�W2�s����¹�o�~���2T���ϛ����ȍ�-��ʓ���wo!-�tϯ7{��yr����̅�(��$���&��d�і�ͭ�|���瀙ݮӺw���u�^*P�Q�m�"�G��k���>9��1H�_��?(���8�Jz�
�6�z��3�Y�^J�*iz9c�ՍEV��/��9!���S]l��0hy�6SFYx��;���kL@���4��8O�6�W����v����V\{@�Vp���������Aϳ���W��m}�g�$���lj>����y"��|�}��ӄ�o���D3��|yjri�N����:��r�T�R��ڮs5���RQ*k4�]�Hk�AOy���M5�kF��ˤz��/��0[3�M���
����Y|�JB�3ں&��kmS���m��S6^w�`e�3 �cqF�_�L73�[iG�5;Yt�f8�%n�������:3Z2#�G,D1T,b�9�fZ�5z�x�jm)4&�tq�^B!�O�U2f��R��} VW�@MAM�GO��zr�ݧSv��>�l�`���0!��C{].�*{Ҽ4��ҷ.�����S~/�S�j)���iR��V�m)������+�q��!�_�𨥐�y�+�� �G J 1%��{���2%������)������U�����ܮ��{����}����ٰ�FC�q�5��*�)�Ts�8~�BF�|+�WBL��$u (~{D�)Vݾ�e��4̻8FL �G��:$��W����p=��X_1"�n OM��ȩ�Qf�w�2汼S�2~Vj��<�\z��h���kBxu:#|`N%�:+¸�$����Z�y��J�`�,���5�@�S�O
ݮ�~��8{�����~���խ���ֱ0�sc�4��Ȱ�_Q���)�T�Sr&�>�"�O"�o�Խ�^l̫��T�#���l���8�͹�mL��Mg�oU9�˸� �@"�p눯_�
�=[n6��7��,�čo5�#^�Fl��d���"���z����°!l���q�Gёu�0�u�������/��S2�r���ǘwl��/�E��(���4,f���F6�����H���M�噤|��#r���_�F��]t�[uv<gX�m���f�H<��Q�IR�������T�Ё�?�8��+�+C��~>��8�|�����R�u�t�es5���%�͠4�xr/[+��I�K�{�ϿϸX|��3͂��Na�_@��N_U-�_�vAS�w����"�:믔b����d[ӗ��n�#�XX0�t'��K�����1�,*��\��6j�؞���Q~�(8^ad���0��`~O �� >�5�4���vn�X]{B%4Pv�R1�Ӿ4���/����X��� ~���T�vۭ6�bZD ���H���|��(�R%���̮k�b�u��%,��D['>G�Gb�1�����*K�Me�,�z/&K�Q��ى�S�LqZU��N�-G�٨\fr�Z�3ݱE<V!&Hw�*�i"�������C���������Ub&ZJ"�������&����F4f�����C��S��P��䀯hu��R�/ym�E�Mz��=Y:�����vK��ܫ\%����m˸�����q	�	3Y�kˇa���:���4#�4\��R=Uif��:�<88�u3���V�:u�kZ��:D�Z���m�+=A3�i�]�+��z��L�;{I���1�Z�|+�o�����Xb"��o�o�x!_URΩ�ʎ�L�dc$���p)��|��X�ꐬfKHd��t�9A#�I��L��g�ڷ��R����o�a���q�;C/���%�TH�'�͗F/
�h�YA�`QRX���V��Q�$~iNiM�UiCk�$k؆�n2۰�ϐ;��IX�6w��9"�F���� #*�W���7SM�1^h�wMq��q�$&|?�M5K���ϛ]��h���߭�����rQ?\���rut�x�ZP΢�I��Dt�v^@<O@Ў�����1@�2wm�?������DBĨ�6��[�Gc�J�&V��{�li%��fl�"f��E�j��j�.�m���|x�����9�u����&���ǵ�`����&�*��x7Ǧ�T��"�s@V�\�^�e�̊)�m���4��M !��i),E0ܪ�rJ�c6r�z�,�Y&傕6�bXz�������y�>�sz�w����zV ��-&KS*˘F�*��b�!8���?��卨AEi:�|��H�'�+V45�g���TJ*l��»M���kn~�b&�3|<� ��Y������|�Pp|��v���[w�B ��r:��OG����L�M�V~s���pu�7��u��
I��K�F�V���ۤD��K��Y	�����KA� n[��EH߶���+cԼH�V��g��X�j{�o)���gc�;�W�����~Q&��t�zYr��E; �:�,2���CݬC]>�]&�ҳ�w �Q�F ���I���ǘ�!�m���2�K�)|����D���
�"�>��/��%��W鐅<fpt��nk>��@`��
@�����ZD6�K��/���Lb���6�p�W�%����_v��x�8�q%X�N��Ò���V%�t);�W���y:�O�l�E�1����XhY%_�)��.T��>9����i����b69Kk4݀��ɆKQ
0���Βᖯ��$lc+9g�~U����R�����ckZ̄ϩ�$�����i�9�@���Q�Wa���3�9�#����3gs�B�93����⯀gJbZ@��4�gd�	�q������1��M�P[�ɪ@D���:�i(/��wR������W�
�ؑR��y6���T�
�ѝ�� !!��:b�@����D�1�d��cC�%��^F�EP����K�_�r7*b�Q�������i0;�[z����/���W�������'~��+�5ԑ���oM"�B����X���OK��䦭Ř1t���(��ϥ w�kZT[��[5���;{���p1Qr����A����6������YyX~g{B&��/%�m��즽�i31�V큉�r�Lv��]�h@�`����|������@\i����"��WM����|�h$m��f=��-1w��"a���`8��l�ѭ��MB�kY>��<�YEBH��4ES�O�V��]�&=�햐�"_#�J�Yۖ9Tꏀ��3�酸�=W�s�n/Y"�*&Z�W�qW.6���7U���?�T(pl�l�p�~���[ �F�L��D4�~��=���O$������父y?��g��߿yy\����R�;�Վ�}������yT9?��OQ/��ܸ%�΅����l�+�ܻGa+P�"���oj(r�[F��oV�:��=�����\�������]�Rt��^!ï�1P$�#�N�����C�c��Be+�2U��v��v4�6y�1^�MU<����W ��p�n8���zƱ�Yi,,MK������O]�V���	t)I�.MR�/YYpY��||t���%7�J�6�������_�u�*#�����(j|�0K���g*T�[��`#��\�D��_��N��	�\�Q�f��B� ��O��zr���5����ڔڲG��5�7�yݡ�sT�m�P+|m����]��_c-^/e�Uԋ 6LZ��;Wg��tup4)ɏ+!�@bk3T���t�9������q�;O�e~oo%L�{�ƍ�ap�?=O�T�(�*�;��~Abu9�YV�Sځ#�-5�r6.����B�t��y6!�ë�3��8i�]όڔuO��<cUm
���N�کs��5��Nb��3�AG����ӭ�u(=��9�	�����X(�t�el4��1�V�Id�]�(��[�A]�V*���L���5�k�������%QO�r8F����2+�8��};�| �N�kzS�*�8\8�m^=f!�3 �r��� ]�SHKϡq�ukɹ�?:J�S��� ���,J���q��`%�Y���ړ���d*A&�_�K/��Htiz������k$fj	��L�tEQ��=�9�Z��3������n<6Cc�?lV�)?�V��ѵe���/��96ƚId�(o���BI�xr
U�v�+��'�~��wA��j�K��n�L����
��S\/C����0Vp�������>͙Cx�E&�SX��<Z�<a2��� �YV�1U�b~�	��XBՂhGK�FsQTk�P7�jU�W��&��W���d��N*�PU��&�KM��8�w�1UM-� �G�^�w��7���c�ug�'�2�&m]&$��Oʇ�_fĮ��FRI�f ��(�l��!A1���������'pe���ܖ�ŀ�Բ�5��g��ѽ�zo=�r8�-�k#�R�@�
��x�j�|b����pSݕ��'%�T3��~5��$Ӏ�����Ņ}Tc�����E)w7��|�{NX��ב��E��)#�J����w���?="�� ��Y>��{�/�'�԰4�&u~�3�Sk���o�v�ȓ����r���d�.�)-.ap�l�壖�z��l�!���r���
�
��r+Ҷ3P �:�w�c����$BD=8��{�K���Y�����Cb8�&G'�yi礡 �\�3H;��$�&G��갥����Ҙ�p.V�	�atЦ)�O�~kU�D`3�p�BP]gӏ~�KҬamL����`���*9�L�9���)�U��q��8�Hq&��x�J�Z3�g��N���$�]{7ŝW0�����,o�k	�me�R��O=�-_�H��
�"w Q��������6��\6���W�C�:�evFV��돩�*a��9ۿ36��f�<߼x����8���!������=�k4%ڸ�9���Yl�U�@�h`SC~��������Z9V��XAz�]����M�>�s��,����EX�=���ȭ�!*�W�h|Xbۢ_�*���n�bJZ�෢��WQ8dx B�5�j,$o�x�ܟ1ߓ�p9�Ң6DA�mO�~���^��'��fV���\���.\��]��fڢ8��n'���Ήҳ�"���4⭤+'��=�U�:U.KC��A90z�͖���ѯ{&�������C�f�7��<3x�̀ڀû�N\��<Ф���[bz ��ޯ���^����@ �p �!�$s���:�'�x����?�?����$�@�l-��(��-�a�3Vm=Xi�J�r	���������D�vN�|��Rä��K�� k.-�g�!ֿ�h����~�-Դ�g햌2�П��/�9�>�k% `=�����Q�Zk4�f\�������U+���g�a���}n���C��xtzҠ��O�͜/�`�Jʹ�l
QE)�5�` 8�����-�� (hmHڶ
:�H�sڂ���<+�3۷����Z����ٽ�[R[i�����{``tv![Ԏ�d*�S���/�І��ɂ��E�2}G�����}��!�3�O�\�}��^��ə_Z4�_nS��B��~��Z�r�GF4���)b�����?(�+s5O�X�ˑ)�
�q��*�!c�ֱ�>=l�+�ԣ	�v�~�b�����^A���>�*��x��'�^m�,L��YQKW��� �r�"x��ҨW�ȞJ����� ����5HG��{�N{.�����1��������z�=��H:�����Xrي�(�?8��8m��������R�!���'�^��Q��"Aa�̆z��H���h��d[�ĉGIǂ*�o�4��-_�T�&���={Sd��ci�xV�p]�ײYcG�.3�b�f���3���տ�{')������WU�rKd�f�J)@ �������ɰ���Gb������H�oRkʕ���i��*m����#X�|�<8K�7��Z��d�~7������;9)�����0��$C31Ϡ�q Ҹ嘮����oL��Z��q�\p���>&�2�G��i���uDq�0�-�h�3�T֞Ҭ�`d`A��ppf>&��@����ܢ���w��l��
;��&�5{D9��L�/߯�2@��!VR�`�3P�Ԗ5w��O�&�P�W�y?("Vq����6|wOUk��4 "ez�*���V�s��
�`iՑ��*X#��EǅH4B@4 �{��
�z[_4&?�
=T�8Ѱ��{LC(o���a�Ǘ�u��U.���1�dN �Oq��L������Jؚ3f咨G! �u��f�Լ>�x�y*�w9���^���z�#��}EQ��2�[���,/��S��v�%s���IX���L�}2�"���+JB�D ��k����#<ou�jBƇ�M��$�o/Ke�qI_��Ķ�N��[�M4�=�1��P��T7'�3lpr�+K��F)W���^��ٽ?l%�]�|����Ə��Ց�tu�{�jȃ��wS.A·�[�����-� hDA8�ҳPp�yǴ����0%;F��D'�rwq�"D���P�Kq�)/+"!aQ|ꗐ�2�v�M
��bxW�B���G%�����x��&r���}��WA�и�g�)7��/���yl���V#�눛g��ǭ�=d����uj��ڨ���L��H]�Bʫj���s���K�2�~d� :�3�S��������7Ȟ�!���ϒ�D�%�]&J��j�淘b��閑QInIK�|R`���9�Y�S>٘�����R�q�#ñ�T3���I�iat=�<��W�߫�d�%�YW��ܫ������ϛ�T3�mn�k��ٶ��g��Ԏ�j|�(bO�)�4ޯ=Ӹpo�sa7��0�k��ea��n��9����y�U������Z�vB޶L��˴�zw�į��#V�{����@Z�,��8�����2Q���}�#u��6�$fi]���Ǐ�G�����Ȃ�.S d����#��ԯlξ�e�F@��a�q}���w �ǌ��v6��#��#>���D����v�B���֑Ӄ�N��?�(��h��I��Wӧ���x�u�i��i�e+�-��E���
��Hnǡ��}D��2����6���Cb�>Қ.j
ػ&]�����dͶG�n\��/��U����rc�"�2��e�<!v5���lڟ��S軣:f=[?0m��ok��})�+S���6�~�A�q(�Z��׹�%^��(Ej��k#�l-=�"������|>V�I�NSPؔ-��,W\��0��K'e8���4)��p/ �A��T4��+I��-e�8 ���/ܿ_�/o��xx�7���h�s��j��yp�bJ�4k��0#�6�t�л65	�f������pX�d�CC�l���TX����������2D��KB�o�U��"���j�+�*߄
g�7&�~��Ѐ'��(F t�^���/s�j���>|�,TO�/��o�,��Y����B�+��`�Ve�mz�=���r�جG+x�'���g��UU��}����S�B3dx��ve�\N��V5�7��8���,1�fWl���<��d��'�"���;5�S�H0�C\8�q��Q�YT�������s!v��{�z�u�kB�V
�����PBv����5��&<oY<�/ۉ$�ͬ����b�	���\���s��k��wiV�w�ʒ'�Ŀ�iy�ȣ�ު��A����ѿ�&t�պ���>��������Ō*��:D�ׯ��������R��o�0�}2��'�.m.ׁ��ܿ��Yc��}��I����|���!i��_[���;�w���>�]��	'��~p::	�k�,���OI	Ab���&GN����7�*��a�O
� >����wb*��T'���m���Qb
�jQƫ5^|�V�����	ݲ/�|��[�ى��	>�Tƞ����r{��?L����k�Wru���>)�0��_-#��=��%?���S�}��1O"d�rSy�>H�a͚�����p�67ɾrg�a"}�M��0�:��A׊:J�~A|�hY3��PA��Pu�(�i����vwo��Ѝa��B�"�� �7Ld��]��o���i�!��[X7AQX����t�þ����������q�)���m�VҊ?)�;p�4�*N.(S����0
�$T:�Q�R�@�P�W)8vX����l~�inX�N��M��W=�>�������{�J�s��*�f���X��C��&�QŢH���^�䑂��� (���I ���XUWBT���f�/�i�둜L3� m{�qs-�oة�5[B���
��G��� �5��S���a7�D3�l��%-��K��TDx���s�^*g�,��� ���y i��l~k�j���dL���޾�0���i�-ս8��g���#�+i�-��3(�&92R-�j����4+k3��Uf���du2|�	�t�_�Rm�ϋ�����,u�N��*N�谢���q!%'C��:I��>h���oPH�4�K��B\�b����[�Ë�,5�|&ܘnB���,<�i��;��~�:��!����Z�5Ş5���������ܙ�բ�p�1Q�۷<��}�ÃY��a�ZQT�$�ٵЧ��P!��X���y�6��;,� ĵg�8��G�)\��'(,�������5��?h
tH3�OY�A�^�1*�[x�
����x�tz�B�ȍvQ@�ZN�,�����3�䕜�)��M���%ۦ<��/X�kQ��x��/+4��+����̅2�|\�K;���d>n�n�!?�r(q��R�!�}��.��������C1�߅���P�����ŵ�1XGl�&@߀>�a���8��#x
h3M-�q�U{:"3����u��OI���x;�ٔ��t������Znfכ6hm*#��|��&z��������@�/��:0"[qw_��r�{�/�Pϓ ��E.L�A���ȧn?�߂މhi)ݸ9�0���%����;5ɦt����[����"��!��ZCY��� ;9���p�ĺ�K�=�oR�X�p���^)�z�������LsЀ�]|S�c,2�ALY�	��\! {>=�܅&�Χ�n���/J�!(�^���Oh��^�ztcm-�n\?��TT�m梈�NoҞO?eد�5��_�2h#s�����;�Yͧ��ۥD�����߻�E�i��U'���X�'����恱���b���<����̾m9�V����ՕK���g��3�B}��T�y
_Eb�6*��Jc��)�W�_J�nپ&�P4���(�F��w��ABTC�¶�f�+�?�-�&��3�4K�=�����}[�:�C�H�h�K}s��l���D��Jk±qV�:��.���V�X�����&FN?{�!�QL�A;�yƓ(���u�յ ��p��[G���0��0.�~�sMx�YcSq��3�:1 o� 4��ĥ@
Fѹ�����-���H�5T{����.�\�U����bo`��7Z�Q����R�Ϗ"_��E5�����0V�ܸ���ڢ�ʎ�|�������2�*�Y0�e<$8�r��E��5�C�pLdD����tz���!=�ؾs���gN�^]�
��F�3��Lp�U����ǦDA{�/a��$J`zR��b�?��ѵ�F ��fp��U�	z��A �U���U7�ӗA0�sX6)�}Kh
1x���g�#��e�[Ô����A�ZU�Q�<xw����O��X&-�F	����h8�k5�~n���2�]�&�8T��+������Ձ��&�Y� 9g�^��W'[��{u�v��^B7�MY+� �;j1����A���O�ݣ�RK ���d�BL�������]Z��&+�i|��������\��rD��62O�\����"/q2��E���Oܩ�)��|����6�o��~���\�&E~����S��m<?�'e�\Ǘ�����?%vW�����AaiR0�rܷ��}	����D mY�W��[Y�t�ёܐF#P2~���~j&K������j2��[x�F�է��� 5�����"�˽o�n�'�L�~��\S�"G*��d���;�V���iw9QC�]�6]�����wg��w�셃��ؔp�Aھ�W�
u���r&7� :���ƔQKXC��x�}������{ؾ��CW��g��<�i������Nv���W�/���1(fz*���9��8�sez�؞��G��D���]��j�e'�f�r_9���X~\mG�V5�p�	VĐ<C������K���J�aU�9�T�B�<�֭�*�������5��EJѓ�eW�� B��o�*6��7�#a��9%$�xa�'��vW�^�ħ��@%��D�S9W�I!"�����Tm`NE�uʻ{!�֤��:T�����H((ƺx�.��b��4ƁD`k����֨�
���K�O>���"M'�w�� �܊)�� ������P��}�D��s+����o�����U@e6~�֕��c�kRٽ$xz�c�}ò�w��1��Ӥ�Q�Q+�}��M�d�j��Ȱk����6ꚺ��"O�3#��Y]�|4�,ޓ�}�
��PG���$���W�"~���3fr e�^��H�N��r���k�z�{j��EI��Z���fhLvZw�ҧb@�"��p��}�;��ZS�mwC�z�Kh�pE`��P�"�e���S�A����0y���h�;�׊���M�"sl�EWH4���i|�tu�G�}J��.$-�t
m9�C͵�	�##�x�c3��_t�}L)�jM�d[;�ݞ�Ld��g×���'��Y�5ȑf��4�@�o�^�XD�UA@@�=�D;e0�0�^�t��� �l<��B�% ��=tp��s�(�\s�Gk��+���>�������Y�[�%R[�?"��o����!#�*�)l`��p�-���1:�a�������Zr�Rւ�m��rQ�^u�i+�ryJ%"��v��~��'�<��Z͔(�5��z�,9�p��rX������Mg��2:�VUR�`�5��%�5��~je����������i}�*n����nn���ǵ����1!�x�]��������7�dNj~$�$M�՜*d�����L��Pqu�=�|X0��4V\�<[��Q�P�J?�'��|$G>'�wO{�$�\*T�#0D�c����_�V~�J��2��u���c9�V�!�L1 N.�H/�ׄ:8^�u8(���H;,��D�_tJ~�%���$Е0���L�
���<h
x0$V5�B�S��L�R�Q�>��F9��U�_�3O�E�	�6�q���
G	�\��$�������:e�sr�����l���Qy�̏֣�ach'x�1��*���ݥ��Q�y�i�ZJ�e�;�`Ƽ6!�0�}��Æ��WԎ?0�7��t��WR.��ۇ�	�\y �S�.���yn�m]td� 9]f�n��4O�2<���vD�ώ�����~ŗQQh�C����K�L�K|�7�����X��4���5�_��-=�q�_������z2�ğ/:�'�7��Y{V$��uF)}���*�+0�%>��ZR0\�,g��ǫ�+�鶯��������b~qF�Сh�^��w�c`�A�[����3a�+��4��)kt9�����%�_:�R\t�?�j���]Y��m��������FOV�5"�m�������!�`�(17Z�Kc����P�unX�b��|�9�H�ү*X��aE�ǂ?3���,��/,+f6����������{U�
�*Ă��_O�6��Z�X��I���t���hz��0��.X?�iw������os�W_�Z��u�,�
vcQzX�����Fl�0|4�_� ���gݓ(�r
(/�h~��%�K�&�;��ɋ��1i7�]��XS~f�M�	=�?\��M������^�0����w?��I;�?�� �,�|l�gm����mDќĒ�������^�9���D�~�2=��mUy����7�Ȗ�tv��{<���f�GUUG���haOo?m��P\���D$�/�޴6���L ���O�'G��W�{�ָ�r��3a�����/�����7�V9��<�]9o_����7whDF6�op�\�ο^�q�BrΪ�h�G/��>������m����1b�E��|�K>����Z�� [홮|���n
�Z�E�|E�Tz�s�qʓ�{�)�$��Xa�����H=�j��S� ֈ2ٜ�B1�&@���Oy�籖F4"R	�(K�H?����X��#����[�K�i���jR�ۃ� /��ʖri�0SE��:���~eF��m�`|�{,ӛ_RO��Q&|��R^x��}p���գ���t7��[Ƿa}յ}��<���@�����eԆ�ܓ3�A+��=�K�Ù?幙(��S�n.�j�;��|q�Ći���<�I�C�1�J��^=r{JY�����T6�c�{i��	��4W�`#�q�xSH��+
�`�pМY�9���+�ya�k��������ߴ�|V��
y[H�i�3FV��>h�"��� �VbM��ۨ��i���ɂ3#2&��3J�	u�"s��&�9�D���+���#�<�=��v���
��l�h_�������u�d=^`<U��FK6,�1Yr� �X��������f�pccFf�eh9�t\NT�g%1���b��	�p�N��G7vB�h���Vz-D�:�����q듧1�W��M�tU3g��C�^ V�9d�S��E���͇S�΅ễ�6"�>w��'���BUp��:UU�H&ӓ�xӜ�E��ڳ�t)�����i�i���%vK�A&Do�fo�J��9����]�*Q���~����	�-�L�Z�@Q�r�ə]�J��5�%D�\L������,}����lqv���
	=� �!Բ�[�����d����� ����,q�Gϼ�V��3��Ph��7	+��߾��q&f$�D�˻b+<�2lu�9G�=�偲@�L��z�X�c�Q���\�j��� nj����|b�{��^�z�w&����?E��
��#���Z,��bqcK:�u	ݸ����r�<��S��X!Jߴ#?Η��$E�V�d̩�=@f��Z}{C��y�Q�Ʈ��>H@1n�'��)q��D��DW��>��]�.@�$'RTK�|�1Wt����_��������ݢا*���V�����_.Ȅ�eD�����_U��/��\Y�s���ߺ�=���h��l���Ȩ�L���*�^k_�G�j��/��m���NH}����B�Z���t�)�n2[�g��:�g������!S4��ޕ�6���G7�Չ>T�n(��:cS˯y��gr]{�Kx�+�^؝]_�b�+��5���u�����+5��ˑ
r�g��(�f�{|]�F��e�g<�'Y{�U8�ŷ2���dfv��73q�W����K&�Lf�P�|�.����i�ܶUtE�/��x�{aM,:�%ј������B1
�뱳e����{�6�'ESg7r�0�D�to`�V�ƻ�ty���8�
l��/Y9s�m�*`��cLw(��������CT?��ѪQ/j���|��;Q�d/>�kk ��H��9�l�B���0�-��z5)�(��@�u1�E#o�_�,�գШֹT%����*�]��:���M��>�ҿ�{9��^5<�5��Y2x����5�E]�����|���������*K\K������Wgs�0%4M���������4,��g�-��NwK[������� 6T�?�.t߭��#��x�~Bמ�r,q=�Ϩ���8��Tj�\?�<La78�$��B�Ld~"?ui����m;Q�'�"X�xk�X!�yoE�ܢ�=��݄B?k�AK-⽨�U�������7��lw"��P����%H����p�X����>����F,}�8d�r�X�p�9?>R�,�#!1ơ����r(&�>���aoS���^�k���:Bد!�V�Ί�!/9�K�8�CR�.�*Pƴ�AY�Kw�=y0�h�i��=<��^>���9�xm)%�ύ'���{��u�И��(Uh��u�_���5�~���]w�a�l��g���Y���i�{�^����|���J���X�հ�ûɌ
��A"^����prp"�8K�A�	"`%���S��ʫ����@�?�{Kc��AC{ԏo���0�DI��&�Q�Ұ҉��i8wҸЇD�L�.��L8��m�J��P��0���71B��3��Sen�V]�}ھ������t��!A0�TzE3��]BՍ0�	��搢&鼬�I�v����!\Y%�Z�8�#P�0�~� ����C�d6"�h�,�-YA_"�����3^	��d����2�yx����)J{5�ugM�5��&�˦�����aX��`�����5�e�꽲�pW��e��*���.m\53��9���>t�O`N?��A6)��^�)�lt���F����d��;RU<I	�1\j+�c����<m�h�X&��n��p�ŉ�� W���I���+��U��MUB,��[�|�]N��U�S���M��E�Q����U��=��M0O��`Ξ�h�La��,�^ܔ��3���[�$�E ��M�X�� N*<�0�$ߨ�5`|�ZZ�IΨ�u�h
��^y+,$6�\׎� 1ӧ��Ϛ��$Y`�*w�L�M�]�F�ć������vmH�϶)��5@Ìe�f�0�����9��Q���Ma�=g"�p������-�Xs��b��p裺�!چ	��~v��t�6�D�-,T\ゑ1�Ka�v��z1��&���������� Lo��5V"�nc���B�f��4����]�E���A�G�L��7>�e�r�s�!]�'�W�rfn�Ȩ���os��	_�`��k�������/JE�ٴ�BF�^/�&�w,��mS�k/���r�~�Tl�idg�R5_N�Rj7����\��$��q�)��͔�q�+���T��-s���7�Ou�R�L}BR��9���\؍�����yD*v'����;�����g57��vmA,�L�3D�4Un��(�c#j�̅:�NS�C�m��9�B0�2��O5r��ߥ��͒��*�@������q��(�|T���I~-��o�#��+
�����E�`E`�;嫒���!Z�B�B}�S��9��7R+�����%��k�cl�oV�_�Pj�ָ}:�p�e�ޮˬ��󢟙g�i�[1�h�
�rR2+%۸������2���X%�p��v��X�ə�좬y2���Y�ij�!��`8�n�
eP����섞�����Z����I�����Uf��K�6��܎LeJ�Q�6�oC�L�o4:��W>�]�̾[�օl��2R+�%��T�9�ڂ��X!��y5i1pU#w#ǩ F��\X1�1�2�g�(���їeCD��Ѝ���q[�P���b�tĭ�Ȧ��_�T����v*��k�7H:>��K�L�R\*n577P�)�q�9fy��9��_�H�=r�"���fe���/6�=���'@DJ�Eqh��XrgE�Uf����b�Y2zb��Y�M���qJ���%��S��^7�'���(���v�;�E_S�P��E��?nU;oe����o��v,N��AŪ�x"%j�݇Z��~#�_6�¶�x.s���2A�8S�M�	��s�������'gײ`Bx ��j
(�9���q@���}�k�k������N��U�i	����ePpZn��l�k6|v���D�'��X�U�,(=�d���SM�JX�l*զ͆����]�{����X^��q��G=u�(�|P��M�T��������$\��e���������J��o �Ld!\ ��'��}�u@	e��r��Ƣpd�ދ{�-Y4$M���}U˵�����A��|�__ˉ�q��0|�(��'���]���\%)̯>���AU�ܢ����pvO�%a^"-2ږz��Kbt ��cM��b��5�.TuP>y^?��A�u+���ݿ���L��5�~v���IeCò�����S�KA���q�������7D��v�k�P�b�]�R��~��d����(��2 �u������J,Լ�J�Pg�ҍK&P��fpooa�Q����C� ����P.M7�$��?�\ �������W����)\؎���t\����n n�%����]�$�ʿH�m�}�{�9�7��!�t����Ԋx�5Â��ƿe@֥$1���Ў�}�o5/\�{�㫪ĳ?��?�|�8�B��Ϡ+���ވ�D��m�~�_{�\zõ���V���&W�KV�dt����}^]	̬�M��0���%�k[
�V���%�p��Hc�'�;������8T�	�y��kR�;P5�� �V�r� ɬ_?|�K:|./ْZV��Hf3}��ĘT9T���<n�u`8��;�Lf�J���'G�yuG��b�� :��Y5S�B$��)�U����+�����-�8�.�9�ug!	Q��(ֹ�����ꉁ����f��C��B���5�:��'.�.�M��7H�D( ǉ��]&1����
�ڏ���	��X�j���N���(�`���CS�W:�]��|g�.y�}��8�]�|�3\�<�r�+�O+��G*�Q/��1.���.W�v��d �S���D�"�pOԶ����c��f�)sô�t�Ii���s��
��O��"��r�[�	��4�$���C�J}ɿ����N�p� @
�D���V�_i��cCK���ҕ�O^N�����ض�V���	?1`����L��X3QSsW?�C�'A�|�_G��.K\�G�J����Gm��_6J����h"m�4��~������[�&�lS;���\uT|B8�>Q�2E���n��Bʉ<� ��s��_Q2�xb�(pBf��{ǇmҤG��IU�i��l�\`����,?�kW��3S����d���+[	�:4�np���N7~� ����k�Ӏ�_��3�δ�o�Xc<�&�� ���j?̨�� e�Ds�u-��*�1�[RBiFb,��IV�c�R"2��[`��ɃB��v@[AҠ���^�BI����.�6v����l}�;��k-�gO��UJ��]Zз�46����lB�j0�U33B��!�+�zo���g�/��� ���.�A,i=1�K�(B�l��&@KP]��uj�\�MA0J��b������u�4%bw4Z�B�Y�	��״��/�3~��7�5D��X�د�}y�1�n�9kc��>g�'��sh����ԏ�k��z�=�/n�B[ν��$ E�Y�Hl���fv�ٖ����,T�"՛�Ir۹�>�����{���na07����R�ϖ��^X2�C�=�)d�X(��@̿<,<x�c�,[ꐛ�p]�s80�jQG���<{�t��PL_r�����Lh��	����$��7d�2O�h3����� z�+��B������O��2-;<�'$�a�[�����3A7��Ǣ�IP�]������@ B*?��F($t	���NSA�Qڗ��M��h�-*^�H�l=�P	L	���ni�F�T(���##a�ѓ/:p�%���St	[��3��{���"eK/?���I�Y��q��aim���{���HDv��jc��5b���
�u�]9��Ə�%�>�~��G��@�Y�4�:�u���v����F���
�%l-�J
j���m �a�.b:��F��	�\��l��i���i�yZ3Vo�2�a�%�z�zew��cOQ��B�[���{���Y�|r���r�_͈
������ߏj7QB�|�ύ�]��ٯ�sZ?8�]�L�ec�ͬ^u��h�q��n[��]��Ĵt �
���7
K)�)�/�����׈����s2����4�W܌�驴/S(���>P�T��W�όɅ���&UŎE����}�.k�p1��nI����@	�tw*\A���:%�Ƿv��YRy�����
k�R��T�g|
��4�Iץ�\ee� ��Z�\�d3���Y8��H�;]�,_�����#♒�b�ǧ�}ɰ�dK9W�X���:�knт�ߍǀ��A�&���z��a�g��{��^s{6��	��η�+Ñl[����o"�[�j�h�;��y��ݠ<��.����\�̻�o�~�w��v�x�>{կ�̦��%� H@���m�F�g{�~��k��18�f3�3�P�����ǟJ0=V4�Z��0�cj��ӠЄRazm�&1F�j�6e����[Z�C;��{��e!��ː�OOOb���Hf�B3�=v��f��|�;=n�w R����	��ȒR��!�tV�I>q��p���I^GK�D��\�p��1�]#ز��Z%&4���{�*&E�<b�4��{@k����n`
�\����|���Gy��,o��u�Ō�VJa��<�������N�X;8��"e�c2��E)���
�dՊ��]��J�t]�vM�C(˦��$��c�I��dA &Y���;�!���)��P�D��_����Y�AY�ci �RP;���
XU� ��N[c�O�e�� U�,�#��l#�)�0L���]����)��$0�Z�Pg�xS6R�+T+��)XՎ_�l��:M%��&<�)��F�o_
��M�UR�o�J�R�Ժ�� ��R�9�E.E�BK|��-�Y����'�ʲ��-��B䦂k�zy�H*}�J,SV��e�R!���SA0�Y3`��D�'�	�׈/@Fk�M t��#�P	Zq��Gئ"�S_��<��� ����]!k��L��Y9D9Zj��!4+�)T�� ����X�Lp
�鳉 ׋��#��
-�La��q��I NӱH%%X*>Z���
��j�<�S���B�c˲J����i��􅨭�@�����
@�x ���)O�/���.y%▐-!��^S�p��"(�+�Y⑥,��p%h�T�9e����,Z�m'�SM\Va��<�G^P�f��⁤�/��I�y�q,,�v�Ь]]"$� `�%��S��pBj�#״��/V_�E
��e��"��B��)��e�m'r��J)qWk��6eKA��9����,O�`%�ڈeG'+�y�� �Dl��B*)�B^�bוO�Y2|��� �,\�|.>2N�Z�ڏWG�z�8&OY�ĕ�-��^-o�.��e����p��u�:9�pHd�XvQjGP�x�iX��oɒ����OH���cG��'�!淣6�wQ���6�.��7���Ƴ:�J�lL}-C�LJ�~-B"��-�q���eL�eo����XVg�{�kl3$B�#f���>��8�!�8��:D�o)���٫���"g~��(��^DS!��O_��G�4U���Q���$�"�5Oӆ�ө�۔85�L�J�j�L�1|�!5���������f}�THYc�G!UG��41\�b 2d���şNL�̲�`�t�K)��y�@_�P���)�3䆔+l/NX�mS���ik����_���nA�
�j�ŚG6<A�i� bUN[���v�9�^*���`h\�F��,k�C��2�O�>��}�0���N��k$N��̖L�` �x��|`
U��v�3�R���qx�
�my:�P� �eW��R��KÛ�ۛ�F���x�bJ*Y��&�MX�0-	�7R� �P� �
K��f�,d"���u����l��R�ĳ��-����vw�)4�-�x�M�9XG�����I1�#f�qH�o��&����,<���N���/@���OX\�֝-o��{7���|���7C�q�9ݮ��S�{gp'{{iH��K �nQ� ]��k����RP�IA�|i6�1�3�d�_�t��
i_Ԙ X�6�V������ɾ}����T�q���QD�,�'�m���)�0�	�q�Chܲ�A� k�f��(խ�	!��]
7��S�U�'B��o�J,y���'M���l�f��6�̦�J:k��!����L@�i���8��)��Z�K*&?c��A�K���r����駬ܮ�}�>�Nq����wo,���:d▲|�T�v4�� -���EUVygW�Y�Nb�@�r�چ������{��!���S�7q���_�l֓�f�<��b��"[w�u�H�Q�X�2%��l!��b�鞩;��UN
�62A�&�v|���bK"
��!�5-/����\4A��#_������
x�^ܢvg<�!�:(�xxR�$�Gsi�0�^��S���B�������5s�x��
���D9�����J�o;�9�N�#S��.b���y熌�eHYl����<ƣ,�&��j(���F��2{����7��צ�߿�f�����yv���ӓ��F�����������SR{y����|@2��t�}Qp>����Ի\/cG^,h���v����P{Ą��f�Y�:�.Zg���E^�TS��v��Y&���t��b)��4���q�D42�ؿ���8[�I�+g��f�����f��녏ى	4�3R|4AK��Z�!ȉ�i��`"�����L^��Q�h��{oMt�S:��������6m�r� e��T��^΄��Z��+ҙ#�J�a�IA�y�&�ڦ���ǭ�0e��j`xU<�Z�$����՗ ��2R���K�P��-����,�J�I�%)��	�gp�ւF�6J-�Ym�%e�b�� �娰9�qhNID�8��#/Uww����J� ^;| 2�#B�4��8�j���K�.b��M!���xs�qXA>�n�m����l���V��.f�N_�8D�b�d�jC��f"�b^��bj�5v�F��T4�̵�<B���M
���2��%Aq`G��@V/L�8�nh.\cO�lC�m)U� $��ᛊ��ۖ��]I��3�&�JALv�b&��Hy�"e�f`��櫭�b�b���ĬPL�*H�|�ܾ�d��3L��0�J	�$��j'F(��MUH�N���@66f��G,�[�D��n)�^���&X����A|A�R�KU�l��q ���+AK�Ǳt�U��0##Ț�&�X� ox&/�2�/��a
֥l:��R5
��d�$��x1���9�C(ħ#�V��)�0���~�����7�NCV �b��3 [\�P�������N�0Fd��N
�m
RS���v��L,di� D�*�ݼ�K����fHǨ�@�q�P:W��KY�<<>H�t�[B�J��q��7�r��J�!v��{�e׺lqUX�3A0X ��,�6[��9��Hm�8��O<D<�.���,�ĉv'A	�H�2y;�n��#0_;%��@8��J���@ʢ�:Rp�LVPӆl��H�|��^<�kP�@U�T�?gF�T�`�`�^	�1��|������8�� Y�l��)h:��Z��i)N!$���*6!0�e)����?��Au��S��@
n�K5�>8}��q�p�}֦�Ծ��+W�:K�T���>p��M��%��-Dz�mH}��I�H�� ���Wa]� �܈r������Ykq�H�t���8R>�3��څ-�d�6��GYCZ6@�Xƴ��H�%�F&kAئ2x�pdx�ڥ�Ǘ�A_�8L�i�-��A��;��3���QbfGT-���6��phR��B���e��Ųʻ=p�5kW��U��1 �R���:. S"�CDSs�6h�@��/����(���}/�
N�c�7����]�����)i`�e�����JBp iBX����t���]�`~
��
����,��Npξ�!LqG��0�K���u�t�N^�S�K�k�ֲ�{����m��٪R ��!/��B|�P_�dA1�`Rɮ�r6�@��udb�*4��~�)���p�e�bw�[Α
:�sξ���hToM�h�VLjj�7�RZ\��������Ғ�����e�ը�,�,�����Ȑ��8P�v�X�OG�it��cw"�R��/�|�����w�RD,B������-8a�Ȏ_�~��je�h���v{�"�E�pK[�׋��o��)(�[60�_� -S{�پ�����X�F�D�S ��d����w=/�w</�����a������.�`�J��ih��H��bY����������R�����4	2}"tKq�A/��$x�ƶy�Z-e����])�F%���2�NcR4L�@@��*�������Ď�3��Xy:^�FrI�C#�ac:�&����%AW��.}[�W����ɐ��Tk�NS�&�@jmT �j�}�{���~��A���I�@,�Mh �t7�1�n;�Ɛ�FA�al�!(����az�ڥO����7�� �*4��՜������R�N�.�$ �����I�R̦����" ��'"E�Ra�LKC
tdb��A�J��3)V����Z
�k*�YJ9>Y/�f�K�68��^$&q�'���R��oI	���m�-�֫r���?�T����t�zq��~{`����U�n�{������C��h)Cpi<��n��"��a�Wl=���F��~�ڋ�-*6���ݢ� �����	��ġ��D�;\����1���KCL�����Ą�Oܯ��D���?��CC�4�����8K ��1	#n/pO��cTK��<e��B0��h��<N��,s]����m4�,IiJ��BǱ�e�Q`�ԘF�F���9�)w�4�����8dLxX
0��&��<Jx���Z�(q�BHY����X��vW	W8H��l�`�َ.��3�\�Q%�/P3Pl�P�oI��8f�r�Y����-Պe-k���jg^	&q[v	x8K�#��L"0�vE��Ǭc7I�u&���M��NvE�v��u݁"�<�-�i�ٖT1�Qm�Cp��$\���*>N��۩yc�mS�|-�mdU͙�� �O����W[^���3����wR �*����o����q��H�:��6r.��TYU��	���u��nHMy��?��}	�vk�bd�F*�
�tX�q��I ��������pA�@��'�`) �iF�!<�U(Pxs�-,��n�U�\R��5�Ʀ��r�W8�6�	�<��(t��mlU,��� 8��F�����*�&��05)��R�� �W�Z��eMkaY��UŔ%�{�v�Է�Ԝ?2s��h^ D�i�Sw��*扇D�\	��a b�J*o��MD
ΪJ!P�f�#��8p��X6�m�
_\����SF`��<���%�`:�-�&�7�Ȗ���*������5	Mkl)����μZ- �]���7�e'a.��	�(��V�e:��ud�#ׅH[�T�=вr4U;qj� �ɮ��t��	9�֎dS��2AM̀��*�dJ��m�ż�9�JQ�i*�jY�Rq�r�-Y"��&"�X�cT�,�@;L���!,B[h�@N�`%�W(U�,�xU�uo��yx�,�%��/J�׮S*{W?�S"]n%�� ���Ϫ��xuǯ{8�N��e��I�)N_�F�e��T������,\,P���V�R� j�t��"d!��n�E��
#7g��jd�`�mG �� -�����*!��N��RbsYx�����Ʒ�wEj���[6�I��Z��:F��)hT�>��2�O=}�$Z�W�M�xK�)��[�%��ŔM���|x��@��eS	,I��P�j_|z��,���pZb2�r���y��Fz1KfLG���@��cZ�D0 ��F���m$�V�ο��NA�@jCZ��$�0��	4%�u�A�ͣ
�H{O\�ɜ�F��W���څ+���ڠv�6-�G�T E�����d�7���;:���b�&��$�{��TȺ��T�eU�bB_�@L���.|d]"�B�bU�J��7B���oQ�$eL ٬���!�`��>��/��g����4&Ś�g��ư��H�[V�w8�*���X"8R�R�đyY�R�����%�&k����i���!(�tn��J�Bhpq��8bA3��.�RVm%�)��-�I��Z"&��|�4�ߥ�b�%ҝ��B���!,Bc�P.X/�6�Iz�J9|�/3}��5؛�����
����^�8++�,)�)�mJC"�W�R������Z����+i). �����3C�.��b���p'��_�o���؉ۋS�;��{t�j��_SN�� i���t�4�bץ9�R�R�W�r�$d[�����i)v3x3䩑��R2�X�D/���R��y��Ap^o.������k����5��SD3
Ϥ�@jL`�d���Z�&"FP�]c�rd�}O����8d����mR�A�#5�)D��__'�bL"�i�lf�$��@�S�Ev'��ґU�K�ϕ<�0�M��9L/o�⼋��Ր`�sP:ڋv��ļ���Z�&�
������D��4M�#M Mx�9H�z���i�<� +aD��KYǲ���8����B� P9�v<Bf*:����8(Q~��_y�Au������_	�/�z!hM\l#�R�������X&ْUr�\
�Q�(�:|��D�Z$����h<�b�bi*1�g�|��<u^,M����q��h�A*e��]3ǩ/&YR�D܍h�X�5R���Ͻ�F��/Ȩm�޲�9�u+��vA�{#"��ҝ�]�>s�=T��d��H���;�������%Y]t��]�ǟ=���M���@�T���7!o� Kި�0���V�4L�l���4��ڈ,)�tzE�����}�C�#���T�HU�X_�##��ҁ�D3�*������y�Ô�t��ُ@4/Cg�2�)�i����H`k6���.�B��'� ;U���v���1��ӓ;���$A80c��_�2�r"�6�FrEpL����ͮm�2�v��
���.kr������H�R�}�:�\)�x�Kj�;�Rh	B�3�"7��	:�n]"fP訥\�3��A����]�v�a��YH�`L 2�T��#�j���B��pdK̺�8"���H�p�{��]�8��\ ��8Nj�����2�    IDAT fg��\��%�`��og"fR��u"ɦ\���)i~���+��:�kW�B�W�x8���f����������#�\��d�7M�Ȑn�����.�hL�T�����)���Y�&��+�B����5ALFĴ��@�=nپ���q�w��.MG�(P��yd`[���w���d�tf@�V��o�E���ӉI�G\U�f)0d�
��B�@xV� �,�������$�vtԆG�6�b�F-�oB���l�"��m��i�vGA��y��p��^���4�td�Eˆ4d��ׂ84��M��>)Y"%����S�)W�W55�~�VU��j�к(j�������I�^�R�9�&����6|�ھ�!�����C�'�����QV�X-��1�s�.�,r�m���`ٴ��t9�7�q�р�J�fل��H��&k�tBɪ�7!�el_ulN1AY��0�����62�K��h�"E��sKY|4x��B�C���`i��lL1���r� )TҨ�cV>�hRۋX6ZR���S +n/���J����4�,�?���S˺H���AI���^_�c�L�MY@*P��n?�T'���p��0b���؜0Y����P�i�P�8�S�؛oI���YS�"�9#� ��$W���4m�A,�=�Xs&%k`K-^
���Q%�;
��\/��A�8�ɚ��#�:&E�-6U��L�� .��@՝Lhٮ�P^Ӥ�Q�����7�&T��6�e�q�w��M^�|Ӻ�>;�/وO�}(k�
��׽r�Og�O�.�v�H�d5K�,f8N�)h�)�
����
 >@1}�����z�4	�Kiԇ���S�F4rb� �/eT_���l�_}�U%R髥d	�5n#�RƐ5gY�u�)Ƅ㘟Wҕ�{���hF���.l�n~m�l����#����D�~#񬗭��	S0ɤ���9��:p1�穑�W@�] (�X��!X��,� (������f"��r���;gY:b�,5M-ᐆWg}[%h0߮������KC�pn��@�7o������2�[
�^,e�Z-��G����9A�T[�����)Y'��%+�ܮ@R
�X�{���Ӂ'ը�L�������ȺR�񝆣���B1Ad���q��
��Ȕ�4!Pk��@��o#�!����YIj�J��f�V,kY�,K�y�������;��y4��%��/I�`���4m�<n���5s2|1D�|�5]��d)��5�"�C�_|�q��O*�e�ɲ�ZX�K@?_;
����H	���*(D�t\]e1�)�}��׶���Ƨc6W�okD���Џ	1m�����}�`6��L	�Z���k��Z:|�H֨��$V^PQ���#�u���Ul��^�̖��F �l�ȾҔ�ͳB_A���駟:LU��~�H�3�ׯ_�sN5ە6Mi�l�z��ZJ�R-~�p�41�^�v���ڡ��]�B����@h�N�M�ZZ֎O�&�X��%O��T���z�b��)3P#�ٜ֨|�y��J���d��<p:�����5��� h.��VXff���N�`J�?R�&�����!���J �9��\��T�A�f��Wk�!Jy��f�L�f���+ӧ��K'Đ�+!���ͧVw���p��l_|�˳w����6M�T��BK�] [�%e6&f�ji_�W�3^�.�M@��%�%1c��A�d���[� A
��!Mg @��[V�|Q�)��em*�W���!�� ��O2��]d7B� _���;R�ӓu�i��<�Bs�|��gR�\D{q�h����r��}�)pѥfv/����t���Mw����$pKO�d�Ț��>Q��0�BR��ڨܢ���~@]<.55��P93Tn¿���ĉx��0��)�A0�r�p�*m�I�7��}Y�l�;�%Aq4�Q@�H5����t( S�o�ݓTؑ����X��y��Y'7@�X;�F���P�j�#�#Ѻ4�9�W�^��?�KA�lLe�8�޽Sq n�J�&�o��C�2�.�p ��T=c���~��s֧�'?����*s��x��ā�i��p�q"�+BJ�,\/f�U�MlH���PG;���r��B��yBx��Z�BUpwD��&N�TK�#�2�8�N�љ����";�^_Ʀ�"�Fj1���[��Ql�hnW&K�����?�!�	G�7Y�D����p�H�,Mˮ,�a�QE��T��F<۲ D�/�SS��&�ix� YmH]�I*e�NQa;��4�YE�2�J�Uh6Y֐._�Y6�5եFyS�������Ry@������Dwٔ�U���3N��t�6G���������c
��R��am
B�%>�<�>d�U�LP��C`å����p]����uA��Z�dmj���DP�3��85K8�J��iW���%в08�����R�v�/~q>��t
d-�����4���Nm�4��K!�Pk��l�}�i�.�Y*[�ʓ�Z� K��^j7@Y���
cB��j�C�ߒ�#(�)s��.MS�阾� O$Y"R�!@�a2����̋�'1B����cg��W�o��q�YyKz�y����Y����7�e�c��9�8��B��.�"c2`-xʼ.h�FX�6K
p˘@K:�Z?�n�W�{5�l'���L�ֻ1B��͉�p�+n#J�@h	�-/��{l��Dܽ�GȫJD�ɴ#(��jmx�WIW|��������w ▤|M� &�u�£Ŕ�A�,�l�č�B�%.�괫��]S`gg��	���8LL�ZR�7�]q�v�G��r)����ӶR�Pm-��m�h���;���E��8������M�Q73�H:hx ~��UiL\��&WHSy��QL!Y�,~�eY1��٦�)���k*N���] ٖ�Mŧ��xQX��b��� Z�6U�t�0��I��g�ʚ�v�1�4�ח/^m8���h�⎋��h���Ϫ>��
A`�������[��B�G%�b8��}�irx���W\, ��Q�D,������ŨR>�� 샹X����#��8}��3Y oN��1�Rb�O��I���o���<>�7/�+��� fv���>�ө��hSKMŝX�ukM�25��\�:�2��m����	8�td�D*���DVI��f�&�Ԛ� �O�h�"�P@S̤��-�u� !<k_zI%�~�� �^v!�\mU�
p�>)K�I���������A�g��4`�n9���J|�w5}�jl�
j�F_#Rb���굍�+��#�a:��6Ί�MJ���Y[�#̜ NK&Ƥ��
�v
Rs�:I�vVe�a��e�h!�6~M|�hP��2O���|�Ơ L0&��ZF+Ƥ����\����\-�=���Ac+�]A�/g���Xʲv�LP	0}4�킇C�C�mm���T�F����ڂvttq[�>/�W�T�/����.	�v���g}Y"����`6+�:vL��'h��pq�H��9�&HY,�GCh��8�eļ[�ܮ�-��B��$����L|Y*�7�J*l��hl:b��ti*Kq_���!����:j�Ȥ2L"z��&�@��f/y�@1q#�Sŝ��9�Q�������i(�d�ݦ��~��W�4)��П��������s׿��G?�mC�9�����ћ^�&C�?\��K� 45Ao8v����8�2���b���>�j���&T�WY��V�e1m�d�LM��3�����G-���ߡI��݄jy����h8�/���`%L�1x��v~~ێ�g>4O;�A���EK��Ӏh��ɳW���o0�F ��T��O_d%����ׯ��܉�t��W_}���_ݟRu����?�Q���?��ϔ۔���(ӧ�f�Z\'x�!P��le�;�؆ؠ��6�fu��=�[�9ؗn��ͻS2���::嶯�p-�3��a(��恴4�]��祘�H���L���o$��!
�yq���B�,L*O��4B�Z�R����J5�F��`�D`1f��ۅy��
!�X-L��6 ����\;W�i��dRޣ��ý��܊o޼q�����Dp�nK1P���ۑ������<w��� ^�GGO�м��d�5��B9�V�~��B�W����U�v����p�6�{�������#h�5K )cX����]M�-�#L
���X����{X���ޕ��r9��^��I�V�i�� E��^2& �ϫ�x�:7)"^/u���/ͩ
�c�-N��Nҩ��3K���`%t:����i�2�N٨p��F�l�w�����V_��1�[?����()�Ɲ������������F:���A�ex1��@(+�3:-!�2�� e�b�~[JP;Y1�M�zU�ib�h*k#��8mi6�H����Q�񯹟�s�^��|��?��O�:Y~ߨ��y�:p)+`��M.E�M�c�"��,v{�cץRJ�x%��-��g8p�f
b)U!�2���k�y^��I"S����Pk�fn���T��J��&��v�PɎ+�8Ș|-�.�2�(��$��x����A�mM�)U�<Cn0q"��,�Q��{� ���x�*/P��֢�lݻ.d�²<P�Bq��t��N�hZ�
��Y��8bd1����5��uTB�T�Ԥp�
ꛗR>�Z�U6CU���e��eU��ٲc�j�p�z�c�pd&�dS�Ǆ�!��d��d�%!�2�V6���!ې�)t\�R��Xj�6i�ċi3�Ut�D0�R�+�Դ�����J,��{?��c�|弎|3ČP;�,$���<6R���xw�=��Wкt��e%��MBM�c9g%T�竬	��N��hy���i�yx{�E
'�f�Fv�o�D,v f��C*q��PaU���	�Z���,���wD��q�����_#Y�U(�ڈ ������?7LY4�N[�x��,Hª���bR� M��󧌙щ� �i-�N>��Ii��yVI"u�R�<YU�+�ɓjY#���SN�2���}�@�'}�^�m�BNA�rH�#S(kY/��ꨊ�"�N#<f���d63f%~Z��V�ڍ�P_�%$&�;�*����D�8D����L��1y���9��ͳ��8_�����]��/(+��tp�s��h����t՞���Jx��M��1&KJ^���q�e�фl�Z�*4�՚_Ό�~-��%Z[�5EH�KF9T%Xk?�|�&������ŵ��B �6CR�x�>���I�R.ՋW�`���>{��� ^���r�*�U�"�3�O�����х����)�D ���"&ېRp3�h�����	f�qL�bN%��F;��d�vR� ��40��VҦĉ㓅��3T��p��d���!��r%���Aq�h*��*�bje��}f;��j��+��ё���!jC����31���2�B-�c�1�hY��p^J�Kif%�B̀O���B3��/�(58r��囥�j�̪2�@l�6�l۹���q{�$�-V%PB�cv����l>�T���Y�IѷA'�l��guw��8�;�ߒ���f����!k*ff .��_���"bxL�f�kã�� Ȗk��W�<�T[��G�u��U)3�x%d�����	"�#�����)i<�5���i��4!�.q�e����.�L��@�8�T�L��-�5!��!��|}qb"4dw��RZ���w2.P��Z�`b�іA�ީh�z��ޜ~xy����~R�"��5j┓�G�^ϧ�qo#R�p��S�����["kW/�a�B0���N�0�Y:�CS�[R�*��]	��T-���u�)�M_���`Z:F�b|��朦���!�g¾�n�qv���SA���m\���	b疶�2mz����|�ڳT�DS��������j�7��}�Bӂ��o<b"5U��HaZ�1������� M������x�t|��_����� 8,�c�����m '�Ky��4d;rC��B��Q=r��q����!��	wȖn}֎�أ��F������.��_kxcx��Y�B�ٲI���z�q�������i����?��/4mgH�:��lŤ���_��0�.�T���(訵5"ΟWnH��jI��m�gH1qڑ;����_}�A klcԨ^���/LL��k�����e#����*[�Ԩ�/�1 ����k� �9t�/�D���Ԙ�Բ@R5jH8���@�πb�Z�Y#��h���$�~���O����6����~�r��q�Xb�nE���eu�����x!�C0�8��á�Vw�j���U��8F�n	/"�+����ۆ,2�*���sn�@��G�A;1M��fY����r՚��)S�Y��	���ڂ^6��?;h�^,@���>CĨ^���ub�;�6�c����5S⏼�{��WJ�)�ɥ�,M�gr��M�I��N1�:��uT��X���
��3qu4uvѓW%�љ����>���78YL|�� ����S��WbZ���
�H��k*1-e�������p��Ĳp�,H��%&$�i*�I.0f���w#ɊkG͒[*A��*dR�p]��&%pV�@|d������ ��xNН����,_w��E�^ι1�0�Y6?r�r�hJ�?���Zp�h�����h�t�
����`�D
"0RHUV92��i6�!�Jݔ�[�DN�x��vD��)C�b���	Z*i��l	gM�a����Ʈ������ �F�ע�B��i����)�#G�*ߝP�$��!�XSA��H1�� �ۅ+�^ m��hM��S�v�_?�
��A�d��#���������Y"+W!D���%5<��lA����,��B�BӬi|c��Y��$�\m�!�k�N#��o*k/���iZ2�O*5����eC�!-K�D.nl�����#��>A�B���5�v��s�Bֽ N�ei�2K��@�8MC2"e�!��V�,����)پ�F?�j'�p�F�f�&�1��4�T`�2X�O*�E�¤�RV9����X�*��-��T��%�lu��* �� ]�h|���/+Ya��g�vL�����<&/��۬ ��Nز��Nj��R�eʆQȏ7$N����+�PH>e>�~OA��غ�ٮ"�=�z�c&��^��!����c&ɒ���2��;�9��Z>}��W�X{��Y�yn���j�D\)K�;bG�`��6��v���eu(�Ȳ�[R[V�3�mJP߼l�|�b�
�����Y�
��Ip�v��&���|��.fj��@��|��� @�Y�o�vD��Z4�e��.f��.��G�y,5�b��9�+�j�U	j���ٴ-�1V[U�h@�8��C��^����gb�<��X�yB_���REM�i-.�zY���G��KU���B����Zb2`j'��}���kaː�
�C"C�J";(�J�/�'�YV�Y��d��&�۵T
bU���yd�>����O%j+ox�������Rͣ��i@��>>�Zv�ऐ�e� ��y�ZM��,�H�9�,5�^}���%1߄|K��mh*�fI�"�k������<�v�P/���i!f�Dn�@� �Q��<N���æy R�@fYl#� �\�l����ވɔ�e������7-dM��g�ƣ�X ���6��8R����TLY8G�P�cyW��b�K-%m*O����	��W"Ȳ�O�>����E�C���kǧ)˔3���m<%��A���/�����n��	v�t��*���
�6���� ޲���T�a
,ǉ��)бkW�%ZU��	��)�
���ۂT
d�"�0iz*�6��Ɖ�\LAk� �<)�,Z�mL�����z��B�4?B��Sņ�0�z	�����0�R����-���S�<M�{N�A,����I!3�C��+qY��ӎ(w��d�_%���L�*%�Ѐ�hxq�0-\!�����;�Cί*)
�'��$����Ĳ�)�z	�@ޒ(�R۝i*g�-燗7OL�2+@\    IDAT>_��'-�<B�Gx[P�Tij�&��u񢾺����{���*'"����	 
�o˖����� ��YL�R��w�b�h�Z��,S���'n	Ƿ��6�rYG��lge׾d���W����\����q}������:�p3�����o�� ��`�
�e�p�쇉yU�b:�k����-if��c6K� �h����`� 0;�毜N(�:�� �D0�(�Mk?J�&�_����?��!_%;"}���05u���$n_7.빦'���_%��j$З>Y�����{������/������wH�x��jVbam�8�4Z1ٷo�~��ߧ�Lef���!�FL39M�~�x�����/�{Z�ĘK�X�Ң�+~��9j$��0�|�����ۯ��p��ff`��7��R�`iT��I:.f<K��'j�����h�/��&f�@|K�-
�B�4�Σ%XK���2K"�5�e��4�%&�Gw�=�3q�F���l��5��d�$X�#闪;)H�0-5��ø��d���])��=O͍-Fv�������]z|����7*5��Dp��m��M��ziz��4�\'#��_��G����۟�Zณ��{YyQK!0���,��뿈�%�A�M���]����4ܱ̃Fq"4�Q�xΧ�3{|��^씬]��`�J���)��?@K�Mk��Dfd)���-�ܦ�~uDp�e$c襅�P�Qț�er&��m6�!u�)�_G���tqzΰ-(�
ZzG�Ա��N�l
�A�������-�x�]���]�Uy��������F�t�Yk���vJ���j{Qt�I	��bj�bU5�+/k��pjO����#874��- q�R8N�K)�*kS��uq��O�� ���Me��Y���Et�����V e�� P���0m�4u��Cd�y�^�*w��@1�v��<B37�e:RwAj��0������ܥ�2��
Ŏt����ZA��34 og�$�/�3P�`Zf�"[���p쫔�&�ɗ�>��IQp�����%f�U䙛J9�ƛ����k���F���-Q-e8��H�D��X(m�d���5N��j�&��Ł�h!Rx�N ���wt�b^��-L�&����V|QϮ�f���0kA9D!~��R��"�jŧ�cZ1�y�-�}�H�l�đ�*�N$NM�"S@�
��aȲ���U�o�4q�}��|�{^�"M�L������ò�@4��;��ƉD#F�fB��U�VPB�j�F�%F��҈Y;�ԪM��޵�Vլ��z���p�}�9��s\�}^hg�G�D���EŌs��C�������9��h��ڠ^'J[�)�!�*	de�7�?;��3���{@�����n1����3�pc� �� ��2�|M#���h�hP�
҄;�ȅ`8K�KčU@�@"dF/��r	'5�V�X2&�b_duz�����U8�c�$ ��)�w9jG5��xl�9�c#���vI��w����`� J�ZOȸ>�t���8����F�}�o���W(�O�k�^jô'��S$�K��Q�T�g��mI����U�8���x�0�ʰwiw���z��jT/|7�}��!�a��h��B А����}��K�J5|8$#�4Q0�SqC��>�W�Q3���l�L^eΕ�\ǃ=o*���auf�Q����~��Vh�EP6����N� g��1@s3e��T�9p�Sbمļ^K��# �5���Qk��-�����y�����4Au� �����FZ!�m�+'!���:Щm���{��t�7����Ī��z�h-���wY���z�S��S���i�V�4�3�Q��hE 2�3�֛������9ֆ��qN4�xL��h�f��8���F�׷K����a���p �j�d�^V��bGR�~��K�mE6k��^�ǱK���}x3�VN�B�Xv]VP竴	�;��<GH�}n�Y]�����á��j��ۂ#�]�75Nh�_�����Vk��_[�P�:+�l`b}���h�mV�ϕ�ݜx8����KR;�=n9��^[N3�akO�f|�ã��q�}���yl�yw��L+Z�{mp�d#d�9ɚ����}�}���i��QM����MM+N�nV���8���=͍�s�"��l@�d�AR-�.���go�/��+�\�ԡ�8c8%#�%�O=B�f�]Å/�u��~�:�ncfh����������^>-�g��6��֫@]�9����ސ:��6+����7xR3+�HҊsJɶ���
�˾)��C���$�E&6B�E�sd�b*��>N�spR[�c%uMgh���.�T'��g�fμ���,٨����.�p�sj5"# �����!�FLY�(S���J�]?-�����E��)	�ӥ���~���O��oCM~�Ǵ�X���3�7C�~��T���'�c��WS
�2IY����EQ*q��5+7�*Z�� ���M]� ���\�ܦ28´?�.����J}}�&�##����۷'���-V���䀨a���4ț��{�Cu�R�1C�����sO���~r�I��}��j��6�p�
���{�7\���y�H�N�r,�&�%����g��,V��}I�
�=��+U�ٕ9+��i@��)r��s���}���W��j�V2��-9j��
$]�g������ �c]>V�S��M��U�ϥ\OxشD	p��(�j�W ���JJ�D]7��p�'��,�U��z�)yGԶp*ʲ���	,�<\��C��&S�8T���c��()1��~�'t���F��.����X�h�� ?�~������Uk���w�J�ǭ~I}v��H+����Mp��zK@���nn��_ݔ�>�_8���S��j�[Cv�p�����}w@����6��Eҏ}�Z�ث�=G�mU�����U�f٧� �K�	`���Z���,k�F��<���Vi���}f���|8���}�u�$|��(L��eT�E+<*/�V\׮t8�k�֢óG�Pc/�'6�)g�̪*7��}�����C�u�cw������rPP�{�`�K�#��N����[�n#�e�%��ڇ��P2`�<c�:�Y��6��<JX���8�ȋ$�G�Ct�p�H�]0��"GO%gݽ����dZ��#�
\���& ���Y��.T=�5_l٪�c�����3i+�h)y�Q��l�%4� ��F	�Y�F��s$����ʜ��Y�B9��.�8R��s�,�*�|xE��z�y����ۤ^xo`þ�ض�!�R�KN��ܼG��E���/b����(���`V�2���.%��M=CA�M�P65�A���Ȫ�=d%��l~�M0Щ��l٩� 
'9�$O6eq-�|l*����c��$�8�߇w��:���N���b,[��0
	����ï��T�e�Om
�k3~�<4o(�'ڞ��j]DY̕	Pa�����o F�~����#)c�U�����&
q�Sύ��~�yY���|�H)d�Z�t��G���Z'�]��]�X8_هGlM:暄����Mw�Ւ\{�%�_"5S���d�u&ZT���tZ�.�;�0��Y�/�(Y�Y&�8<�d����&O��Ƃׄ���~�$̋�<�&�0����S��wŐABNĮj&���&�9��G&=A�'Lg���Ay��vXا���lA��|I�rpG���^��V�D�P�{�B߽���>H�)UVWrA�	����k�0p��	�2Վ� B'$/
�)1t8U�^��/v��-�Y$�"E���H,���G?6��xj�x;�1	����
�xn�}d�6�l�D�a����$G@�.����~CBl�#q�ǩ}��o�H�����-�0���[�eՍ���G٭���9��Q����������5��u�ҕ�ޛ�![,#�k�''�κb��c�2��c�{ٮ��<Z�ۮR���V%���z�k���3�$
Wca"b�������x��v��B�/ҥ���R�_3����|M/���|�E�n����wu��ޅ�WNW^m�Sl����~�$6�̅{�k��Y��*%�LH'f}��U������oNv:��v�#�Ӟ�3,���c{��4�`���O� p��T��sU�~�8�
�v��e�&W(��q!�Jw����n���4����fɀwrĮ�Z�r��c4�q�5J�v��V��k^~"���2q!�+���ܜ7{���fxg���8C�k�9��� �,��O�Y�AbD��cz��O���g�dV9�O:N�6@����'�-��X0�y\�1�e�����������W*u�.u�7g���'xE얶Q9�E��׸5ش�˧���<��-�}�z�ϸ=ė&�l/xd3�6���R�T,[��Ҳ{�:"�GJ9G �N�G�J:֖_������Q6�̊�СP'�bO��d��cd0(�1�..�f�����m��ĄN�`�p�`U����� ��!�j�4����1xċ�s��;N�}Y.� �;������,Ź�9T�K-����j��Q�[�����=8 H<��6�͖�m3���]���oaJ���>�t��j��%�k�45���S�)X�E�?I������F:_<�u�{����������3S�*�%ïң��%�n6�X���VV��`�d`�4(����J姏��D�r���bA�CL�d��ִ�[�8���T����O�����yaj�é����Ē�@@��(��.�<;Ί����^ņ&ǶE6\}ox�����7�!�=u��4ջ�)�ʬ��޿���,�+�ı�'�k��a�3��:zX�3�ׇIǼ0f�k�{N�9���]s��`Β�Ux�~����L|WqbSYítS~>�D �~�H�"tCv ��=8��<�{�����䂿���1��ڴ/Q�E Mpt*�?�?��0Qc,�ɗٛ�!��!����ñf݊&Z�@����h�:Ď�ӵ���.9��;�O<S�ܶ�#]4���vxp���9�C��K c��z�m!����#ސ�n<��£�e�#.��-q?+�
b��s�A/c)�$�B�96�8�;TB�?wj2A���}�@X�,��.��J�j���-��YM�>�@��˾q8�T�O2)�
��T�*��zoV�߼�����N����+nb��t�������
�Y��I��/�}��\Y�+���䜗��kv�S��W\ܾ���=a�_�⨨���v��[9a0@��?��j#lՅ$���/B��M�qe>�Έ �Q� ��|�١�t��w;"��<$ *�2��.�Vo�-H��;������t8��;&ˤ�W�o�ɒ�m�:3}��Ϸ#����C���٣�y=�ȷ��E�#m�t>zټdp�%�%�u%%�lp�I,���N����^'�Q�2����G�f�����v��oD�B�6�h5es��[��(a}�9��
Z��}����ϸ��,�o����`)�� G ���p�@w��� `�XMz;������j/3�#ޢ�cp�1`�X.��NH�gmee���,��&����9���0ι�R�b�x )箠|Eq��%��W~ U�t0\�xрg��������{F�8�����)!�ȻG贬!#.-��6��,Ǯ�k�F���E�����-�\�dE��K��h7���ɘNS��t�|�����Q�N���Y�:k��z��?�������O��~/N�[�����|�thr׵mw�
I{��b��?�C��i-�������R�6��x�KD}r�/K��+���#���6��J�r�C�.��N���$�BIwυ�����^g~��V��R|�y�nω��Bf*ґ�<qU"~
���B�S� 0}��mԄJ��l�������d�8�|X�����26|t/�%��D��۠t?�m�eI���n��|������M�㿟ޞ)N��v��"���E��H�+':�C���X��Y
Yߟ�I�q�Z�ʿwd�O�\A��z�hN{�.)�W�V�Cq�ci�$]���ݏʃ�D��_w�>��{����u�%����VRK������*�MB�<R�K�d�.��e�Sj�	��sNZ�7E��#i�Z~��˩��zM��י$�w�+^���-öh��k�^Z8"�
�Enq�QFvzA	i��z�H߇N�O꯷��	�����%To[⦪�Ϳˬ(�y[�<�M�q`0������l���p�2ɛ�=}!P��[km�i�Z(wd����]b�T�<����es��l�:�{�(�����rc��X�>�c��B0cX�U�ș��[^�c1|��}���k���'u���eϵ(�-d|ʇk�qy
����/���c%|0�?/�0I�lẕ�a�����'f��׊��܂�D���Vi7�����^z;����s��w@�@S}�s�6�[��_B��al�#s'�')'�j}�Uz�l�Þz}g%J�.�EDDӏU����s�����xDyvN�[�P0<��[��W#ޥ`�y�,���{�~8�^W.�fl92(�m���dVXq�!��ތUZF�u5zg��������]9c���0(8�Bʐ�^���U�oUg��$v�n6f>Fb�8�h��ޛ�EG� �y7�P�q����*��k�	V����@���MvY�,n�>������r��O:���+�9���O�5�.�c��������X���՛��J/���{��(bG_I>v�fL]�B��)� �8 ݾٟ��vk�w;�n°�yX������;ݶNWO����9�Q�]������/�gm�����������G�d⹛����&B�v��!9[�X����a�o[�1��������lrc�FϛV���aӸ"Z�Ⱦҭ&|$z9N�[I"�����d-4.o�P�)�LXb2�҅`��+�n�U@Y>�x'��Fo��?�� ϵG33΂�Ր����^m6��t�����v�1����#�z�d>���7��
�l`�
���w������+�W5o���r)H��Hʡ!�i1v9�ϑ���ϳ�~�C�C��#J��o��zW��� �s����b��C�V�M)������2����o�K0l������O+Gpmwn�$"�t	{DJ��]_����e'V�|*��`�X���ĳb?�W��B��Q�Q��������e3ҩ�����_����#��g�"Y��7������M���ٔ��#}�گ�9z�����#��h`�R���:�A��r/K:�$��/��|�w�{F���#,zVt�����'�kw�[z��G�*��r{�ߛ����AՖ���N�eu'5��	�,�'O�8��]��6�ۇN&�)M�U�ίH�a�!��;D�-+?a��_���|�M��j�`Q��7Ռ~ᤞ	s��9��3W�y��_X,˧
y��"�U3VQ�����/U�ߜU<��P�*Z�v݉0a�C���֧�~N�k��gC��Rޢ�m��-���\و�a`�74!Kt<�+?��%�,CRFU^�~G�Yj9����)�2vO�e��co��$��È�0�7�CG�c4����i+�>j _$�oT���b`����	�O��Q�����&%l[�����W9��V$ʨC�t-[{A�>�j�;�j8��x9r5������#�X/+�u0eY�оU��?�᭬��w�d�{W�.d���:V�ǉ�n"�b�E�|8Ol[0N��p�V�6�C���َen�ȤKi3qT��b�iX|TY(��1�(�*� 㪤�^#������lIvŁu��S�_k�	�Rjz.�JPM$䔰A����ƿ�"z�2}a�h�9f|:9qb>�Q=/mg p��A���]�v�h\s����$����F��`�p\�!��Y֨�� r��%�SA#蟯�4�R�D���Ւ� ��^��Sģ>R�I��q-�pDo��I�ce����@�iZ��N�G���A��i}�x6T~��v�M-UG�)�If�����)��Q��q��ݒ�kl�S�T�I���az�{Y�i/�NW�'{��
������E�8���L���m��R�0��X�Pp�/��QfN+�~��%�)A ���s�^���s����Tư���&G@�����ތ��j�&�SύʗIb�)�Z�/��2��Ѣ�'el�vw�6<D�e����$�%��fY���J
�����Q�GD�";+� ݱ(�h����2�h5egah�q6�?��UB���'�E�V*�`,v�惸�E��CU��d_�sEO?�����	��E�\vQP�/����z�wcI-��:Q\uQ)�K�6j�	�zUp0��RgSmENK��ߩ�T��;�2N�7/�&�u�:�1����&��EV���@���Y�匈F���v���*���eR-���]���̅�|^4��='=��y��[�h`�@7�ڒS*�K���$��c9s@x�@]���sy~��-x����� o4Mz��i�G"�M񏼰����~��qT����;o���b���^Zsl'�����{�����'�)"������ǟ���˱+rp���-EJӤ�$�8.��O�İ8���5G6e���ex�h�ðP/���mS�c�'��^��#���^�M)[�At�Z.�|wXy��Bo�h4��kC��߈���L݈X��a
Ѷ���p��@�#�u�ɲ��xͣ�:�������XF��l�R��JW��b��3hWٹ� ��M�
%L1;q�����(0$q$�u\�F�����ⵟ��d���r0{�;�Z u�T5o¨Gc;:����`k�����B0)50m��~���S�9nyy��.��Z�J�ۊ��nfJd��"��ja�tmh�*�����-Jg�D$^�'������6�K��Ɔ B]>y��O3��N�+��5�f�2baIkV�&����<�9�"�xzUu�"�RGO��@��1���}G�(N�#�њF�_N[�8Q��>��7*����Ƕ5cy�˹o����=�Snrϓ��-�#.�����~{-�d��|z�C�x�Mގ�>=w8�P�y��R�ѐW!�@�4���Mqv~|�{.]×��Vj��S�G'P�/�D�Fc�ڵ�e=ܢ��u�4��OlZ�!~Q*vm��ݞզ܌i�k�k(�����otZ_��fۅ��5�g�����Dsl�;V�q��f~�������yR���Ġ��W|�Q���Я7�
�c���;u�v{).���M��7x_j��:;���[�?���G~��J�|������	_��g�ݓ6'  ����G�����GV�����-��.\�[��3��]n3�٨i4�XF�!�,�k%�0��f��:-g�~��l����j3G�3k�*�Sn�Hj��A�"�9YUz�_劣ӓ��)����-��*�l�aI��x}j4�x���
�n�{�ptҠNu�P�������D]y颀߱�h�a����1������� ���㉹��.#mN&n�������ݙ�[.kO���8(0����B�q`� �i� ���͓��D�o���5h0���J{��Qj4�I�v��n�S���<G�e,�`'�!r߫��Pc���~=k~r8G��<��>����׼|X�{�����Ű�٢J��?IGT�g,�>��u'�$���֓���Bx��h��um��"4u�&v,1�Is�Z�nU�DE������}#���@�	�3��
*&E]���"�bUU��;i���^��$��n�0�8�^r#�=H�7�/���d2B�m,�}��aB��$��vE�a�Ȥ��Ww@��nu=}׍�]aY�q���Qeˉ�|F&5K������p�r<���������pj鞗ɼ#�YO��k�m.�����B�A"��`V
�1q �:��[l��>�g�8���vq�����&R�2��N�Ƽ�*��g��Iu�tJCM�n�t���%�Vh^g�,ވ_�=�m~�c��
5![��֜cB�O���Z�����B�s�}0�V��Љz��r���5]S�ofڃ�-}��nvEdJ&�$��q���^�0=�u�mZ����ج�k�)w������x���ҍW� G�<E�/����F�,�&�m�W��~����?j�.�I�xǔ.Q%[f�2,����U���R�/�M��Nk'�!�%5j6�g�dq
Jq�o�xN.�z����5�ۚ�Dl_C�;� 2�މ�u��gr��5�q'�<	�#�K�����"����χK�T�l.��!"�.���ּ�ڿV��UC�]r�k����qi���*�kN�ě�*��6?�`�v#۾,�԰���
�ɵ�TD�eU.B��u���P����"�A�ǡ�%x:��Pp���nl�Éaw�h{����Ɲ
f�O�7��{iqku9�Ñ�r��RE�)k�Z����5��4s��8~�d���q0������ `���ඎ�C�rKo}�fB1wq	ہ_{�l� �6N0;��T6�?�i�4o1�֙��*<w~q�q{�q�Z�=��c�By�$#K4��1�\Ph5��a�'I�hP6q-J󕔸iЭ�ծ��s#�_�/�/�E	�8�W������(`R��p��.78�~�̖t�e=#�2�;������h>���]��X�*޸����@�dQ�EQ�i�(˥�����c"������~4ٗ��c�Za��/��.�g�Ň����Ѻs�n��3���qs��+B��8
s@�b�u��ML�'E���&�Y���В|���>��lYm.z;��,���Na����c5m���T�tw��
�s=ĝRk����"�Ki(��7�5�}�@0Qj
ˑqy��e�l�5%�«jN�6A�1mm��E�-s��P�@2�*j)��m ��g�e����z��P�]���#\Ӽ��
/���"�3d���F���1���| ����m2�`����9�֟5��S����	P�GP�q].Qn�U+�����Xgy�]�B\L@K,)�";��ѷ�ms���^uD���s����uԀ�6�˂����}+	jy�n?��}�g~ak����S�IQ&2��.�4] N���{��d2�z��z7v٤��Y>�ќ���.���r������(',��3�}�*��a{�R֟���X�7p�GP�O��#CC����Ծ����/�8������`�Д�����`�xm�A�.h��}������ͤ���!�4�sp�-L���%�ދ�tJv������U�k�?�p��@ʦ�0�v����e��ٛ��0��=�|�4�����~��٨8�lr��H�GJ��j�.Xj�e��gr���>DZ����&	a��XV94~�}�_��"��̑B�&�[�=�6��W[ܩ�x#�u�D�y ����;?����=*�s`Iܡ3�����$��>ǿ�n���k����(���S;�\�i+Q�f�U�hm[�f��
�u�+^	��Y���N͍o6�a�i�EiŢ�bDYa�3��m�����h�4�d�G7aҟ�Ԗ0)���r�>��^���ݐ�����Wz�-�9���m��W%��`Q��Pe|�>�WKź�O�G�ͧ�_B1f���Td!��}�B�g�F��f�?���~L�c��,�uW��K�\�j�"�/�M��J�!E�/�Ƌeq���'d��>x���=�</�'��<P��a�����v�9�ئ���Z��)NCԙ�����~�>c����\�.y'�S����у�Zv�v�(N��b]���,w��C��'%}�)��+��1�1��E"�ȇߤ���;d2z,L��{S�'{���y�^oX�N-j���p�kfs�Z;�EpJF8
�ܘ��Ba�n2l@d��21�Y�:���mAk!��-ƾ4��_Co7��Ka唾���Vb��Ci�sxl*���u��L~,�� ��H`(���W��ʑ��9 ;��P�{���!��w%sڌ��S-�R=8�q|O{�a+k#�㬃�t˩��魮#5�b搦��XKV�U����]��&���l:�3�ZK�0E"ۡ�v��s�<=+)�r+zC���	�=��`��3��n;�	vkh]]�o� �-����m=�����c���Z�~;^�K|3Bռ�g��E��VK܃b<=�,Y&ɍ��{�j>Q*g5��zΒoC|����P����;�JLN9E?g�٨y!�y)��=_*�<)��E._t����7;���g{)�?�R��$w�B���jY��Y^����1�b���x�㢢�!+����츇k��@)���{�M���,���vMLB�un��Z:ٛ��Gݟ�����8H�<O�4�` ��%>�32k�Zuz���qc)�����������n4�D�K�����zF�ęڌD{X��.$��4.k��;&d���Iyj�lX\l���q)F��|w㳇\�^� �'��Ӻ��/�|O�ߥ�N�i�����.Y/H�(������m2˻$���;M�x�_K��>y'�R���Л��p+0W�޹A�"�w�Ȧ��vy�4�'p�������ܾ�ě�P��v`����0�D�K�=���*0�$c���ϼ���B"j2^h�g�U;���bJ�@7�c-
�XT\df�)�}y{�;E#�<�r7IB��!e�kc�h ���X~�Q�Cl�$ٜ>��)S��C/<�������F�ѓ�J����}:
�7_��c�4����G,7����+(C(XS�۫������c��0��!rՋb���/MFH�U�j�Y�z���h<�j�q��`��#�d��n�(a$|�h5��4���"��L_�L���.��*��e��\/Ϳ}З۰�Ȑ#on��J���S�j��
_zK1�E�������IX��	Vl�.'��~
�@��'�H�G�_��jTk�ak��n͍���Vxlm��@��n�8��*p��3'G�q�A\A]����c�hV�U��bf�����(�]5@Q*��X�Vo�+�(����{e@H9�"�J�׮@�I��߮��R��S
��!K��_�8�<*!Yu_��ۄ��*���̏���]+��7	|�gt��i�U�s��T�����%�XS:8��vg�C��Eކ;CQx��W3����Z�X֋ǉ ��	�󒅭���Y=s(5{�8�����\��.w���9.ԗ9^��!�].]7@���O��TN�IvZO3�27���4o���밺�GA��a9�o��u�Ԕ y_ވ���̎/xی�l��݌��'�u70�VNM���ʊ\ו'5/��<�Lb_7�=��z��Y�"����J��+�_��S,����텗��7x� �|��i0�pC�!C��/���WW��MA�ϋ32�s���;��R?�+d[,X�ݾ���(�Q̛h��}��x$�oO�h��JA�86���ə�N�&���;co�v�n�q��g�`Q�T���T��&��������b	���@�|E�de�oA���A+�Z��i��ָ�e��u-��P�����O� �+Z�Ӽ�>b��x�+>�_d�����Q�3���߿��@w��h�9�ݣ��(��r�&������	� ��Z���7�9g�~��T=8��(�_U��ѹ��?:�䤘���+"*�XW�9��
J����u�'Z3��S�GkЈ��vv�2�a��}cE�t�Ϡ��Y�{~S��{�����;��Q����K�å.ZL�Ʒ�s+�j��k�=36����AW�����ȋ�焫�����%��ts����F�wm�<������e�1�WI�.�S�|8�\dN��(u�u\Ԉ��әy����b����{{S�{���!���&�k��Ŀ���-��*fq�z'so�V6�s��|�
�����
�	M�-�L�o����r減�_Qy=��5���I��������+��{vR
�a_KV%��vuP��x�6�Q�
3�x<��B�Ġx�x���`+�d�+�ǶR�x�j��� ^�o��
0w�r�"�x�z� �v���U���z�8rE��+�MB��<�g��X�|+4r]�&�;�m�pĞ�������<���(6!V	V���E>�"�PZKiNa9T�].dQ^F񌒡�eT�s[�b�s�*�	.u��B$����J�bf�<��yh%eӑ�s�^�5�I�<�v�����p\����Q���Jl�%���!��������r(�����������^�E�HʙkxEވ~cUx��I{�F|͠��B���j���y\q1b�*d<$\e(��\Ɉo�Q�k�㚍���B='�T�#�*m1�0�������_=)��e�Ɩ��]�9��|�X`пԲ�S���7d�Z��
��I/��+࡯��^H���@�RJ���KM�q	
��T	u�L�䷚�
�|ǅ//�tg��TN}�9z�d}�髻�9���7�I�Qޥ��r����婣�&Lx7~�Xҋ��#W ��Q	t�gIgVDO��P���'LVGx��Т��,Fu�O�k<���'$�n��^�u���l`�����W��fo�L�L�8梻����7
�m֛�"LŽR[<����	a���=|ƕ��u���ъ#��	�>o3��O����I��z˩�)�-W�Z5��}Cq�I�G��M8bp�ҥf���%YC,��[Ejߚ�b>��=�_��X��*�S9�c(��-��U�a��#�#z�Zr�G�n�J5"�ł�G3E���23�	�����ˡ���I����4�l�����l��.X��v�'h6�Ԓ��t���{���q4\�
{<~����T��Y�8�H�s5gm�T؅	����'�>�6���g�FX*�s�z8�4�C�kR��4a����O&6�w��W��]-�Va9�Q���آ.�{,b��S9K˫��[XJ�*�. �CR$���g�hF�,Q���?�X�nd՗��ej���!fW&�-�okN�6�1�)�wzy�O����LH���MS��$�e��5f��lO:�9�}����P�[LFĹ)Bݑ;�H�����hcR�bo0��G��;��5_���Ԍ��_��yZGO�S)�����|�U:ZC;(k�euI���#!6�����mJ�fU;ܻS�t%RY�/�5��pM�U��`�
��_̾�DQ��O�n53��`T�p�	 p�Cc�����X��$L��־�ߐ�@8�V>^�\�u�̤� v�殛��I1�&�Y��i�VE�i5��`f����ol��Ij��n�����e���x`���Ժ�Ns��u$���"н�=��L������r�F�ҲK9�����3:U���7~OZ��ٯ�΍?�x����y�^��ɸ�w�M�n��}�Ƿw�s����Z���i���&��&N9ab�#Խ���Qȳ��d�50�x�;� MPI+jNE}��7������O� ��������H��(k���C���.j�������ݺ^n�"�Z���f�w{�,o�{1���[�}�n���$�>�q�\KT����~'��*1F������]i���0|�L&��I�6���X�AUB~>�{^0���I�4Z�f��J����N�R�L,�����K�f�
P�gx��E��L7o���yw�C:_��=s�ŗ��ՙ�=u��
_��Ay��}���`��G)�����c�q{�*���<���Խ���͵8��)��i{�^y��l��܏�P#��8 �«4���f������������X��<7��M��f}=�"��}?�J'��!M�G�K)k���&&Ә�>1&�B�cd�l�g�gL#o�c�+kN���S��=�=���
��"$��-^ dz�a����O����@T����i3L��R�=��I9�ҝ:����}��C�ƫ�}��}�a���EU�G?]�77tN��dO���H�:��E�_;�lzB�<��̝�o�%�ߟ�~~��_j�d��|^��Һ�!�g���c��s�EBϥyN-4'�d��V���o"j�c���y>��ڄ���\���ޣ�ޝ?-A��6ۇfkf���"4�ף�б/��o�%����Mn��H+��,@[�K�ɵ��z��B7
�NjLsn~�u]3���Cb�@F���Ɋ(�,fs����Q�P?%LG�ƥڏR�1�O�m�B�2���o&�d{����ܤ�?�����]9�hXaص�E��o=?i}3L(��,zǸ�{3���D�U�fhBM�|wO4^�4cH�Y�1�����M����N%v�Ix���0!}.s�"�$"t:$Yi���{Q@!+
�@I10f����6:�\�v"�~�JȅQr�lET_��6X0��������\�5)�/�,B`+���8��B�	F"^�]ܥ��}�E�#����m�O��.��hL@&^qHX�H?"T4j�&83=�^��@%E�1������en���Q�D��=��� �������iB#t�b�e���xq����V(ȝv�ښ �HmȻ�*�5�nЈ�ͥ��y[]k ��h��KP읞):�j5��x�g�<�TQ�:7��J?|��b��)g���f!�:�EV{��t�:ئ��)�K�oD�;�8-w_���v;��I�i����x-����{�#J̥C��)��n*��{8���vo��<7,�Zٷ-�8ª E�W�
�����s������R ӭ1c��0pc?�D	]3�yE�wļ����tK�B�����~�w�� ��%/�pc�L��������ʱ��O7u���1�Q�����B��>�Z�3�Ӿ��A�4�ĩ��;�2J,�ݖ,�ʻe|�>�f�:����9�F�*����A�҆�4�D�&��
9�9�"������,��y:SQ���F���.RC�/~u+�" �q�3X6���S?>�A�.W�����4����"���?t�:T��d���&���:5���n.Q�#��$*�?��F�Q��n#��� \6�HcH5��?�t'	�W�Xh�~�d0i��ɖ�e5�\�A8�Abݲ�碮x��X�0B��݌�1*�7��w�@��o�s9���A�/V�N��k�W�����������N��/̔�&��m�>�;�_ՌI��׶�i�D��ӫC�D�{���bW4�5�PG�#H�~	�W��)��*��\ DbDR�R��'�
�l`5�MH�I�b�2x�Wʕ|,�'��b��O��Q�ᘫ��Htvf\�6�r""!�Ų��!/�GsQh��Cۍ,�8_�(ļ[��}���fR���m��<���e��,�?�Jz�<c�K��y�*��4V<��X.D�t0��=X��0�)�߾��Ĝ!XWh��b��׮;e�,k��5���1�-2������M*dH���_��t�����)vY��rl� 4@˿4���ҁg���;.n�Ԙ��u���b�Ƅ�C�|\�$�y:;pq�\#4%j1g�-�+�O��z!NY��䯒���)w���Ƿ�нa/�m���-Pp��W2_;��j�#<�� G*bH"��.�@(�X���/�?��s��ž�����侗�]�/�����R�\&i�d�aX{D&�ܙt,�ᴣ�:����X�aj����ԾRk�6e��T�4��vp�N�O�B|12�B�#�t�~�lh�Ҵk
L���Tj�p}�8#��@�{�]a���u|8�`��fJZ*�� �#�C��C�����ԔJ�V�D�G{����T��	��R�� ��@_xO0u��}�U?\�ҁ8,���ӓ��"�E���,��/D��ѫ����q��]3��	� ����2�����h��/ ���I" C�
bR��r�����ƫ���?P	���o�讣-��XzQ0�Z�I�c;I!��<��H�;��Rv�����?hS���*o�	�z��
]�k&lOBG�� $��]K�	�B���	$�3\L��e�bǂ_S�5��.�*��*�2}>%�!�k�H�yFAy1~d"J��rsE��f�b��X��9�o޹d7![��O�����5���#����/v�ry��v��E�������2�+�ə��� ��D#����w����x�4�T��*+��Z�~�p�^V�z'���H�����9�,����7������ �֨��T�$�����=b2���m�sM
_~�e�'q�~��A^	j�sL���S�®;��i�vmYMU�JP�R�� ����:RVnB{�A�bًSR�m�id
y�˚�0�K�x^ڮ�M��Zx�	�4���32eM��]/��A��8R����E���׮��q��,��$��}A���pvo�)8~YL�"N���B����a��I��h�&�rق����Y��|Ƴlg��K!� �e��r��BJQN�7?~��^���hn��w�])j�.�c�A/LdV�*��4?�2B4�4��� &+����Yx�<|"�J�`Y^\9��]n��vW��@U���G#��+ޅ3O�ۙԥI*lwb���t�Z�q���ҁ��Y@>Z�w)qU<NMח�y�����YۄT�Zq��[�I	�d�*n�b��5�K�b�,S� 
#X�e�vr��{��qd��4��pˉ�e��wq��Z#4U%<d}C���4��G	A1����$Ғ��e6ܨՊg��R��bx����HwEH%��5R�&�I��k�NdvW�7`qUh[:���FH�2Ac���@�6[j4����	��25�����C�F$� �?��.��$5jYOD�PvH{��Y��ի����"�;�aR�jڕ�bN�
��3T���}AV9��-���7�8e-V"�00Bc�hI��ƫj�Y�;g���(t���u�r%L
��y�#�<N�~56��a������ShSњ�Zׅgi�W���M�]�J��
��c�&!�e��_�`�P�Zۚ�pd�M^������FUw)k�54�T��@�̲�g�ˆ������IY:�`3X�b�mN�ٺ�Wݲ���yՀ�H+HB:�G)*ZjC[�ۢ��=`	��ֽP^��H0�|��>g���N��\c�9�\k�g�s�SUV� F �T��i�Ί�D���ƿ�����K15�P!p�iv�UL�TH����H������NkD�^|�
+)�/����o�$r
n��0�;�`U���G��/
���d�D�7�j;]�����#��Tx�.�]#�vM�$ȫmG��
�n�F�DH$��c�ep��De��v,��x�"��|qS��ߑ�fNd��U]�<\������Xm�HũD��jmKݍAA�'0A?���/,)�ډjq*ْ~j�����?���Fi`����0:���F7�^�!�
�Z��gȕ�&3P�8J��TbcS�ｇ���]���ʁL|�G�'K�ٲ<�-�iv�6�� G*o	�.����Ŭܟ�v�E��,�E���OM_ٕ@�eG��3��@ h�	����QU���?{�����MoQ�߽��O�>Ļo`گ%����#��c�ro��>EV�=�W:����oh4S�;̖�5�-(ע=��bFP9>[�$��	R���oGD�}1�b:%��e�L��H�ǗHU�gF��]�h�U�/�l���Ya��AX�!��ʝ��$hi_b
8l
iZ���]��<�%�0A��S�w��hV"S\U%;mx�F-V�r�轰�)�� �<P��a �!�̏�� �1�� b �ZCRCj�Z
,��ڲ��e�T"�R�P�U%(��-���zDx8D~�����`-|��C����2ć���ګT嶩��❶8d�p��iZ�L=ah*�0���_�"�MU��mG�$�֒&�K�7I�:R�^��<����`����< ��A��=��	=	y��X0����ګj5t�����dDm���i���U�_�&���7\%8�݋���� ��34M�8��h� %�nm`����S��1.��ɧo�߹�b4���]�՚N�FP�q���[ǿ)A;)�&(d4ۑ�TW��#@�wJ� )[�<�R
MŻ_��v� R������KiS�ZF��
�Vw��4��!���²du4 ��p .%�ﰪj/���`4��r����]��|�������d�j�Kf�[%_��3�!͆�u!����S�*���v��.{u8���*�<$/H�#��(����z�����m��iv��5��>M�b�@q7Nx��,�K`B�>A�BtڣFm�2�\\jh<-���hb�S��M
G\@�Q���fP��+�vX�p8�׆7�� oTG$v�|�-�گhP7?O�l.�F�c ��*)7��7�sv��^���0�
M�[Uwc�O�����dy���DS�/��؆�o/J��ሻ[t�omz��\9e �v��̯��Ҥ@��*%��|}HM��BOcd���y��]�t>]4'�@�*�v�7�9)��)�4<�|��|^p�B�<������ɩ1����e);4 �i�/3-�����5���L��9m���m_lS���<��<��4qqfNc��D̃\��qPa \`٨��<�bFS�� ?[�Rj��&�?��h�i�8M���Z%@����ߴR��D�-�j+�T5�Ydޅp��
nHK]�J���i�9O�R@f;����!�$�b�ž�<��%[Ӂ�S��ɋ[�T����Q�h�����.��~�	��rQwTd^��)�ϔ�g�� ���j�8�Z�|חŴM�N-�!��db�<���L�mJ��xx�
���pKٙ,��Op#4̘p�65Y
<�{@0>Z�]��T
���HL�	;��	�s��P�\V9����N"��P��/����y���O�ݺ��"��ׅ��.R�	B���,<$ZH
˦��"��ʛ'����A��]-b�H����*�#�w�q"j��� I�*�"�Ym�z _ �R�u)�B[�����*�5�Z̔]��.��w�;P��8�g��!�i�@���llKց7�彋xCNY#:M[a���/]Yx}+w�gO��JR@hi����i���*F��*�����[�U��Ѻ.�Z���Ƭ�� MyU�9q��j�-���"X&�v��*Ua�C�tF��噭�J�2_�F�w	<'�-+��NO	����Zͩ������]*��r|L>D�X� �R��O9� p�N�����Tm#j��O��n#�*�T-b&�ڵ*"���c�{� $�.���jG
��T-+ı���k�p�b��m$�J ���G���+O����8UH��{y���T� ��#;�fh0�����X*q�Ve��*�hpY���!Wg�J�[
B*WY�+�WP���>C �	W(&���e��1c��[-�T
��3���$�I��K6Bj���V���MN����&wϗ�r˚��g[n�)A����D-�N�IZ��!�� �ecB���}d��i/J�e�#Y�@q�8�0Yq�f�!�@!P��&�ltK5�2�Re��k��!L�4�!)X
+�p�}��<�F�^�>>����G�w�=�����ǡ���h!ӑ��x�:�J��b�����{��m�U�1>N�I
�����j�����(d�th�0�)�\�@�8D� �!�-MKG�apܮ��������xс ��t��(������.725�U����R�Sy�"K���j�i�"��:4"����n9��Dv8�3����`jbY��@��`U�7�X��L�ZF�Y�)��S|�fG#��D�*.�Gf�ŗƃR���G�B�B ���u�T��lr�,M���;[ޒ�PFh�o�v��Xvi���p Zjb�Dx�Jmj[��Y�(�/f	�⭥&%���R܄�2�ƑTD�#`����L��Fi&��d-/�� ���R�`��*�X�؇:�w�>��*{�yg�Wr����%"��hr��V�w:b�������%��}����Bǻ��hZw3xz"yQ��������\q%d��s �[V�g!�bd�x
�t6%���K����^����Hl}�fxj~Ty���bp��+_����햮�#9Zԑ��)eY�g�V?�A��[��� ³�Fy�O;WQ�%p��(�"(8�F��-��Dld?��B��1�x-����L�c���w�p��3mM/�sD:�i6{��\k&�����Hʄ�j�r� '�o�o���@U����!���EM
L�?���x(G��i����v� ��4��;M�F�.��P����i�A�)�k`*�A�,�0R����K���NB� ����ؤf��1)��S9�b43C��!��<�d�c6����wQ�J_!_�a,w�D�,�)k�X�4�8NY]ڠTMP��{d#�T�(����� G_pǂ���(�/�� Um�ꢖ,&B���u�qr[���������ݐ�k~�fp���O����M�`.��������cD�\���=�����D!�ׯ_� c�%�3����������)�X�B:&1�� P-�ؾz�i��Jʏ���Ra�Z�%>>�4?��RbT�4��4���q�������˗/M��n#5�#ű/�Nh*����R�GcG�7i���Y�l����;Ng+� 2C];�f6���I��t&�~�$Eͅ���7����J1R>�f�u�Z�!N��ˤ5�?���R4���!1y8G��d-�fXa��j�!x|�p�<���&e)���	Ǳ�/�v��M��YLǒ��R�fN���\Sg�ڹI��wԮ��ۑ[
�6�f3��T����Ȑp�Yw�Sse�����RH�����%&o�
 �֑�%�"BH�S����<В��Kx�}��f�`j��BjI�)Y������t��Dڈ4�c�j�T�X�HC�o8�0SP��]"�(ڡQ��񢅐�^b)����� K9���촓m/!�*\ߐ8q�4�l#�e��s%�ъy���.q�Є�S�����Rw�O�Zo0�����0<��!L�Da�ls�"X\9rARN��!3Kd�{!�x&�#/nL���n �Ab���<q����ʛ�B��,SV�N f4-@F��������m qV�U-�]�ŐMԽ�i�h3G�@60(��ZRh�@�-�{�R
�-�&��������5%"���kB1��{F9��F����a
����c�&aU�e�$����}�!4-ַ�j��ŧ�jddY��OD�/k��.��LҦ���k��S|?�:ֈ�D0ǫK�,`R��y��㫍c)���$���y�#Tn ~ � ͖�]�B6����ve�k-�l����偲�̓Y>�汼�=-��J���T;B�6�8�.bx� ��D��]�ī��@�0+�X���D��[��v%�!-�lNUY��~�	�DUSU��*c@�M'X	���:F��o���.���!�,)�M9AL���i ��l��U�%^�i
�&@��?чo���Y���	 M�� �)�,�5>2�*o��b�*	�+�'��}/@�hbc�ҁl ��B]����Jj�/˪m~�K�-������L��Bc4*���A�P�Ѩ�k�9���P�rS�n�wn�����q�酰�T{`�y����	Ǆ;�vdN���&TR��I��P_~L]V��|P)"����}�٥DK)�i�.��3��d6������D-%@��6B�օ~:���DN')1�I\֘�C�sݽT1 ī:LU���w�	ڈ�樽��h"�9���oN����;����K 12���`JEh<�7��)������>Sp��bqK{�>�篐���j6���ֈx��-��>����:4�	&�\����EÏpm�<u�;[�e��6��4�m�B4�)#8����@V;�������!>�TC�V�� � �D
��\!p�)P��E֦�m�5-/��*K�Hw-�fZ�[n�p�N�ɻ�G�j�b"�����@�n����m���i���6҂j;p��p�m���Z/�駀l�b8���b!�
B,qXM-�����D�����p"m_P��_ �d��w����NY0���Rs�L���&�R#q�\�>����M_Y�h
_�{��p�x@�ś�҇��)    IDAT�@�7I��gϞ�DF��F��w������vb8�d�6��aJ���4jY�*��z�9�3A&��,bm�5�;�[.e*��O����΃Η������yAm���-mc*�5�q����� �g��)�y-!�)4�f�,�J��v�(�J1�<�K�j�A`�Z�H4</���M�MЉH��˶��qR�u�{���o|�@Y"���P@X�C�pן�|S���b48O�񩹢N��-�Y_�������w�<s)��K0��Qp�A�g��������G?��{�a�����)�~"�կ~�����x�����q;2ï�k�*��RSfr^�](l����kx#�|t&pޮ�C�lxG�>�襊!(�����94U���0�v�Y�f�Ȣ�55��!8��J,�Zk�@
(H�T]����Řj��gG��;0}A8�R͠<���@^V!>�"�b�>�mt�����9�H!'��[���RG`Ӣ5�ZW������ѥoȤ�~�>J�Q��x�r+�jj�+dݟ�pw�;��&�y��I~�߸X�͏�کr�w�I���`Dh��H!����R�x֙��Z�R��}�n<{�$�d�j�`�:�����_��C�Tf�"51\���>�Դ�	�LM�Qu$���~y�}��o'��;��N]�ׯ_+��.���&p���|읅 諩^&��w]�Ut��{�8+�5�P��|pĺ��&�#W�6�����ϴ8tx�'���LY��4|R��^�ctd�,���C=�	V�ђ��CR�YF�B  Ϛ��,���4�Z�e�]�C���S���d;�p�����!�h`M}���<�r��>�T��x�t2:ʕ�e�� ��5��!��O�Җ��<�8vD�G�H�2�#�&���{�`�������ؐ;�a 5-06rHAwQ�5�0�!�8�4��bM�+ 7$0��	�D��qA,q,�w)�F+�*2o ~��6�T'V��EUouI��7	�,�8���S��W6�`�e��RxZ=~ �#%�Q�B|U�(�(��A� 8��t��G���#y}�����#m9&ߜ[�Y�:&��&�`�N�}U����^�ni�h��q�m'�z5��U��/KdA�X��w�-����<[����+�p�Uߤt�1DP#�G��SU(n�>����=
)Y#ח`4��1�J��5P�,F3Lxj�͵$LY*�J�M�ܖ-�Z$�	\;K��T���؄ 3	Z�5*ŧFpU�@&�TP�����}l)"�� �q;�L��	��B�F�ϳ{
��BA|���U����pK�-�ZK��|�FE����_an�dUբ�i�bx-��yx��r1�{X�F��*�.�Z1)~�W"6@�@�* �u޲B>>D�+䩙��f���L�#���l��ѐ)�ΚZ��(^3�������D�ɕ��]�/E�ձ�! �*��Y�J.VRU�2��u��x��9�UE0B�B��zA�n�:�f��^�B��1�T��\MjoZ"W�f��ym���kG���OD�r�v�t�Z���r�:�M�l�4ʥ�Ȳ<�u�G`9f-�+o�J���?~v �)p-��_J�O-B8Z6�v4)�C�V(��rj���a%�[�b�ͪUBВ7�@Ǯ����d�j�I�:�L��j{�J���[����N&)��b8d���a	�yK �>��� .hkkl#�b��)4pd1Y����b������N�2�1p�i��F�F������,�Z��F���3�J�(�iFj�ha���(t�d���<�j�̖�S63Nc���o����C�w�z�b��JZf�1M���A��)U���^S�{��񗲦�=ҷL�T���6-�C�9�@�J�[��*)�����C��:�]k��O�{~�@#��x{K�m��0�c�v��)���p�8Nƫ3�^Fa���|��?�Ñ2m��ɷK���"�;�]M�ᥔ�L�mU5E� l�� ���D>��vq����R
-�N /U���K� ��gT��D���R��Y��K!� [9MK�#�
G_ �*j�	^u�i��tq;��1eS$�'�R���� ���啤�߱Tx�\�^��X�ܻ��,}V�k�Ɖ���ZJ�����^�55N�X^�f��.�3~"�&q�f�q���ɦJ�����^�J)�녩��O=o��z��;�hvoP��jڻ\L���>��M��ՋO��v�m�)u�S�%o)P�&�=�H�*�A���zX�y���k�~� P�aBl�Q�)�/�߹��5{����U:�mhIi5%]�ƒ�ȐmOyK�9�x��@4A"�h����S�7�3��@�[��@������-e���QF ft ��qj
Iپ^n?����D�J)qb���$5���A��"�-q,�����7j{�$(�%�3�Bܲ�d�ַ���/~��T������3�u}��>�C�����#?�|Ea���gϞ�T����T_4���B�l�.М�y�	ڏISi�Iʒ���� #���`�1���DS��A����ɸvb_�؂�qߑ�h�8NM�)���B�g�̣
MI����
�ϋ���(څ贋�y4�q�d-�)��#eٖM�� ���Q#c*��a��1�C`�Ru)lU
 L�SOVPk����X��o##����Ȋ�?N��e�B�3W	�-�M����d�w�[­�F�q�2�h���솱�˺�|y�C�Ph���T�����W����ڮ���jN��.|d����ܭ�fH��4��W��y��¯�8��� �����Ĵ/]��v�
UY�M�r�����>�8�:�1݉��v�Ta*��B�]_�@��K/�.��iG�@��ِ/^�P���h 1�)Kd�1��Y]�6��ct�t�;|3 �\�r��;́���Q����I�,��)QHb����#/�V�uQn�F��(�,%Ap�ʁR��ɒ*n�@��]�f����T�3\U�j�K%�)SȨ�-��N��a�l�.�;�s�1vE�;������4eD�"�<pq�<���I�f�a)]�B�,o�H�eAG!�UΤL�KUhg�K4%��ul�B�(�>��v�͜�T��FJ^v�A�������K�B���R�+�<��m�T��m�R`I�	*4��	�UY�I
(fb��;�x<�u�� W�?B�-�f^S�Xm��~�[ʊ)x�t��(�,?�*҄��l��E��tz������W�,~�ᝏ�t\�;Y���i�U�{],ӄ�)@�����kײ����I��w2�}K�l/5E`�c�7M� �VU�:��8�yǵ�)TH���y�M(�B�(1�3�0_I�1��W8���V��v! ˳��l����H5OM[��\FS� �ߎ�K�OG/K^U;m%긽[bҩD��B�ȋ�eSNj���h�@�EY1C�����y��5^�t�C���*du�T2~R��LsY}w�8�# o�d����-ͯq�b�uO�t���D���<�*�j��A�Z�"�!FmK:1+��n��Ph)�o�hR
��%�|pYURuo�vM�b���	W�,%�  ���'m���)T�x"1!���p�󵶜��Z�W�_m:���46�tx��]\�٬%M��8-;@��)n��4!)q)ޒ�D�`�7LcT+��i#��|{_d1e�jc�C��@� �TU�	�D���x����#�e@�ℨR��NǸ� ���4�v'��
b�Es���k�!bU�V@���k�8��)@K�R��Z��|�o���ʛJ�,K�3��"1�Xc����%XS����	�]��L�o���B�bv�.h �}�.�q)4?oZ��<�����!81�#��Б�,��_L���ê.x�h��n ��Snʫ%��q<�)�#0'~�N[��9�<8����F6������E��S�Ɔ�m0�'«�Sߤ�ێ7ou��� �lv!Ii���	��j�pW�~�����ыm�*�9-)��I�nBoK~��_���F;>�^�J�B%R���iMe$��P��}҉!h�u�)d�s�NϫZ/�|�?m�f���X��]�O�����~�f����˿|�����6����?�o�޳9�?_�;J��%���m�^(Q��N�{V�t�FY[`h�tJbYˆ,!N��-��RzA�|����K�;.�2
8
��h8jq��ӏ��&e)�,�llYxF�R֕���y��ւj
��^�Y8�npˉ$�	�N��2�|��U	�e:�X�S�c�d[�eJ�ű}KD�������K6/b�D�%#+ַ8f]�,e-�r�V5��촹�-��R,K��6pH�R� �
�6����ĻӞ���v�J�����?|�c���������~*5��Z��g�^�zG���K�~=7jg��Z��Tط6��]'�=u\/÷�n`sF�9P� ��6d|1��D����9��g]��T!=�!J,M�3��izBz{����?�)�}��}�m˩���g$z�
GHcA3
u�Ɗ�A�d;e)��K�e�T3��14�
��[�� �Z���A�QG��y����*L:H�E�3"�KV�L���ު{�FAf�p1�iz�L�sw�h���lU�6�Z�ZW�Y�����pJϞ=�}��E��7����~��9���)/�#�}?�|�����` ��ش_���}㧠C��ڑY��u۹�h��t�թ�'�HR��cZ�Qe�,ED���BlP`0�@h/�-J��d(���z��L�*�^hNG�'�{ׂ�1:s�� ��2ys�ԝ���xjY�ʆ��E0s�R�Ē՗� $�6��:45�C�\/�*YK`�̖�0y����)����!�Eْg�zi���y�;��K����v�[7��L��.�9�=��K��,z�!ݍ<A�~3�4�[E/M���&��R��=���S�;���L��_�|~�������gwD�|��cn�t��_��D;_@���P9��f	:C�r�Ԣ�7U&FCPhkMk��?�q�6�߀y{<�����gWk;�0��˜vmB8s��N�����8��`}��'����v������t~	p���%"�Db�6��P���޹I�l������H�9��;(�~��I"�8�j6⤘@����Af�HdY`� ��;[K�Aс3*D��c�Y�:()�t�R���*nID�8Y�Ő�!�F0>M#��r���+qE�O>��F�g86E�-�Y!�(����N�s��B#En<��R��fv��6�~y�t�
�<�����i���
��)F�@(@Đq�4�J	�b�{��m�jGC.{�k��:�u!I_-��h<�%�#�%\<� r�w�~Gv3@��	�MΔ�
�p:7��(����J�(	_9�v� ,A8xrOVUXK��������l�|8�m���M߉Y���<��1u�n�v��ǰ����)d�>�ʋU�K�S�����ɊyHAZD�R��!����Ac��@K��V-&D܇z[���*�l/|�"��.�t�@��nG��Z)V!3��Q]0��,Vh�71/W>Mx)7�'R-������\/A;R�/F�ww�q L��\n�J&e)+�&K��	T%f�
�e��Z�
95^�I����T^��p�rq�M���Z���$�$X n*�]����X�{a���O�.� BX���]�4w��)涠�%��q�������pd%�F3���S���r���c�_
a-Ҭ�OY��-��7�T.僐N[�v&ĩ�/��Զ��ֶ�Ē5I�UB��yR�-��TEH��G!K!���@
�^ ��Y6�
.�>H�"�U���V4<SE0��<��)� [Pʒ�q������e�qd�XaU���)�lx'��Z�Љ�;�t���qR��4�)4�81�&O*e��-�h<�3	i�Ū-K�8�j$ٮv>��qU5����y"͓�p"lT�&�l%4�OM,�/˧ u�9Sh�) �3��SL�l}q��L��*H"!K	2��ES�(���;ɔծ�v�L��?j�-�$�K�ߞ�+�G�W1ok�!� ��p�=C�UK3��w,@�I��+`� ���"�M"6���z�7���Zބ)#h���,x
�d���W��s�aJ0qJ�ۅMk�5?%�ZH�m.�EjyK�p�2P��`OJ	e�>�)2)'&���7'��*-1��\�|����h�� ��#��W��H�( �M����!/.l��v��"�\S1��7-�ޱ4[L��-��\� ޖ��m�?���潐?��}��*w&�R�/j��nG��^��������[��/_X���8�����MU�&	�+�t��T����-[���B�8�H6$?��p�uWXw�,�)Og[+��_U"i�\#��n�8���ٱ�h�%Na�t���(+ 8�:j��������AKM!���4c���>=Ċ�J�jU�Yy�bx><�t�d�SgNo��;�w�RēJSa����G�<�y�RR�.���^|�}��S�Xg�j��Z&��c>�8>�>�^�A��sc|�i�ʣ�4������3�yF��o�U�����3���Q�-�w�ޯzڈ{�l �i�C��%�Twx���\/��R��kgZ�#鋑ݺ|�S)R1�#�H�TY�.D�	��2S���<���cTu�����	O��ʊ1�4czC,Ih@�4�b�H�-ͱSk��L��2]T�w�,B�l�.-����G���^�H5O�wU�k
a�R(�k-��Ѻ���G���g~qwf߯h���Fw*�[��Ԕ��� j5�U��o8Ժr.�����C�U�F��4�O��-׈������F��Ї�T�:��ig0�p:@:b��0f?\���/���rGg�,��[�K���R
Ak�P��A]�x��R߳�� �vO�07U�P�c?���ptqb��x��8Z0�UЁ[��#+lB���8��u\�Ȓը^�@( "[�j�A�m�dk��]L`1�iY�f
��wi�*Ą�]exR���2��nx��-Ř�-�]%�Q	��C�0��Q70��/���Z��'E��a��F޵�ۈ+��HwEߌ���<�Z��,��i��Pp�}M��3�{�����2��:��ER(��^Ҕ��&�#��F��)R�tt�#���QkT4�_�C�8P2e�2���hN��/�b�5p�YGJ��R�fy")�N�8{Դ�fS��ܱ��D�IS��b$�ԹxW/[��I��P�����۵먩�Z(1�	��R@�׾ph*q�V�&�q�3��54N�������"�R��2����Q������3ĔjHxUѴ�� P�~3�JV� ���v!(�PJ���,��X����]l��N	69�0�х�$�����5O�TB�$��gR��T7�ZFǴ�UC����턈IV�W{g�d��N���[�+W��*D�ʀ[.�.)|���H�`HU�b�������+�S�Gf�R̲�)7 D�5� g�!���x�bd~415��,�`c�|�/�CIv4M
8>z��Z�{�^��R���*�4FU��������
�*�*MM�;�8���e-���<�|�vg�-yK>582DU�ʓMMv��Ä�g���5В�*|K�L`�(��@��o����~��D;�� �$'ҽ��Z����7 AdH�X*B�o���l�D�L!_ӝՕ���S�I�mj��-Y'@d�
S`ȫ�lA�;�����#�w���Z(����5�,�TdHٚ&���Y��T�oIA��!4F}��\��O�^+�Ɉ���L����bZv�jg��AOa���Z�F
!����dM�)�r�!��pK��D��{"J�tIm�}^�"ׂ��z:���H�<�\��	n���X��PI��Q��hę���N5�2M��ZKYAHY���eRZ쓂�2)&"W20�cǩu>~��BdYq�lx�dWX�{a%���t�    IDATm�iB����i�A�M�}ᰚ
��;�@e
�޺T�gU��5�,����EԀ�C�Q�W�P��l|����Qծ���^x����D"�ˢ�+k	�)��^	��n�m��M���_�%���Ru�y�𥢉�MUG4���@�Z�������EaSI�/�OnoS���S����F��O6�*��+�� �N1�ex��
p��y��_V\I���d�'e��g&~�t���~�{����'?�OȚ6'_�@��S֏��i����Q}~�-ᬫ\a �HY����5E��ڎS��a�(�4����,q-";���0D�������1���mP@hrA�����?����y�R�h�g�;O��#�r����VS �p ���^4U"�������u���+�����B
R
�LAwS	x��$�<~��͆���8Z4���-�^U15�
-3���>����S�^q��o�%_�?��K����gϞ��Y𶄸�7����fFd���	����}�i*)K��[�PS�⺛Ͳ�QX��j�������t"�*�#x��J,C���Ua�)���r��K�5��C��!8"K���(d���b`%f���"�b"������	BXR��d�p��#�Cv	�@�!�|�M%��P�x�Z���#D��x�骆�2?Y�ā�]S��c-Z�������#��`�]��D�#4	���C#��Ip�)��'��w�h����B��Ӈ���O� �kU��/������p������?��O���Ok|"�!+��'#�'�ǔ��E�7ؼ���*�V�ӍG�f)Lʒ'(8q}R�÷G�E��B���۬�CX'�����$}�~����Ʈ���?�K���)qG�V������[Q�d��Sҁ
(2BL�����y��@�JE6r%�`�!�� �Z%1��8LR�4�G͒���r�h;��*�UT(�PR��6%��9�){�S�O�ɺW޼yqJ�7�̈́LJ�]�L�hp��a�Q�ie�Te��ͳK�dM�}���b��%��@t�/��m�`6H
�+̾m�L\z�ᛍ>��Xk�,;1R�
mG�A�6ϟ?�o���.�Yd
����li/�1-��<}�R�KbY%�;Iq[�C�u1	�%M��R�N�7��&�H	f��@p����ȓ��J�H�)kqubI*�bY�6r�Ѥ�5��Z%�+���Է�U(��<8�t�&4�Wn�8�B�tT�W8e%bð
}����M��=��Ӎ���'��/��� ~3��g����K!��g�oc�dZ�_``�+����w{Ӂ��� �G�0k�A7���� D@�����(5�9� w���"�o�LS�Mh#F2d�@���� �d���8�b:�2Y�B�@#��̯��	ڬQݖ��8R��*�1�'����٠F�b�����|"h$GD\Sq��d�"�A����5���%o��G�az��b$�'"���ޕ��P;*��HY�N�.\��3Hw��\dY���H��鈙X9�Z%vC��L��G��y":��NR�C�y���X-⨂�B�����>)S%"h)`.�s4����H���x��4̓��!��u����Z��H,@su�@��Ԃ�1>��@��.o�&GN��КY ˇgp3����A�+S������A��%+��[�W(K*P܄#��()� ��l��V��Z�(H3�J�d��X��W��\q���*}�+��Tݽ��)KM�^�� �H��N�[*��2~㉝*~`:[�����Q"H��R�	Õ�>)�;�5�֎�"���g�ݨ�F�.1���c�������%���u�(T��6�
�HMȀ<��ZAʘ���l�:VR�#q3`�<��'���4rU�h�)��e�<%�qxK���8)@Ҕ�QM�@�
^*�4�C�t�y:IA�-)��!����H!��+��B]�u!S�����H�$A�*x�b��H��N����� u�n��S��+qxL)1p��4
G�)/��F�t����`��E�W��C:.�^�S�y̻�U��m�̓����w#�̥ �`��OGG�/e�<�i�	Q2x
D�X��7��wq�����es�'����K�J�/r/�	W[y>����؎�I�b�!(,^�AA�;�]�6��4UU	��z�����RL��/�ǭX��v��#n����TɊ���&�g��eiJA�c�J�YS%�>Dv4��u�������h#��<���e�����bx�e?� jį�tj'�+O.������R�Ka��@q���!]?�1���Z$ŧ���#H�T>}d� �::���NG����� ��χb^���-ő�[�y�PI�X�{��y�����!)q��X�.��)y
�e�X��c�J�!�������#R�v�d�h��ċ}��r}'菸�t�v�qH:	6���q,���c*���X2x�D���B��FU�_{D0'Y�
�_��͓H�D���7 O�^���@�S��w&� �BG�Q���^� ��Q���/�ຄ�j��f� N
�H��Y�=h{5a`1A��7O�0yVj�d�\�%�kC�@�ҷ�RZ�f��i'` Ga dK�
I	�?��t��~�.o?Ď�kq}��0ʛG�lȺ�������_�����wB�Sr,�1��;3(���_��[S���tM�̜�6\�R`���L�lU�w�Xr�i�-Ɏf�,#�Ѯ��aRl�B�BqZ��ŚV^�m�=:�ʧ�8r:��Ŕr�b�� [�K`��/7��%��\�}ښ���9�q*�kG��J�i��
���͐���j��'e�, Xy���y�T8ߜR��ײ�
ۈ�@
?�%�S�o���)�d�r�w����<Y�n%u_	)�	"�cS&�#��5JA��'����Q�R�L?���������`����,M���;�������?��O1�={�u�L�U9;ꗉ�7ޕy<3��ޖ�B`7����nKU	�y;�9C!�4)��J,+)�r���-먁�#��|��ҫiG�}��"�O�J	ir*B�S�@���oJ��R)%pH��e:@s�y�l�FT^JW���� ���)LD4�I�	A� 1�X��b�D���jѐ��~srR@U�~�:;�g0���� Ԣ��B�|R���^�Fxc˪e��v�՚	���F��_x�]��_\8�h��y��63���}�k�`��\h?�������l�S`:}�џ��g}?����_�;��fCv�8ߕ�)����l���`�s�c*��592�R�2ɚb3S��G����V"C�)�4�������)�B�w��T���q`q���4a��j1��P�Ԯ���b�d��pXy���XU��t};����H�$.+�� �R��g�����	���U���:�������x��0���=�h����粎�Z�닦�!�qo(�d��hbw�]�R"k����{^��u�(����>�#�_D#�#P���x���ׯݖ>Gbg7�7o� �nQ���]��B�"5~�,����|Y������������!�����Z���p���K!K�7�;��1�Z�1ڸ���+c�kS��_a�(l�Ԕ���f)C2�Ȫ��>2;.��뗾���{~^��q42��#֚�]��Ck��2��1)�^\b�����������l���
Kjp���.A��<d����4�!�@f��[��H�J��@�滾h�0��(���ڎ�:�9�)rK4�!:jd	tVNF�ܘr�hZ3�ҙ����07�ח��̅�	60AL�B
��ƷDc><��5���q�!�t( �tJ|�)"���+l�q&�$�]mC��d�"���G�Iٸ]D�i�t�'"�B�f���O�/�a)�A��rq����\�&,8�@���Zc�Bm[�m����u1�e�lG}.�c���\������D�5��Xg�l"�&SX�u ��e7�B1fj�b���� �j5*[��@jf9�>������g��i	eYC�-K�5\�xc�Z�3ٵM�u��15vWC	�U%�7a��~���u�h��X�qg+�,����HUț�Qq�X�N�}�ǿ�jT�H�w�]-˜�M	�oC*�Qkفlkhb��@LR@R���Ch^����J��!$e�
�Z&��?�?�l���N��)b�\(.��Tٺ��h� 8�4�트��I�6��^�����������ȼ�kM��)G�B
��٭J�@U�&����㭻��3$�x��0)`%���-K���6�PНiHd㫲;�q��!�1A��<��"�R��,A��oI�N��q 5
����H3�
T�М)�[�&.B�xR�V\*�� kɫ��gb"|�	����D /��~������T�C��P@P>q��O �$�Z/��5��"�'RGHAlr�&>AH��T��S(� ��B٦������1�K kj��+Oʲ9k'��Ŭ����o�Ϋrn�c*L_	��/p�R ����I6�C6�J��ͶM��9]���ul������"B��[3K�Tş~W�UK#5�8rW�w�v�ӲZL��Z`�=���|������+ិ�5rVh�Y�dś����� �_7<�� ����^w�}Ge��v��X����Ѳ��]>A��8B#[R���|3��Љ�D1�Z�]��'�&/�w �fPK*�J��1����8���uKU[k��ǲ?�!�������yW�a���9����-��q4�%�6�MQ�H�Z|�Z76�%r��{����u(����JM�`|��pf6K��hl��ׯ_���YY��5"�����N��r���^�D�	q�����ya�ͭw_h�Z�
4�Fthz+%�f�����߽T'��J�I�Y�^�CS��U�HUbY� �0�����R��*I�׋Z
]�d�MX��@�.�h��c�����#�d�ĥ��!�U�UU��!�ɲ����^/B�ֲ�SS�����TN�]Eg`{�HR�fNbe-,�` �T�]�#��N-ZN-�/�&��to�t�
|ہ����K�0N�����C��O����d-M"�k-f�2�
}r=|Ὓ����)?�����U~�s�U�e�������_;���=����4��ʻt�g�����{{YGP/]��iQ���%~��<Ȕ��c�4 m��)��LP��I�5&\ �@��D/d3  ��� "�ʑ�9���DG����o��%�+�m�y���@q4��_�
�o"JD
��0!���A�EJ@M�E?���v�8v���O�'SH���U�BW!O�O��}k�焣觔Em|�#[_�MY�!v�
�e�T�'���d9�@���~3�ݚw�,\#7��el�y��t[����]_UD༦@�`G�!���-}����ޏF3���a�Lk�L�����J�������+D�q�;s
@Y�H�!D��f��P����M���	����Z4c�S9��X���f�M��z�jH��R�
�L��BkTd�r)sb���Y�����n4岘q�v�
e!���n�M��2"b��6U"�
"�W(eɛJ0�>�p|���aʋ]h��G����0]5חٝ���G�H�����j�׊`Y�ً/~���)�|����N�ǃ��^����m�{�T��c�k����7*���,Y�t�*���}&�Ψ8���������@��ٳw�}����������}
>Y��A}H�~�ٵv�0I9.��M��òƦLAGG��G�g?��Mu�8v��ً��]:��vV<��6}���9���w�s	Ԛ!)j
��I%�P;U��!kH%����5�b�!�Q��F<N��R�4+�_��ԠI�~��#��6�������}jd���L��O�D�A�a�u�8��.S���R:M(ND���ix�%�Mя�My&�o}#�q �b��mb6��:�R�a
�i��<�f)0O
Nҝ���d�
�U؜)S���Hy[�MU��Mb�2NS	���.��.�[�]���1�*���Z�����ԑ���
G�V��l�R�&�PG>K���*���/��7R�j��y�� 15M-��@G��ި�YU���ј���Z��&��'�p].�s�p�#NU8�n6���<���W�V�j�[��T�YJ�ҿ�
�!�M1I�[�J�E�0H���]�
��`Rj���X�#}=U��e#�Z��
V^���kGZt����;�U5FY�z����#A��G�<��'K��(6C�\H~M�(��5e�eץZ)D�ZFT.��X�$��D�[��I���Nyd� 8��hMRy�D1��&�>}�Q���O0f��#x�n�;GV�[^;
�w>A�f�ֲ9�bU)�����
K�3q41k_�Sk��L�CV( �)!4����
}L\�&�l�5�ׅZ���n�a���i�D�ul0"���Am1pL8��ޓm�xV�Ԧ_*�����ꃦJ�,�Ū J���d|)��wJ��l�<:����$��
bٺ�������T��H�-fcT(��H���:Bj�y�@���U�	)N���U�Tݛ_�%��VwH����<f����9w�-��Q�Q0�
eq��2AȎG\k4)��7��~U.��M�f133C++���SӢ�W"��Lv�I�eY���@˦-��-�XK�KS�m�#L�o������mĒO�G&(��ȚM�kT�݅)P�0�ڝ��X�J	��K�ŌL��?�m`�,>�h�&�e��k�@�!]Nc[�c���׽4�uk�RU�.Y�@wǉCc��	w��0`��1>$C"�D0����-5�����.U�T�[�_J/DG� ��O>���^[��J�7|��yʛa�i4;-5� ]?��_��S9���-�"�Q�5�V�la-�#M"ͬ�!���y�b�i�XJ�b���t����"��v�-e!�b�,A^�I�kʧ~.cђ'�S��!D#j� �&/��5 _��!��y
��e!+���U!NO$�؎�����Ɋ�Z��l>7hS�"ئ���d�q�"��4�8���&��@�.��hb�
f"Ļ
@�Jh-�Ȣ3���#Сi�'WG�}��c�P�����f��/%ZkA
�K"m�w?���m������Y?Y�Gi��g/�9��TI���k�V��t3����%�9�E�4Z����C ���"Xf�΀�.L�e��;\�K�E!�Z^IU�M5e����<���0��ҡ��M[
8-&h �8�O����k'`�T�.�a�v!`�)��v��*�>�[NjF�T�
S.8�@˱Qo��c�	�E'Bq١�N7���� F����|�FM*���oK�X�G.�EI)�挽�^U%n"|�>�*f�μ`e{8x��}��W��;��A�[��|��G^�Dt�$y�<(nܸq��Ϳ��/^�~k��_���,�� �!�4����H1-x���	�ќ����p�!�hL�h��bN������)\گ�J�����^>�뭷|��@<=����}v���~]	OZ'�mLKB�pB�d��!��t�j+�1Y�٧��(a���I|�_k�c2�l &��Uq+�]��Ř����eޝ!nS�]��a��
�B:NF��w�;C�ĝ�D��Z:�/�)"��œ��Mk��2S�ow
;a8qH��)�Ʒ��q{���9p�z��e�.�� "�ל��O�
��R:�(�!�o�����G3�	ӗ�R�̼Z��eJl��IL��?�(�����=RF�7s�XRS��M�����(7 ~�h��J
��*�f�R	$�`Ȳui�d��rY�.b�ʥ�p`��`���@4FͲ��@��G�u:<k��T�@SI��u.J�ё�#+�p�rAA]d� ^;�@4��#h�l�������.���Uvgvs��j���.5�4��˽'�&YF�I�M�MT����߻�B@������a� �B���6BY��7 �/����+����~�A��]c6E��Ǩ��<=>�p#]�~]ߟ���ۑ�<1�LB5    IDAT~����4���{��q�j���C�8�ǎ- �kn#p؋���X�N�͝L�=j툾���y��"���e"f�=���yW�/�:s��rM��ڻﾋ���2��0!=x_\��YU��(��`�(����cw��^C�vxY��|/��f���҅��� �t8e�@"<ñ�|Yd1O�0��
L[�6��bhpK&�q�2A����d�� �ZK)���0�Ҿ�mY���!�)70�9;=�u��uA��Aޭ�/����⫭���M��S"k#:�%���&�5���;�@v�$��4 �l�t���^նT;6d33��Ƈ��ӟT� <q���9������?�/�Z�6��{-��;1~�F�b���6���,h;h��5U2�2^���7<�؀1��j�i�&H*��jm�}Ҵs�р8�c��I�E��a*)����˦�<�a�|�y�Qx`"�K�ӷ{"R�BB ��J!,�mV�Ѐ��z�l��)���g��BU�]ܜ5�v�b��#Rl9w��-�cBq�TSс仲)�E��)0��&���Km�a�k-H<���B �B2�v1�ӷ.h$H�Z8�T�f;��T"Тl��(8[��cz�t��R����l;3Cۑbhp��oɣ�'XR� RA;*3_���e��b�Y�<DP��[�Dp�%�҄��ʊ�XƉ0����w�Z3�u�8�8L��CٖR�fN
ؐ�Ϝ�T�P���B����@|��e3���ř�zM�p|6
�œ����ӌ��l�b��T!d��K��w��X
���|�vJ�}5����S��&.Hp�fY
�֖���0)�>��򉌏�D�
��*�`&\���� ��0Y4A�j���"��;���Tw�:"��#�S�}U�-��
k�˦Ŗ �W����Ip�����J�R �5¤Tu�K��Z���,3 KV�ɔ�G��4��Zq�D.���c;���
y�R8ι.@Aj|�g��0��6_�Ӳ�
��Q\���F�9˚aR|4����"�ִ�L�K[IK,U�kW-0d��A`�s:����F��g�(,闚*Kqd������T�~������
����4-GYa@0������8�R:Uc�� !�1e���	��D�EU�
��\8�&�+O��Z&X`Up
!h��d���a���xs���b�Z�1{'��A��RbdY^�%��#����hꅏ�)�
Tut�,�|8��:dLY?�v�[R����͆�5�����,_̔�GԝїR"Ejfj�S �f�+�م[�_�>�X"���*��)��0K����ߡ7��L.�C c(��il��/�Y�GY��@wn�����ᣇ���s���ٗa���^�&?�;F��}��ۻ4�g�ʵ���D��qg�c�r,��K1��OMj��������)��eS��?�3� f䤆֒w�@�X�=��_���{z��G�Th;u�5�W����&��Y���B�ʧO-#-W|�{�i���8r�pA��^�KALU�l��̹���IaZ��+�JyU��xZ�D<U�'�P�FG��0
��8��r\nr1\y]��Ӝ�`[2���+��^�w���B���v�K�SB���UlT���:<>z|t�s�����&���ϟ={����p��v|��Z���7n���/~�~����7�	�3U}L���񢯏p}���j��z��8JX[@`���)+�d���+@G�Ĝ����v�/5d��B:�w�y�ؖ�TZ6�@}��	�8�2۠��^�=/n�(G�!�fR�5�82^�"�"Z���E�#`j�X���C@S%tm"�-�ڈv��KM󵀫��k�f[.G�}.p�~��;�����SKP&oISw�>��ѻ������-��<h��k�ܐY�wi�s��piL�1��G��� Z�j�#8y��m���W���wάCvb�!LL_@��4�c�o<q��w�f#���D�8q�Ǆ��qh���]��W����8��f��K/L�jۈ��83P� ��B�e�f���Ίq�$X�##Ll_8�L�0uFƜ��� f �]bj�Z�\Y�6�k=�6'�#EG\��p#	 Z��P�J(��@����~����4��i�S�P��&�T�FnEhw#q�]M��\.�%&��sY_/1)��@W���V/��n�N�Wk`�F�;��Ώ��o}�[Zt�ݴ����1�|�M��y�P� [k/��߀���&�L�ۆ��&��߰o<�(D�w��Δ���M�/\}��m�	 /[����������e_m��AG'PN�3ǻ�M}����m"�7o��7�10�wb�������w�KD)[�m0�U��:���?����.J��k�y���s_{=�����8jޱ��d���}�) w�0����u��&A�؋%3U���5@Y'S/fj����8P6����n�b�j���N�F�AA\&{��m'�@�&�)(i��n_<��Pk�* Y�ZK�b�Q^���!)4���X6�������P/��&�d"M_:���IA�NR#LK�Z/4ߛ�,�éĒaBjQ�t�,y�iO�.�Iav�o����	�"�p&&+˗
	D��X��Z�8|�,m6���!�U�TBD`��*��+)�QCkS�k�������@bv�(d�*���V��OA��+�R��-n�)G����@6f4�@�	��u��ŕK!�j˳Lp�T"�/U�xlƫĒ��XL$� |K%!����2#�_U4|)���I�7|���TuuR���V��C�6��2��[� N{����$��l��7����9ӏ&�6yH)U���j�����)[S1<&)S�$+L�N�w��9�Z'e�jS&Kae+�W-�*`sn/(~%�!N���<��pMӏ)�ȋ��T�f;vWV�x:��K��iH>�T��i�������=X��B�
G�P�N�V�g���2�Jܾ:�t"̨Ç k)K����`G@�4Jy|�*X��n���S"��0q �\Jy1�Ib&���`{���ݍrjR���YfY�9d��e�pd��Tέ��IYj]<%k��)����@!}L8��dG���<)4��[��2Z�#eiR�t �gD0Y"��M�!#��yj�LR����D�K�w���ϋ��W�g�O'eYBW-˺G�b�];��P,�3C�0 �wŖ���ZAU���*����Rf�bb%HgHȀ�Vli;R|�j�@O\$�B���&82�<�Sh�RuA� ��p��T
�ibZ٩\J\��8r	�BY�k��a6OK�*�*�$�B1Ǯq���� �s���#	��"t��C��	��2��u�,u\rOP��������Q�����g4`j����$��d
m�RCc�!f����ND�t0S�
��avb~�TRJ!Cn�����B�����lSp�J��0���O7�c?���ZUW��Y�����p"3�@s215�F�"�38�H+���sh���F\�k?����8A1S Q��cNq ����`�/n�(ƾ�Nw�Ψ>'Av���zJ���R�۲¥�_�|x�����'�l�x���ΓG��z��>>����W}[#����$!�$�gYX
b0 ��7>[�'V�óJ��.M?Rk�)�`��y(�C<����)�D�E:b"�Y	D�Z^U� �Ԓ��+�5�v#%%vA�Z��S�,in�-�
��)���[KD���,Zx-�5-%��Ԇ9x��NJ��Z!�7r��c6�eY�Yf��tn�5�� s>[R�u�淔�y�ӯ�x����η��F����
,�u	lN1~?]d���^��<�<��C�S��;8�[��>~���w����K{���<~��}��į�xzػa^z�u��>��/Ox�x�{�0����yx\3�l�}���r��΂>��#;۱����mH6��Si����B��W�5<�V��)�Edjd�9(���d���jѯU���y'+�T���"�G��'Ė �=�bu2����{t�a�-ei{�)1eY⬇/�$�a�Qk�)�;�,�f�B�2)K���l�^9���R�w��+�i�@�o;4��bw�����;���o_U ���ߝ�K>Љy��U������v8s_�l0,����� 0
�Ɠ����T��I������Z�ZI�x�w�:R"��>��i��A�N��A3ؠ#����K��Ȗڡ�)��W(�K�p�V����%�BAd]����H	�U9^��������c)V���脛A�,�*�W���<|`!�bA��*��a��U;
���I��F�hq��jl�^�s2)�*���q3�]A ���7z�4L��-��nű�'=��t
ܫ���Zw����/,}χ�>t{��@���mC�Wwo����&�oik^��}��KD�p�Cd�����������7��7��HJ��)�Y�k
FbF�Q5��p��h�n*��3��%^��?���^�u������D��O~bl�=�O�n�NF:�
�?���~�׀�3}�L�b��{۔u!Ě�)�D�����n�8�$��|�jT%�`T8�#�] ���8����Ȳ�qbw�%FC@3��c.��a���F*h�;y��L�X6�a8��̺����n�b˦�Ɍ�D���ZLS�A��9SSR_����Q[
hMk��TI��W�rc;҆i���D�07����i|�R��JL�$�Nݟ���\�pc���������"(�ёW�&0��b����~5�����0G��@�0A�Uf�U %f���9���4�,�'��7�̓�L($+v���q����,�BAR�`iGV�0��_�� S/q%�X#����=e�j-�����K@������YAd�Q b��T�y�'�᫥)h��C��5V[�^<�u��$�������Ɣe�� f��/��!���7Y8�b"i�L����ɷ�9�QX��>ʀ��N�	�6��,�.��bܜbfGp:�|)%MU��#�2�k������8y��t�bL��%˞9u�e��B!q�j�r#��#���*�n��@���Ԣ*x�e8d��i��n8Ub�O�A:��5����
(XjVM�֦�uP��٦{��t��c�ɥ���4ӗ�0A�+$b)f�f���9)���_Nee�L�R��(�Ez�4�l��lI�;Kq:�fKH� �y)g���[�R�|�W� 锪V!���lb�h�ٵ�#K͖1ᘕl� �Cn��aI�l�5������e�L�~64�b3w�"+dhJ,�c��T��-NR�S^_���R�TM!�.vg��@/f)�I ŕ`
j=��r��5�M��\�>�rb�^���+\z��Z�V-�0���I*�^54���J�cx��ߒ�m��C1ZNq��~C�����Q5|4qK�N%�aB2Z� �<�jyQ;�е��S����:���'d�:F5����2�Fsf��М���rn<�@:bs*W�gB��*祐��0��x'�&Xf]�M��%ZC�f	Td��Z�%�
R��x~<���8�(L�Hs6�.=�q��t&�IS����R��5�ζ\�>�j���Ki���YVm)�������La��3O�䪤ƫ5@^�@҅�i��Z
�kBU�N�G�$��<�D([
Lղ.��8L
Ζ6�H>6�3�X/L�]�f�_������F��+�Z��O�4"�H6R��-�Y��*�i�v�a���,�c
��ç@��A:��/�������3L��:e7p��`�~r�w�R���������k_x~o�����c"�����s�篜�t����W/��x��K����ó���]�;���{�9?ڟ��!S6�.���-ۂ��5OK��Gq;E+P[ ��	�^YL)jL
�2� X��'$�x��JJ�G��'�z�)��/n�<r &�����D�
�Vi�I'�XR�;�o%�M�H�j�ƦP�."<ZH4K�U��ʜ��Z򑓲� ;AU<2p���v %3��8B��lU��]�F����%�K���~-�7�d�)EPVj;s�]�e���-�;Ӳ9-������U4v�M�4UG{�?οR�\ʳ��.\�t�셋�\����'�;G��w��=�{��K�;�_��w���~������>�=�Y��>�u��(��1}R�S>)(�y^�H�`p%��"����7ޠ`�v)=��ŝoݨ�֙w-�����R�J�9�&��	3�R��e¾��%b����Sw4{�L����(�)�Qk�.�1o����6#� zS��4�6���^��)����U�c��+��,�8BZ�� �<)�w.L"ޛ�,&���[�Y�zO��g��qdȜ��1��ǧ)֗2���TN@"vyk��ok�T! ��'�����2��D(�������R�/� �/�p�4U����p�z���[vɀ��qW�e:v��2-&Cc���`�ZJ��T��i~����Oƽ��Ka�Z@���C�N;1)/BH�-Ӭ�Բ#��څvf6�`�Ȯ��;�\�.A���5�vD�l����'�Cd���&��v�v] S�K��2���!
y�A��WR#��o��X���2�����ju�K2C����M+pO�������X��J�+��KM��wowtDS����A��շz�o�5wE�yp�������FBklW��0���گ}�k-`T�^,^Pݐ�=X}/h����Hɦ����t ��mc��t ��51�ۣ�Kgb*]�d��_~ٯc���%�x"��+�`�M�������_O����f����@�5��W���Mig��`�����7�7׶�3��l���7���@�ًNkK �v~���=b��)�tK8ݽ}j��Tf�Χ��9Ч���4�{�������!�HD��	Z���-�V"HPK1����#����B���p�1�%`Ry�n-KUp��N��<pL�e�j�	7���)%0�Pc�̍jiB7� Y9)��,��:���(�p��o6K���6H9$Z�Y��!������������Y�F1���>}��pt��f�l����O�U��1%�J��k�����:�2�e��A��ߨpN�Q��7s��iZ�����^Mbɚ!qOA ��V��BYw��f���>W�mΨje� B����Z7��~��SYK��J4U]i�-�0�,����Z����ִ��&2���H�������������Z��֊SWS���L��j׎`H�y�$�ֲ��<Pk�ᴤVP#�	�+`���9���TCZ���x�RM8K)6#UI���;�.�T�ԥB�U~q�o���c�3��CpxK���-������)�#K��V��N���o/eK�l�d)Pc�|��f�*�U�W���Au�]����T�+}� #�["�Y����sw9��\�.�͓`�b����*���t
��A� �E؎*f)#�bU�עS>�ǌ0}�K�����Y|>�F�x۷4C)q�R��]],K��3 ��z�X*��v-�$N��_�˱ �H6q)�r��Ӭ�����XyMŔ���B��ӷ�|)�B���J��/�Lv�R�}��}-�*��TK�,��)޾_��Jd�Wn)@h�b2�TZ[ze�o��y
��
��iZ�\ҫ�Ӭ�e}�U'�-'ML�Ȕ��0A)K�dӔ�D Gn�ډc
X�ư��}�`�U��NlUZj�TC���Q��<["���<K0���N�$rqU|�#h)kIY��8m�Tg8:��nkg#:�cfde;�뾂7L�TA�L��m?�v{o�@�i�Z���q���6������@IL�yښ`�~0	T.�)��d�t*���0�
&� �%�~��Sn�
�
>_����&�c�����k��UiG#q9��k���B��hi%D� .�����Z���ϘR
�b�5���J��F��K��Yњ�oi*�����?�չ5�$��Y    IDAT�͆� hZhdf����������$���;��->����D��V^#�ޏ-�ʵ+W|Z|�
��ãg��.�i<�;�_��p��s�w��zx�ѽã���GO|���KWϟ��o�?x�� !kB��$�5^��~�Z
�"�T�f:CA*�����J��`��
���jm�p*_���ԝ��oT�����k��
��bYR�q�D�|
����"D+�`0K�`1�Fō-�OM�l�b%R���C�j���e��S !�\!o9~�ӱ`��4vK�L�rK�p�2g(��4���C�S,H�m��
����)-U�MM1$����4�%Вo����$djż���^�~�ƫ~�cw���>�z���>�����?��ك��'N���5?~⟎��=��|D�u��O�|��G~쟱��>�����~�]/�o~�~�ī�ǭ��<i"N߼��1���)2�Jx��m��y�B��س���v��;1��k~xKU�QKy��A��<��)��ó��Z���#0�q�����{��>(��������P1�� �@���Qp�]-��˚I�d��v�34����@��d�B���eG K"���;���S0*Se�� �41U5*A�sp�|;���qs ;A�T��������u1�Fΐ�2����b�7m�DԶ�j
e� �yk4�B�1��9�h�0�4�*��!�N�٦|�����g
��*�Y�d)Ќ�/��y�i��c�r"ڡq�B!�.��QR�n�/BZv�˛�ё7~M���z�;O�W�J-Y�v�e�M�K#��h���	dt�`x������<fc�-��<<ec �̴fn;�7�)��p:l�]5gi�����T	v�Ł��k�Ѐ��eU���l�BW�wQȶ�J��ߋG���N�(<���׿���@�.sn�M���#���;����u��ډ�����u���;lw������ğ;M�S(�l/�I�G;��T�%���P�C��A�i޴
�x��x="jD�)���A$�<�{zk�|:�y�����i)ؾ���D�K�	��Qk�̙���P�R	}U����,��n�NGcX��}�1�v;^��?c�A3gwѻ��R�y����8�Z�6�����7A)�.�ֲ�3�	��[֒�`k�@4�U1S�!��64�toHK�ӱS˶d� �7e&%��B��@J��ӡ t��4\5ٚ�=&�8.q:��OHG���8�ь /��^��� [�MaۑW���1�хgq���8���xY˥�z�-S�-���[��Hpi�t�b|fIp�&f�e��ř8�<�� q��E 7@ȿh��[����B";8���#��X&�m�,'	��?�Y22ؠa*�W��p&h~4k�0U�nN�R�Z&���5)d��)� 0)�J�Īg�N�tX�q�`�x�zA�����Q�URγ��ߜ�uVt��.d;����C�e-��0���J��FR��ZV>g�Y���e%���H�E�0�>�_�QH�.�ekd���q�.�<�������:�m_�ZY`�-�׋����v-��h8b8�8�%�@����@˔y��D�vi�ʥ�O'>2��s,iF��V��J����;��ΐ��,p�)�j��fx�Zw �N� 2&�Igj�� +��i@��º[NyqM\-AAcb��֐Z�C � �� ���l��n��V��"���1!�9�x�����(�V��H�n������Ow��9���ƕ�q�]�E���?�4g��W�S��Zf�!�CAP��jY�В�r^S�Z��Ԭ?"���GóA��UM���|c g��3L|>e��:�)w,�4�����C)�* �f;
W���5�SkLH�!l.hM�-ۦĬ�U�+ɣ5p-0W�өq��dy�UH�vѪ*.��.h���d�p��dy���LPP�F�� 0x9>OG�rLHg��,����)T�#��
FK�-�N��8�F�,���8
Vm�iT"�uGP�B;��U`�M&`~�S���*��R\��W� ��h����GZ?���Ώ�~���x{'��t]�B3����I�;}/
�%�TXL_��ʥ���ٲ3@H����������qL8M)^LGL�+ei�v�����@�ĂL����?-:+H^6e��R6��EÁ��ll`U8���RԈ�mpFDP�EMqh��pH��tĲȐ϶ii/F򑈟���K����p,}����#���G�9+���gM@?_��GC�b��1{��}�d$ȵk��x��߮�=��hn�������x�����읹����/x�¥�g�ۻ������w<\���r�^��䎿�O�`����W�����Y����ќ���Z��v�J�A�@Y���rA����ٶ�����.��E�%<�R<rU�Ă�m�xq
��2�|���8 E�� �����͹H��`2���Z W"��-dpW�."|�-���;$M%
ŁIU5%�t�g^�/;x�@NSqC�� X��Bݕt �p%�6��u鸴x���i�~�t��cJg���x�FK���6�8>e��� �\�G�H�{��7�=��ѱ��K/��o����_�op^��L?��dw����C���c>������s{�w>����{���t������gv�������)�	��}<�SS2S�!��2����{ʙA��)a�R��V��ӰgZ�3y����� �����W��!��흦�o)&K���oM �U�<3=<�l��`#���y6�1�am�
��|�;�Ј�F<�B���ǧ`z�	�b�R����V�[*f��$P
��-mR;15��	R�K�jj jJq���C�N�`�ԉ%�T1�2�zn���Lv�,oiz�#gN��KӊUSXG;}W��y4�?�UB�u�1Y��J�K�i� i�ZS����}��e�.�-e�AG��R��NP>��B*G��m�p��(�y���V�L:�T_��ׂI1{������7n��_z��f۝�j����J1g��p_&��N��5�X�mNKd���oG���?�x��%��&Ѕ�}mr����U�G��4�R��ִ}��/%�1��p1���;�@%L/�æ]��j�R5��a��2�?���;�n�JH���� �Y��lrc��l��D���&����7�)�f��f��vAV`��:��}پ��׎lM��'��'ۅ��ˑ��͗��e����3(w�i�T��:LK{����~��_3c�:�wJ�ޮ�Z������/� ��<�v�j�Z�٠�^����ӛ��W���#>����ёzE����]���1�<׎9�ӡ��&�zaj!0s?x*ښ9鐕5���ê�W���]e��������T�tz@R��βl˦>3�~��eu�"N
�hS-�@�$!LL��ȕ�MGAx'f�p:�Rk'f������W��N7�d�$�V���l��
�ɷ�AJ�@��E����x�����e3#�/^\�,�8�٨��9�N�	�e�Y Ϥx��%?��J�����Z >�@�*^�Q���� ������D&���BZ�f��,�L�X���Sb�#U�I*��f�І�x�:�Y���`"�dS(^+NO �۸���U	�Rh)��ؓ�Z���:���KaZ�YU��S��]XK�h3S��Y�����N�IZR`��
,ΒlU:�Af�j~D
�2:
S���䧤��V�ӱe����*$f������/���%\�8������l���CTW��i�N�T�� ��fq%���^���<��lj���"�����!@����F^I��ը�+)jMj;g"��K��r`vn��"� ����}H3}~��m���ZDN�p�Y
���M��ަ*lTxK|�*szo��|�3>/UǙ'})Ԩ |�m��$���)�#�x4��G���o�v���w9�$��@��%�uJRMR���A>$�Xgȉ�;���]D:b�#f�� �k��GD�
�SR\-���'��6?"�
��#�j��2`c��_;/;�� �e�<d
��,�,�'�T>=�.h�&6�B�Q^e��@��
!p�XN�dy�9�)�J$��T���̇��#���~�H'���AK�J�D"4CR#��!3�.���;PU3 �|�)T[�3�%>��/n�t��~��F\�
g��|]jM�F���R���A�R6B1�ڲ�bٙv&Y��G� �w+d}�������q���Ҧ"�e��39��R�|�I��#�U��yL /F���bS�Jb� �,+��cZ�����>)��q��,)�hDZ"ǗR;H�켱�U����@L�
Mq�X#T�[p8&�#� 2q�0��ʳ�b�~8o9�.+��Dj1���
mN��vj�
J� �,>��^G�������e*d����a�5M��?R1#�� ?����(j��`�<���,v�	��i�hi�SC�LRm?����_}�U����益�R�l�C:�x>�����7��B�y+����m���G�����G�˧e~
:<�9��O����\���>����_��<���-��޽���ܻ�ޝ�O?]~[��=>����O;;j�����~;���SK4���<$��[v&�y�L�,Z�ʝ[��w9t��rJ8�J�fkw-0>�ow-��0�
�d�x���g8tB�~�K1�����&����Z����)�l	&NA'�e3�v��^h֥B`�&0e~�.��-�(�o�t
�@aK�D�P���������%`
�,b*UIg�朌Tݫj	�$/`�2�(���̇��z�y2������<��'��\��o�~����ut�����ݻ��у��w��=�=�A��/\~𿮝��������߽����+Ν��Q���=ȳŃ�c�o<Y�:�>i����G�g��`^/�ɚ���B��N�v:R��j�J,# � \ ���^̱xJǤ���G�o�d��*4��iT�`�O�}�|���ϋ��7�Q�|���To�!��Q]�S��P�l�r4Y�{I�Y�h<�)�L�4�(��.�FRB�w|1���+�\�+�%�5�*o6|��{ \�Kߣx�����]�c�8�,r�fK_#Yfi��G��)��l�u�Z6���BȲ��WX_x"N �Gkre'�L��w�ӕd�n��
_#ā�:��Дi�᥋C����nD��
J�q4}C��R��J�Fd��1U��� �ڣ����^vgZ����� R��(#T.&�vp,�]2�h���H�F�GNM;�Q!�u�*���� F�,�i��BG'�U�Q'����U~9����*$�T�hô��i^G�FG�B"�B�$�b�B�8��1]Y1Cp���d�Y���E��[47�.Dd�C��3�+�2f�e/-��J1�J)M��W���n�t���Xd;7��F\\���A֎��~�m7�~�+�~y�)�#�3����B��$��[�\#^�Q������G�yz-�ħ���%�M"hI��� �p^,�j���t!�PA�HS"�����oz���2��?�uZ��Jo-��7�F<YM����4��:ʞ-]2���q��R
�#VB����NS6�%Y�%��_ߖ�
e�T�d�Ȕ�R���K��wed�Z�=��a`4����KSIwE�J:O ä��lU�ƻ�LG4R�`R�*�ԝW�E����Z*i*g���F��+������P�JƏ�Mm�-"���N���Ő�HUhq%�w�tID9�J�/˜!_GA��N@ ��S~��b6@[��r���Z��'u*���|-�a����3 OS��O)f9��� 8>�b)�!��W����B1��!P��A �2�e����}�9��h8!`����-��ejv�嘮��9�e�/<e>|�x��e�Tٙ$�<�z-��J��"��mm��{���J����$hG8�A��&n��6ؿ��I�,�8�ȚY����k<�J��Df8R�e�5��ʥ�� -5�.���
Og�R@�Z������<J�KU0H-�lT�>�`j���y��lcC�'�o�R�@�m!�	5��o��R|YB�6՜�_G
1�#%R
��GĲ!���34e�-�O��{&��o����cT^��ᓝ���qd)��!�3�mw�*>|��ӽ��v�bAH�~�Y�AL���T��*�k��`�G	f�h�*~d���]�<�:J5��@y��j�X�MRI]�q�OUY�,/�:�����F��S�[�;���Ԛ<Z��©;�����&�f��R����a9��ʒ!�4F%G떐���W��]��Pף�F-7F��f突�U�dJ�۔���������<D�e�g�īŁ3�b>���UEǟ�����9!�Z�,Py
���
�A"��x�̀L���YE�/���Ɂ�0N� ��6@�� ���.�,k���&@�Y\S%�X��"�h�ܧx:�S��I�/��D8��Z��� o�~�K9M�1���L�`͖2�f�H���'w/��p|W���&�S�%��m�?�����=53�LVa�.�B�>PS�J5��Hc"�Z�X�X�*cX�JK�Rq�'N
�&��8�,�S!f�2 st�Z�XS�v~K8)4��-+,�	�u�q	(Wh<|�W��k��"�U����4�PU �����h�t3 0
�!���B8��Z�������\Q#��R��ܷn���S㟨%k6�.�5̓s>'��C��۷��{�w���W�?8���݃��/��g�Ν�;����n߹�x�_4�r��Oo�כ����ߺ{x�ᣣ�����'���=w�K_���/��3XCvhnGF�1�4����P8S��#R_,[aj-;�-��3L�LjJ��_6�HG$'�¤�"7y:զ�6-8���?d)|���>jD �t��)���uj�ʺI
d�����,�;*D_H34�F��g�l�릐]q��RcՒEZFSh_6b�R�0[h9>)˂�_m`�d8<���3���f�����o�Ē�B�T�v�%�H�%X,5��y%z�1�>�����={���W_<��}p����{�>:9~tt��r�9|��ѽ�g�|��%�����d�����o����]n7_R�H��On���=�}�j�����z.aJ��7�~�Ƨ�~�d>���p��]��!�C0��e��e����p���=�����c#1��R>�4��.�P6�3�lN��̂���v.�KO�щ6O�|��a�ꪱ`9��6�1��1)G�ޚ��%~����#e��$�udӆ�&̫
������C��ѧ�]?���������
�mFA�Q���Ii�c�Z��hz��р�vn�����VԴ��0��ԚD���ŀ�&Yd�1ܸ��o��E��Ԏ�Y�Z^�[-�L�F�N�R93�Ftd���j�&�����e���u�J�p�6��ק[٨t,/N��MA-�#�!B�N�bݽ��@wc�ǚ�
�ͬ��,k�h���ښk�V���u~d�57D`�I�r��@�����Z�F�Y<]0+YUO߭� �]Ga���!��21d�y�(P
8��.�������[ �Wi��Pǥ�z�&D b6H��	�ݢnr73�����(�G�%<w�M�A���@) ���bTW��1��7o�½�?��O-��^<Cs�+L�n0�ߤL"�D����Y��3�{�=�r��4':8�LhT�ڮ���&�9ز����o�[=�#��}k�pdU�ۛV;��0KF�k��|��\�~�����eo̪���o�)���7�6E_��;G_���=���о��e�r3ˎ��N�T(K?�0/��l%�^��
ق)��1�m�R�ۗ�*�)�3x�Z��OV�,&��`�>�s�I:(`S!g
�p��Oľ��
d]#�N���L ���qz��aR� �
Ѵ�
�2' �#�%+��_mԫQCf~%�>��    IDAT�#515�Ǵ��o�U�X�
Ĝ�1�J��Ch�R`M��R���4_VaH�@���	���3
Ru���)OM6AA;�2a6��v�ɔg-q
:ˤ)�f)����KA��3�,~�T"N�WV3���57���'�S;A:�)����D&�r��M��&K�։ Pގ� [�!D&��nل�~�	�Ғ��2��ڤ����hô-XL���iË�::Ju��B�͗#�,٭Gp pA�m#��<f�!����F�04����wK����e�/K�,&/�aV�r�Tބ��"��,e��g�o��p�~v�񁍄�ăԨ��t�-ٹ�����TM�͌���J"`�L�0��&��b
YR��*�O7I��'�c)�ū�r�g�:Z��G[Zu�����iZc�N���*�Ek��\�P��f
��vT!0f�� U Lv&�L2]�ێ��v�ݲ�fh�:��-yL��|��iG`��U�S�%B kS����*i#۔�ȉ�b�7Xq�������4M�	��GL�BM��KaBBLHwN�#o��*[��	��d8b�>B_ /ū�S+�*-GZ*�Z�����[s)����#)xwB1�2��d'��Z��s;5�h�#0�, ��I�fX���y�.*����0��o�Ժ�ȫ�rz�B�Dm`��挀�x4�.]�ā)ėҗ�Wq��Mym�C~-&۲#5G����Qӡ�f��dfX�~����~�R���������.���'��8#�� ȷ)?�T�CdzA���Gr?��A�`�I��`>���MA���a*���'���TY)1���:Uh,K-̀�.�ױ*x���M�G1~��DVRvR�T��F�a
jZK;����Ax � �π:v�G�х9O�&l�j!���a6�T"��@UL;�i����.�B,�-���n��j���?}�ԋ��OZ�O��T8><�A9q%���ɗn��#��N>�����c�����c������G��^�x�_�:�{���?��e�����������ѡ���'��bڏ?|�����[;:���ݿ�W`��I�F_��/�ǿ�!��Oꔌ��<�I��ۚ�#tV���]�� ��yˬsKa��R�N�W��)��#.aC�ńLV	� 0_I���4 &d���4~�-'�y\剛g��XS��v]����!�E��K[����
��Y�x �y��w�	FyNR���3��U[0�2K����=�����Yaq%��*�R*d�];��ӈ��(X�!�eħ7@Y��8)X&"�ϒ�Qm�� Y4Kq�W��,�Ϩ�>G���ϟ�g�����ݝ���'���ߺ�������c/ꇷ���}x���o:���^�;sv���ݓ���]���/��������Ƕ�\��학=U,]/��҇�@Oro���9pU>�����pԞQ�`>d�´���R�ę���
� n.{^����ڙkgw�ٜUǅ/k�P��qF��>!����_�R�}�QZ�@�1O��q؏l�
�"���J;P�BsW� O�;���PJ�,�x-� Ю�L�y���|2�(7���h$��	�8t��#��ߟ�\?��e_�6�\l:އ��
ۅ��)� �������~�D(��Va���Hiaw�Ep�9"Ԍ�6E�¦� RnA��-�F_9��$��6rgD3�_�rW�����R3@ڳeK �i;=���m�3e^/]�⻯����[z�	 �ij���!nx;�}�	UuJpU��,͏�� ؒZ��}j���MbB�`�Ť�:���ttF*��MەR�kQa1�T������;���b�f�Q�#�L_dۡ��<q`�£%��#P(��#��bVPJ/|���Klם�B�@�<$M'?��k���4?>1��jb�[�O�����{�x���^�������x,ex9#�E}S�w��C�)����]�y�o�|h���Z����U���a�/��t,��ˡ�ظ�p�)/X�کup�v8M��G,-�Ѽ�y-4b&���l/�����v�����6$��$�^tp��C��y��;:j�tV��S2p%���O�W���No���Q�B�F��Ԧ�ޓ��Ĥ)�p�R<P�S2����k�|ٺ4��[�"���T�T�%M|�Jj��ZV(6�*|��p��
X��c�و%����T���5��9!h���{�2�5bR� 5�AR��t���a
��6�ʪ�Qȗ�@J���E�T�cꕎ8KD���hKަL��AP����6)U����d�ሷ��>�(�ZI'q�c�z!�T!����N	M�t��6� Ӓ��v�RJ�|dS4Oʉ��Z��e�J�e��Re�F�Py-�F��xzED.���#��aRÓ�!MR�+��A�B��)�Ӯ�f4������S1+ND����J\\��Je�8�#����%3��"�D��w�T�����H�h�ZA1AKU���]�Җ����:��(�� �=�b�\>eSt��R�|�-?�� �ْ�Xy��F�"n� 1���v8k�S�2�.N��t#���¹� j��HU���G-���h��Xj���l
y�p"pq)83L�� i Lq~�:�c�,Nq�C��v�6	N)^
����y`Y 3dS�t˶������fAL��ٕ�;p8�A��ܶ���k���!��!���,����1�8� ���A�S4�=��l#�ul�ƞ�&�Sv���۱k�ڈL/��t�8{	,��.d[�g\K:���|�eK�2U)�k!�N�����NU1xM�%���/��׉U.;:b
U�`���&Eʲ	�u�[���
��
�Z�_ڬ���p�lM.N����u/=��Ǚǳ�}aw��hK��P�kH������	f��Wkc	�#RM%qD��K_�>�s�]�3�X�}�'�}����̮"ܨ���(��H	,�H�YY��ȼ.�5N��Χ"Cp�'�6�Z��$e1���N�Fj0���x{������F��&<�:��J'�P�d���r%����r��jŪ�6�d�4U�1������.�l�&�+�c���^��ˊM5\��`bA0c@����l��d��
b��4��;to�\_�@��V%nrٮ{�#a�Vo�	ǜ���g�^y^������o`%.���L)�h�c�VYJ��q��7�!J����o>R�n�I��$��]:[Dy�Ԝ��i�T��v��g��M��GSX�R�B�0p��h���ڑ��)}q��ZSm�A�Zj�=�Bq+ǌIĒ����M��v�F������V�����?��}<��;�Xڎ/�k&%Ʊ�?�c(������U>�99z��7w�z^<{�3�_\>��[���|���O�����s�΅��]���x����~i���K_������=��}��/O_>y�o/'��}��ͯ��׍�|ǩ#��9����:��h�.Bwn�Dx4)��+�U	�h���[���9�h��>d�[�a�M��[2��*.�m�B��8M�d�wM2UȐ1��T�����,�*�.:�2B�c̇�c!�]y���W?��l��Q$5q[ R�|��@G�k*��e-�)���j��^��Gk��L��R q�|�����1,H���Fӂ��-���\����QO�g6W�$���}`�)���ǭ�}�yy������./^\��Z���?�'�/����o����?��~�3�|�����#O8��M�G�>Iv�L#�9��o�����}�ok���_�oX ���+�-x�lR�8��h���RL�&ff�wO�����	B��eύv��b���{���s����~���,Sڶ�ۀ~N�S-ic���2S6�%&���V[N�*�Y
*T�Paʕ#{�[23�Gh6� �bj�5��UwY%��RPe�X�2[�F�����?����;V��;\7���mA���I���<�/H�3]���S"�@�$��W�	4m_��dp�����u�U��!�o&�V�^8}���{�D�-�a2A_�RS{A@S��K
m���yj8&��w�����jui~� ���-�8ƶw��u-J�Ƿ/�8�J�a�|��/~��HA���̓F���td�n�DH�Z ϓ�5N�YjLvJ�@�=8���#�jI�r }'������g�"�#� &R�oB��[M���	Ӊ/�)	jAS�6�&讐�_������.|��a��9h!`M�v�^�^�m��bw�K/e�L/gh��<7�����Cx�j dR�8���v��Ϩ�:��Y;����dh�������z��gǲg�~UiW���̾�oL�\/�Q��{����o45b�~�������� KDS:f�\/�M�]�W,��ַ<i􂄦��*ۜ��5��:
�p�cf|ݽ�y*�bI�A����p�)4�ݩ��.F��tL߄L��#G&�ƜLUk�T��(�21�7gPk�R�[�d���NL�-��S�G�h!p�Љf)��$?M|�jۑ%k���)�����|d�6F�6��r�OzkJ�:���0j��p�%^��E������r�<�}�m��O�>�&T[#�Q	7�2��&�d������@�fn�
�.)ۅ����U%5���(&D��%С��Al�@�L�3C���ô�E�X��\�l�Ζ -���S3��,G�o
Ù���Cʲ�Qy��Ejdi� h$}!L�	eq-fx��_
����H��0��lbUdzU>H�2
]n)���])1k/6����ᖈ%�fAqx��*(�/�V�r����b�l��,�tVy���+0�<�����R*�Я~�pH�HS��`
���T:-g����mԺ�j�̲��l�Ng:FAA]���'[U�#��`N�Z��2d�SK9M�u���B������v$P%���H_�	цId�!�5<~%k��V�RqV�e�8�AЌ��`&�bNYA#̄�h��T������Ôj$K�@��[&�3 d�pR�b�Mb)f�ZȲZ���e�9�@4KgUa��+�ϻ�S��T�_�<�T�&�x8D�j�<�~Z@�RE�T#�t��6L���03HI�.����R���F����`�d��G.�pJ�+�J߫R��G��ox�"1�X��d�($2U4����k8C�l���*K;�A*�pH������<v�l�D�*����&+�ב���,��f/�*	ĤG+h��D�	������ԦY�592qU8Z �B<�!𖺸�	S�^"t3�%BA�����5K�p*il�,��U����Hee+�$.�����Jļl�-�B"U	�`��l'P�( �jt�8��5����x��-�-�-���������e޹X���B�Zq� 0Y��+Ƨi�\kK&N�=
XY|1Y�\�^��9&��R�N'e���KJ,;� [6�&�	D K�%d-�4S�d�de���$��� ��uE��˚J��x���1�)Շ D�W>} �dM+�M��w8���p�2r%p��٨�Ɩ5!}N�BBǲ�;A�M�@����##����2�D�X����'�>6�	�vJ��ݿ�2���ח�w����O���:����Q���Пn�;Z><�Znճ����[��y�|�����?�]�x�+����˳���qu�=��ǿ�h6�L�� m�.����R]���7C��`�E�Gt2m���kM��!��!��FВY�4�F��r��B��"�ig `�әZ NKM�
��㻽)C��.��R����0��p1��mh��*e�8���
e�;�8�W^	$�Xaʥ&�1�%��ā�ny�#��S�0��@�ĉ��
��x����gv�-��-�J"��b����&����fTA�� &HMaR�~Y����hK�������n��U��Yv����z������v'�|�KϽ����K�������p�t��3�×��^��_dtz����˥����>L�L�C�������~���^�4$��&�DJa���'?�K{��"�
�K/�2�T�A��gQ}�ܨ��#���$va~��W)�0,����N��	�t(z�h�.9��Z����0Uh>+��f)"��	n ��&(@FJY� ��L��K1;�į��t��(X�x̪x�{�O�.|��A��,�;�9kLT腿v� �li_n,��F<)�] �ڣO�}Uc���<�C��n���{�k��l��w�5�Kj8Ȍ�Z|��� YM�B0-\�Pk���ol������2G@_@�˷�d5|)���&��%( :���FǨ\�,2��lڋ]�"��a2=��5)��	�!�.�>M�2|)>Y}���*���⪔`����%/N��x
�*�g.M���"fTk���V ������Ȥ\L����<�,O�c�C�1"�F6��tĪ�noU��ݜD(S�#r���l�R8�#H��������?>�t�!x ��v�w?��S��yS���:_BMw��q4���x8�M=��F3�Z��h���~�{>�
М����`B?��A�65jZ��4�:�6�0@D�_&y�x"Ui7��c��6�c ��ڵ4���M�0�l�FM8}:������xdc ؂i����A
���e���N�g�b4�Zd�3�M��G�,�i&������ �̬v�Yt*�e�h<N%�� D����k��I63�G��Z#���Ɂ�D���w%|��e���^�<1��Z�0Y]0$Y],�,�QkWY)�^�0�W��S���1�F.�;����bnZ�i��4�Ą0+^K�E&��n䲖�5��%d��iM��F_Vw1/F�:1��~�)�Rb
p4�.uI�Z� R�W��l M+L�>��g�#8;M6��~S�Dd�jk'�i��f��F<�rU�8���5�m/����6��VJА�f��O����<�6^�&�Hu�QXm�qEҷ�'�Ҕ)ĩ�l��B <N#I����@�,�e���CԊS.����2�^�4���&R�!3��"%���=W�+g�W�YG~ρ�;�n{%5B"�R�{���ڕB҉�6�/�x)��.h�vK�O�������v�jt��ɲ:�4X�BF\Pw8����N3��W�BƩK"����0'i/ui�yП�Rhd��aj��Bj��ll}!-#�W�e���K�Z��ÔG�1�c"�G\��D iZ�<��(��M�]ӜeL%��"[�㔪���v���d�;���p<r�C����W�O3qc��J��$��8����\w83mM�-����շa M��� k�-�`֑D�㷂="�
*L�Hj��h�V+fvP��|TI�B�>D,�d����j�)��%N_2��ej�Y-�GR�_��E�Cd[Bb�=��́�`B�,���0e�c��H_�-���>:*���u��.����1qU�Yx��R�N�Zx:]�8J,;���R��(�<�=�qjalH���j��w�8�NM�e�Z�S"N�R(QO��T8-e!s7�͐���V2�jY����@��S��0�|V!O2�"=0{;̛GY��{=�t�RmDJ�,�.�['���w.hmM��4���85M뛗��]V�N B �y[�5��F��h �eMUy�CZ�t���X�%���2>��S��AS��2k�:21B��������t�@:�;Id�jk��q��:���%e� o'���Έ[.󭦣�B)�ä�|����H�bb����-ņ�$؜��N��w�bʪ4�Y���N��?I�ݺj����<��ڋ�;�Űw�=xM�󳻯?x��z�����Ӌ=����gw�����vO^�]�_����ۻ���>�E�����ٟ���v{移�ý��s���w�����������];5��l��T�H�;L�}hp�ZHg� ��'��:xRX�!�j�	\+�rH��� �2A�!<3��� q�\S#սC�rA�0�ZL���Tu�x�;�B�2�:�e��5��E�y"�R��+)n@#    IDAT���&(E�]@,CʆC����)�/e76��Ճq�Qj��iڙ�rjR@cC�Ȃ��j ���I��aZYU��M���u��%�5�^�lU�scJ��Y%FȺ����o݁@���D�F8�}��{}�|q|ww������������E|�y�|}�����p~�����ˣ;���O�}���w�������Ë�7�<�ܧ�^�|0�)����C��|�;}��S;)�}P�S\��������ʜ�c`�1�]x63s/R��ܱ�ħ  y���c�ZY1)�\�c��,����rz�����B�F��?6�WP)*�_��d�mkPJ�%k�><E���Z�0n�
�y8���j?4�4+�P*!Xviv�bD������������o��::/
p��^`d���� ^����b@w����ux)�l��I�e;��!�eM���yx����v�/NЎ4�@
�2�a"Cܾ�}�`_U\�_��nV�\#13�%q�A�Tt���o�b���y��n����5����S�/�ŘhL#s���K�j`����}�ֵ���z�;db4[@� tDd�,�Eq,���W/ϑͣ;�Z��Q�^��~t� �����i��b)�J�Y�x�M�� `�q)q�0�0q3��?���8���l	��ݲ�d�v�@Y%����m����U����Q�Ԑ]�����T5�<��Ͳ&�(p'�-vW��ܜ8���������M��ե��wn$Mݟ��)�I��ׄD�g%tdU!���K��-����O��:����կ~��'�i��u2��� }��
��#�`����<���O��*��a�ygnw�:�`#@%v�����M)
J��mZ4|f=�HiM�!(�ah��N�0Ļ[�)ԅ���Z��Ŭ;��K�{f��dbAcj	2`���ml�hy���ܡ�5�v'�H��%YZ��^kr�Ilk��G��E�F�.@�`"��Hb�3���]PU��� h��Fx�%2MR�1`7�{L	ܩVh��o ^�;���t�6@ˉ�clj�G<&����1Z&�|�c������J5��%���R!e%�.b��h�IP��B��(��Y�W^�^j+7� rA�v1#U[���FP�T��&#�F�UB9٩�Z*aՎ<��j9qʪ���&��yBd�5}�_
yd�NX�Z��8Y�ο�#T)H~�@A�,McȊ��8D���9�
j:UhM�Y�2q��1�e1��y)֨�?��X�<��*���4��Z ��~����p����i��Q�,�T�F��\1}!�º��⇧#%@�D "�2|q����2f�!L/�lLd6j�$��=�羂[2��<Y]�I���B�f9�F���0ӄk_{.�2���`�i�S��i�S�yWXv�V� B@��F0M��"7�B�9�fF���iQ	g
��!q��fH70Mq%RYۙr �P���.�Dv{��q  �ڪ�� s�Ĥ#�i��b��#���$I�B�v� ���2>_�v�j�-#l��Mm[Nat�E��,3UH�� N�RG�h�� ѺW�pӊ��z>�L�G৅ �x|3@�Z� Ϛޒ�Wx�tJ�]q���Z	�ڱQ�,P�(��W���*&1�ֲZ�ʥV�EG��&�*AfK��D��ݫ��c) �1�\&�v|�4�V�Lb�Y�Ԉ@f�3N����8\�
8�b�h6��B�jk�h�d|�@ˎNd�LP/����=_��i�u�_�*��ibJ��;yH�mj�4[�%�귯J���p�t��D�њr�9K k����$��*���8<вT%@:��Χ`i�^�NL�\Jm�]�l�f*�d�OęM�IY�#bo嚪v�� ��}�{��k�L�Ȕ�8`ja)�J��D�,�y���Ҍ/ki�R����{�t� 3K%��MA�eS髣�X��T�K/�v�@�����8ZS0��Ӵ�o��t]�4���N�	�Di<��af�@tOp�o��!��<����&�QM�'�}��<~�W"NP�Ch�ڵ�4y)����dMR#���i-��٧%>�r�z�P���n���ty�}�ͯ����'�g��p����_���?����wwt���׎��_]�=}r}v��sߛ�݃��ݽG��W���w�Ǉ�����+��y����saO�X�c��_�^L�ػ�M.h�b�w�1���86e��3��R	?A|YtYy`�#�+�-�m�Ɣ0[ %�#`䂅�y���ۋ*���X��-��΁���p�����R֦&�dt��Y	P0�XR�t��R��j�0M1�!1S�
�	��<D��[M6��V $�T:)'r��p�6B���V��r���
y�.z#u�Q2�qx��vq�Bg'��&΋e�`[~�4���4Fj���vJA<!���ɾ����Ź���[���.�_�>�]������������ދ���>�����������~s|�o������O�=���Co����<��OL�H�3x��{2~���GK��y133A��exH'`#b�����l�r1�ClOGO�ʐ�t�L_��יn��4��إem���2���s��Ҟ�.!A/�
��Q��� A!��"�63W�`��GP�%)|�8]��8��#�$Ŗv:" ыO_-�#��IV
���L������*L�#�0}���
�-��b/�d�F�t+ 8�x8�@|��*�,�Ub;�}?�!(Q1XG�7JS����1�x5U����Rī�WV�j����:@9�hDSG:�Y���~��_Sfvaw�{�"p��� ��1�ۋoD�5>�.�v�u���cG`#Wk6�<�L��H�9��d��0y�������1�i!V�6���T/A�MGf.�."��^4���%K f�X	/+�R��Ib�6��ֳ��Yx���q� -;|̶	c	�(@T%� _�ͨJ�E�E�)(�,1�
�D��@\}��%��tSyl��������=Ż���C�Q-	B�!��������ps��haI�]��<5�._�y�r2|k�Z"������?�9)�=×�SR��Z�y��~�593����f��j�4�4Rhw�욲My�6 N������e�a�+aj�L�<
ͣ����Ա�
zlB�؝���/
�̀#X6��%|�oBٙ�a��Z��u��Cd!<3�)�͜��
X��j1���"�d��[���-UUL-ߒ�*��pi�>��	Q+�5��LH���֘.Z{D#bB�	����B'者o;&9�r�`GA�2��,7^}-Ii$�
�Ő�J��G���dyH^�%�����2�i�͊V��ֽg�Z�̟B��!�
��B���<�m����"�r�D��ۄӷ pRuQ"�/_*r��#Heb)1~�b;^�#�p���h�e��	��y`ˑZ�_,�S�YaWX����t�D��)"~`RuǱd�BR�hM.�8Ͳ#V[6��$�) ���䷵�)L�Z��ׂ��0��M���20Y|˔��A<
�["�/�T;
pfI'&���H5�eCV�\�����U�&|R)~�4H�û�����h$��R��@K��*P؜_�[�2e%Y䆙�鏔*j8�Z�m��JU[PVL'��T�T���	<�.1yqj���1�^�\w�V�e%����jfCP.�/�#���9��9!GaLKY˪��e�L��&bk=�OS�:BģI��u���,�e#�La��C"�L\!���I�"�d�R�4�5���JG���L��D�b����j/��4�e�$��#7� �I
��$(f�
����)d�9��-��,�m9`]�5B�4?)1�T#�Y�2Y�f�*�"�oє�r���Zf� F�S�'�ab�r�iY(<�8�IRP� �E��[��Z"K!b��A��Σ�J	bJ�aJmqq�§9
J�;��q��nN~�ѥ;�&�<�����ɫ2\��Z�]�^�^-D@�]`�C�n�eS�T�0��Vh�t�Eʖ�@L��nBӎ�r-�YTU<c�+Z~�b�Ef��fk��;�A�H�9�đ#T>����v�_i�A��,�9��H�p����̛b���)��O(�����e%R�<�A�&�V�־Ҍ�����0�4gl���>���u�6�w��	
R������T��v=����/�r�HI1o� UFbۇ���U�R��c��h�N 84:L�Ϩ�|b�ο�/�LN���3����J�`'���[&ئ(�3��<5L�X�$N�F���e�0�z�ݛn�m�Ǐ�.e�>E�D��?�h�㋣c�������������ϟ�����ݽo�������g/���7O�|�;:���b�]��ܻ�w��.�y_p��ݼO�;�;��ܻv�}v}�E}���(��_操����`{�����۔�9���b!�4�xf)eY����4��Z��γFe+W��_��D��Įo٦����
�!�,�I�cA�T�4[o���P�#�R�'ȪJdR��@"�hY��X#K&�ITY&8��|����?��F(�s�͊)��B�x[(Ţ�N˘�R|�i��4lx`"���i_@
�ᘡC��N��t�\� p��K3�$)�vQ���D��t&�_�K-�y}��O����]��x.�wo�t߷��Ó��'���������ѝ�G_��e�_���������{w������%��<x�3�?�d�h#��i&4��9j;���E��W��|��"P(�#��H�vWj4��)�ܴ�#��h$|���d-}ho�f�{n^&.��*={����6M#N��>a��S��-g=��'F.�<�F)�yT�Z��	'S���S�3�(���R��pFjU�!7�Z�<�	0y;rD0}@���vǣ����4_,��� �l�����mJ�B�)�ح�,���t <�v5��0B)j���7���R8�K�몗��ܙ��BT1#� M��Ra�ʍ�;[���"G������^fs>�ߝFj���K����(7C�_\@�C�F�x�
�b���B����}!kA����	�Ҩ� �*R��8�u��q��p�w�HI94� ���yK>�^��Y9��0Lq�$�KeZ�ě_���za:�CHYVkdYA�
���ۗ���X�_�U�8gfWA��.��[Rۊ8��S�rW�Q#(��WH�%~q����f3'�R���o��n*L��W�����>l�6E�f} V���)��Fu������Ȼ��Bd�����2���i�	�&�0pH[h���9h4s��7�n*��Jx�My;��ڵ9���KS��fO��H���u��6�yLk��d���H<�TKcS#b��{[E��Z�t��d�جa�%�NR
m�S��#�4j�նl�tx�v*F��;F"]���mwzY�)%�)k|j��iD�u�U��-�����4�LJP	���&e�`� �+�����'X�qd�@I}G_P\k>~�u���Z��)@g���4�^����^� A;�F�Ĭ��!���Ji!��_O��� eU<��Po�j~cĔ��U!�k�_�����&�u&S��tI�oxR���+�d�p������ڶ�s�[t��9� ����*˵�B�}���t�O�X��eA-F�,��&�9��oSt�<�
�f�u��$S���T�ȆC�%���q �\\�2�I��Z7'_*P�vN��jGm�q�NL;W���d@H��bR�T|�� ĉ/َx�8-��R��Q�G�j< S_��l��uU�4q�DU�Y�lV�e�u�#�$��O���Փ���S^j�K<�ʑ�bB�p�[�z�'B��Gk!@0Ico�� �E�t]�MMV �����52mAHU���*OV�to�8b��xw�8�n��h`q�ƫE����Ȫ�	mz�-�O��j	�'N3><��\��|noَ��%�"V����5�ꊈq�PP�6�J4��4�J�2�3�Dr]fS�l~%<��\�0i"L%�A
"�&;{�w8t�tү/~��X@�I,�0�8_�%�/�B\�@k�,58f;�#�+�i���]��rW���%���5M
��ե��&�o#�3� aj�d'մ�jT!N"�V\gY�nF�RNG �/H߲�Ѐu/;w�����d�S_�`�MI�$(ے'iԥr�闏Yk�D��l�)k�f�G9^lI�����X�bU��Ł`��>����d{�[��Z(4Rx&LS �Y�h@K6K�8�[�M#�J��u��=��o�
��{s�'�\/A���<q�R�jYq���?��?x�m,5��ˊ�$�x���������$��E�I!0q�e#��hd��$qq�Ehu�)�/�)6)�&�7g������h{�Ds]���!r�������T�Z4���aMeٜ�L.005o��<�``�5R�褐�I1%���� �� ���F����*�8K- �b
�# �|��s�j
SF��ka�Iā�dD0Xׅ���u�j�|Bۅ�u��H�����r7��'N������ɟ>>{yy��7����_=>�w�������ы{��r��gO^`��-Wa��w�7A/���������W>����������ٹ���8�8��[��_�[0�MM�i�������G
bk��d��WSD�k�u�� ���5J.�Lym���9�P��L�,g�����jyLF����4Zj�I�,ڀF��t"��VRӪ�bm�r����,\ ��r[k?�T}S�Uh<�l�Fzc3���%3c�+�R�4*�0�âPUÛ<�
��`Y|� �rA4~p3�Ɨ�P�dn��@Xw~.\-� �AA�U%H�BL�K�U������]
gW���|���w������ׇ���{>��ϧF�-�w��W�{׻����ݯ������_�V=z���_�$�s��M�^,|�4FS5F3�9d[6�g!���T��L\���{^�,�Ԁ��Y�#)E!)&�x@�)���}� ={ �R�|�/ ک���/��R�'79T��jD�Q���@��2&�[���TS-\o%�6#e�Ca� �EG�����za#�A�,�]�N��d�eM���y�6f������/�����U�ՁP@��גo����/N�F�����Y,�/P�� ESw��(�)Yff���֝g
]�ΐ�q��ha�~�H�r͗��p��`�nR�������q3Ha�����55��s,E�f�BKF�0��`�c��MV-P�����Z
(�e3d�h�3�C��Y�U N�g�+W�,0�T��ɚ'�M���rG��D�l�$ ��!b�Ec�wH�q0��yL���U��B48Y~ۈ�*����8@�����g�x���
�0#��)�]�zYvhj�f3'�@���tx%Rp�gI��a�O��<�g�Rh��1q�)K]��=��n	j�X�7���{�&A���g�d�_%�f����G�a(���+��s&�*8�8߷P�2��_��X=S z\h�{;�s��\�IZjG�<��R�י���dQǄJͦ�B��
���N�){��VJ;L�[w"���.�ꠘ��8.�hz94e[��L� �zYҡP�E�m����	QK�RIם��ł&���U+�&�Ly
�[�򌾃���x�fF�X�9�z�`]�)d������	c6?��<���p�����܁�]��;7���<��j�-�0���L���wD
�mS�73qǲ-/����1z�l����q��Eݕ46Y]���PS�^��W#��/��*�4;@-�b��83��nie��?�N. ��0�i�-�UY�`NA�*��6X/^k�Y
j�V�B���WER,�B��A��5�� ̈́Ѵ@���Q-�I e-���َWmY>�Z���͢1H}c��Y`H#YphSmA�9v�
�t 5*ƜiRhl�F,�@A��M���T>2���,�*;�� 4���\�7w�S�F
�/���j�����ٲ����մ��p�1y ��V,E02P�2�C&�%)&.(�	�r�[1�.@OM�C �by��4�h9�|A#%� R����-�R��.�DW� �,��L��	���X    IDAT�],�i�Ǘ�o)�^��˓j�oZ�2��Y+5��M�|��Bx�w�����"U�oSt2�?���ֈx|j�w/R1�����u)�k����T�
g�r��M�P��XvnR~Y�d�'o����F��s�_V)�2oI�����+�C.����i`NU
��d3`+:�>M��+�!�T�|��l�T�J��T��J�i�f l̆���@Ҭ�X/AH[�&����S���&����+oH���� rR[Z�))�;ZK:�~qݥY���o�����v*���Gk)�nM	#O6�ށ�m-M������@:.ԛcW� -�����#8�8��T�l�Mʒ/�yqA��,��e&N��!�I��56��]hqG�B��4�l }��D(�7�*K1S;Wd�_�@0��t�)(a]M�nZ��h�N`Y����`you�-��� މx�Tw��9�l���OMI?�xx��FX�Z�ȼS�)֫�K��5��Q���L%���Z��̀�2Y%ZX�h�)ｿ�S���y�Z��&n�0S�����e���DF���.ݥ��9=KM)�P�-YUJ�)�*) qo*ql_,��u��%X&[�d����[�]n'8��-���Sw��ZV�k���R�
�)k$��bR�8&����I�.�N��f.�����A�������g�-�k0�t�>���ݓ��ћ�|���7�8<�;�|�`�L���>?}����ԟ�uR��c��K.��˃�'�����B��~��`������ť�F{����>�{��?��T���G}��h�m� ��^_=	�i8"x��U9
K��Ѫ��3�ˁ	�O� x��c��(H_Ё��S"h�FB " ��$���e���PPXm�<A(PN�W���R�L[#�vrK3��§jh�IY�o��i�ƴ4�zџ��#�ˆ�	�6s%����1��۾��y˭/��%a�����6�8�n�D� ���jp�u�#��!W�}LX6D�U����BR.�Xa�b�_\y����O�ϐ�w������ޝ�������������ë���3_Zվ���O��˯=|�_��ڳMO2��<�x�Y�d^�m�iK����OOYR�
I1�:O_�OA`w#��*��$�ԢA��	�P�v8Z[bR�d�������/��˿��O~���2S�\zy�U��X�Dd�pR,�ɓ��u���^~Ę
��L�,��l^�i�1+�+�-�Ty��W�� ��<S���T�Ll<L�M%`q � ?p��~�}w���&���W�����-��3K�h�z�1q�x"p���l�p�^�q��k_K��bݲ.��/��y���~��҉u���M�C�tPDT��@���#�# ڎ�3�S���m���׋�\P�Wh)Ы��]��nYj4k��i�`��j�����v��) �G�jb��	"�mJ�dLyM�<4��FGa�d� J�,�ʛ(`d-��o��E�+���p,i&�F\<��YVA,��(OIㅠ���P/K%�6�]S�*[�3��P�Ӑ�"e���B>s}�h����0���O�l�i�.��]�O8��b�)o;�MG�b��gO�~��n'�N#
����h��R��/}%8ߘ�Ώ ��a 2�F��E@<)LSy�p��Z�o[=���	U^��PN�N�\)�]��&
��{���E�Zh6n�h�&1��������7�ʥ�2�mZ)�H�)Qv	������h��P�n�8��hR�-�L�v$h_J�ǒ%"��'%���Ҩ��C�V
��@ީ*��)3��6�DT"h��#��T%KV�)g	J��g�Ԗ���$$�Y��ZB�T�J�21]��"�Uw�N�����\kAF!��Bpڝ��^p��WBYj&YL�ZX�)WبxRL�%5A
�Ͷ�V5)���R G�__��b���/f(UV
9��)f����q� 3��B���p�R�
�Y�	��GkN1�
-��R�����L�8��h]A�ł��p�˶Y���L�E�2�-e��r��*��n�8I�S5��4@��.������8)K ��Pr;	Tu_���D�ک�D�]�(�Ū�\}��Q��J�(}`HA����j]�GбӐ�f��#����Z�$����ቈ��T���[��7��I��Á̴=j��G��o`R�W��m��Y�#8A%���1mJ�*�$I�Y���5�RJ�pӏd�9
��<Kj|�3�':���20�0�̲B"�JX��$��J�T�+d-�vB�%�6L`���<��Ո�G������/��/�f9'	!"��ZF�O�đ����'�TRU�*<�J�-/X�m�Ȕv����O�^hR�Eb Ͳv�����G�e�Lm�$5S5F�)CFAa&�Z����aZ�OV���v�)$�ij�(�$)�#M�V
R	p*���;�r^U"b8>K�v!|"&����`s"XfucV��y�+��B`ݑ�M e*������1�]�k���0V��xJ,{D���x�jqKSU�J��67�HY:@YU
ŉLg|����ƶ�R�w,Ρ.LqK^I�@A`��t�b��l鈛M0q|���Ҩ]�hp`jm�F��@7d�
�uw	�Z�zMa��עW�SLK4
��3�4�ЩB�rl���
{,xo����+�6}���*[΄��b�8���4�w�J�R�)֎i]�\��)Hg���50��l�p�1)KR�LIUS���ó�XI���Rw}�,M^a�%.�g�|bӜ�h▉W.����	���H�$.hIVVI� v�ޥ������f���CH/)��ܘ�C(ƙQ��e�<�l�y�4�L� "��C�iy1�vQ�&&ܲ���L�#8��DF�iU����K��>hZ?�:�{x��[�;�>�{��������ӗ/�|����ՋO�����Ş�x����Q�������hyu����^���L��n�<<����垏}�2�1�wP�bx��m�	�����G�xi��C:�b���p S��F�QC�NS�l%&L�rKA��9W��us����$ś��3>5��ldK��5�R�qzE�^���FDЈ'�g˃$%. BS	_	|Rh �c���af��Ʊd��)A'[Y�di���7dK��*��X��Q��+�D\v
�b���zz�I�.�ν׳V퀲��̒)���
��a�����<�-}��'W{G~�z9����W{�6�{yӸ�[~��?V�]���g�/�g��ݿ��<��\���l��g��x٩�K�k�UL���	���{�j�R�u�:��p*�Y�^���h�#T���_��ê嫢 ���TeH�k<��������_�������5^��#���P޲A�ϋ
NT�=̓ݦ1b`�bv�y:5�Ak �v3ᨒ%5|1ڴô�>��b�)��A��T�-���[�U�b�'�s��C�:2ߨ�"P@����H!3\�B
���·`q�"b�
ՊV�%��x]�J\&��Kc`)����J���~�^�aB��Z:�OJ-xߋ�u+
&D�_���O��O�����ت#e9M���<<���J��xt%�c�>�0dټ@GR�jx�%Ӆo;6��_�AKVP��B e�������Ѩ�!Rdᤀ�%o)N\# e�ChK����&π8��ȵ�0�D*k�dI�G?ِ�RLL���&'ŋ�h��ʵ�x6k�� ȞC\/7�eg�+WU�^����,Yt�vsh�.%�kAD�`�rC.���_u������y�/�?~�����'t܊nݪ��d%�^ >���(�s�rU�j�T��Xlx����u 6�4���'YǂhG���nƨQUN�i�5Yf6:[���V�F=���T�t*'7��R��<jc��r�x3���?tz��o���O�,��H��Y�G�@V,��|�4��0�c�T��+���\�C�;R-:"
�1�, ~M��	S�;�k�J6s����D�c�m��̣���25`��	y{W�-)�
�BY>���
�֬Z%�)�C�����<4-����#�� ��Sbxj�/���S恌�*K̔k�aE�9�_
M���zu��*,��C�����n!�1y&K?O?r���lm�
۵ !?�D�pY�r%��;�! c��)�t�JũP�����)GPX6���Cd�»���{u�M2
R���\�����"����"d0A��N_֮y�^������j��.�A���dӬd���<>�	�DaM%@�C&�L��ɶ��H�F������Ya�b��'�	�eH����3dc��,Z�=#;�f�	Qۖ�b&�
2L��&Y`|A&۴��J�.)��M����@>}�R��eF4��lw`�e�R�Н)�xh�-%H)��31$)`��7�
��q���GU�nghԑMp�j�7^K��8�'B�<$�8}� �⏔�<M9�'^|��6�-��C�OM0M��p}qϢ��v2'�nז��_�.M^SR�KJwK&��6��Z^*PW�QT�/B�E�"�3y�8&M��Ӥ�E�)Dk~޾J�̕�z�4���j�	��Ȑ��w�hā�uXN���p�s���p>e�~�j08}���[.}j��L��dYj�7���O����[N����ǪJ�u��\ax��-��)���<��-���7@�0��D�h)UGY�R�YH4� gV[w� 2H������Y)�j�Qh�f�KP��D�#�
�z����f��5pD��oE*i�t�Lm��z�l��7^)"
�uq4�Z��F'f)M�L-</���c�R�O�`eUY��30��ǅl6��Q�S�i�3�޲d'E������V�{�z5˺���!�ҋ�-ua�1ͦ�^��S�S��C#)��D�1)T�0�a��T�������*�";=�-�c�I�!��f�p�
B�/ ��Yf�n	'N�I���>c�4�7�8�yU�[v{�"��������;[��wyKRD|���Xac�k�/�<�o����^Ժg|������^��6>�F��8ıe�]CJ ��Y�Hl`���>�5��0�a��֧U��k�_�������;{���w���O�ӊ���/.^\���w��w�|�yx�箯9�K{�W>����>�)���3xw�?Z�;��߻��[�7�}�`o���k�;k�3g�����6�@,�d���@K'���)��{1/��� G�N4���v�bB���mY�a�#+`R�S���T״�Rj-��R�M��%�"ˊHU|�T�Lsc�Iu,�0:���n�������iC2P�Z�?�B�9�▔զ�����V!��|
�-�A��N3Pܲ3Q��e��TpLx���-Rw�@
�8$\��edL�i:d� F�qO�w�S�PS��s�+�a��r�����;_�g2w�������=�����ӳ��W��;���;�xr~�{����ly�����^{��׿���-�C�w�}�ӎo�|��K+�l{^]�/�]l��{^�spc0�`}��	r��)�"v�p������I�s�d�,��vNI�Q�?���
�U�s����?~�����Ʊ��,O��RQ]Ŭ-	���2lY���@0�:�2Y�_������B1�/�Ph�:A#�D��322��/0Z�S`5M�̲@|d �i����5�����d
)ۣ��-�j�_���~V��Nx}��t�<N/̦EKY�� RZ�/K%��2!��f�j�]`���ʒ�yv�� �JDL��u�����_�K��;��BiZ*;L �%��H|���H�>�R�UYv3(�/LHC6v��Klw�k!P%��/�"4O�B0L?��th���dm35Y��`Zq� )�.�Ll6�|U������B��B�Z)L��-�l�j04�.p��B�#(gmJ*eH%|`�<Mx��
�U�N�H٬�(kIA��jr��:g �bx}���e&�-F�_\����/��T������..)%nBH�,7j#y����3��r1��i�!���A�p33Y2)4eK��O���u��OȊSs�0f6�I�R��ľ���3Yۡc�BS�z"Ҕ�aͦ$2�6��ܼ���sК�@��(�`�V ��2�F�<$��u���OP*/+��h�ó&LV
~��Z)�d��DL����J �t8� ���n[��[�)��M<��Z��DB��Q- 
�_9�9d"&��M��I,k�<��NI��_�y��!뾵/70���W��O�e-tw���iK�|�N�1�P�zgNq��Y�c6���e�b%3�F@�.@؂U5����o�&o
��$eK�^�E���}H��6�53K�m�V����@�d������I�>��
5�Y�9��
[*��d����� 1-��7|�4���T�[����2O�)�.��ã���ff�*���v;��B�Ly^ ������v,1�#Ȧ��ް$�x����J/�U	�@V@��	J5 �l!bH�ԯ�L�ZӢ��9��`@V6�:&�X��mh��W�.�u��m�JB0���!���<f�Z�EkB�fD��v	$�ĕO��S���*Y�_ݺu�;�V���S(� (�`���u$�T��U�#(�# �R��@���+��'����g�<r~�bY�8�p��0�U@n^�k�8<�.UK$� �R����YZ�jh�,����FA0S�6��#��#;�3�7ټgF��[l%r�1A��X���A��)?�������ǲ%E��f��K��9�K��N�p�ާ�z�����&�I��g�:*Ѵ����u)ۣ��7�R�^�� ��f�X�l;���.��]k{QRaRC��_���2�
�%.�  �u2q����SX�f�fV��D�/��,:���2)/+h)�4v�ļ[��{X-��SH<"�/e{ߩ��cx��*)Z�����	'R�aB�6sjs;U�܍D�RU��'�,6��bws���LyÔ*.�Nʆ��@VI���C�Q%P"@.�2� ��wK�Rk���^\	��O����/����h���6�ﴦ&��J�8D�Q��� rg�`��-S�L�G�5�*p�܋��6��M�Z�pZ(	�f�V�Y����@R��7y����U�����
��}K��hd�
IUi K�#�����D�o�} �M ��4��H�!mG`< q��}�.�|ЀR�nH�)�Em
�c`�v���傎N��!��%�#Y��Y4�eë!����
+O<�dK����eŌ�T�
oH^
'��i]��`������v��e���%N���A��t���k������(dy��T���E���H�C��Ř����.n�̀0�8�4Ř��8�A6�.P��N��H94��BJ��j�-��v�;���|�b�3���gGǧ~��Ǔ�==?��}��'ۣ����G��	p�����F���p{zr��\�\x7�g�O�^�nvW7W_�]�6G'go~��7~�����3�������p�B�N	����bʲ4e�����I�2�	�~�:����ԺRRԀ����[R0�u�IA�q*���q���ZF�'����(_[�}ARyL�Q�Œ�]P�7Y������G�,�+�h��l)��)���6%0�N�_�wORe	�j�;��Y�_��^�.B��q��/;�ʒ�8S� �M�ע��o�y%�T;�O�#Q����8gL��@֫5����v^@�N���_{���3�fwq���Ͽ�}��o�|�\�Tu���T{�;��a��s���N�7�QBo�u�s����Fs������k�r�5d)S1����[O_���i �	��
-�bUzl��F�o��-�2K
u�mD��.{�Qև_�g�#cx^��5��￯�w�k���Ş�p�}a��<B����X�z(�0-���l=�j�0�.ZP��b�`�	o�p`�I'� �W����۵G�@bZ��z%۹7?�ʇ(舼*�����v�����	�t�n,��Sp���U    IDAT���vO_s�4����˞Ft,������=�7���x�/k�^p��^|Y�@�`pL�5�o�[��-���0�w�恋)��W>CR� #=y��i�A#�Z�#>��+�Ќ�������( .e��l�!A�AJ`��� B�7� ��#�u������1y��� �Ts���#�O�~!<����R:��I�%�NW�R�&@PXS*�R9r)c�!�vZ0�}�h)ÉTeG�r~9���xK:�5�v�^����J���T�-����o0#��<��s8�t�m���z �74��TE`��j)�,�$N�n��l�8AO�~�٣��{�8�l֭Շ��F��v:�mNjL�� �|�%�l���j�"؎���
y�t�cb
R���v,+D0)����d�:g(ei)���J�� ��'?�ɿ�����Gڡ)W(�Ȗ��͉@�w,p���	����ᥖ��J��շ��i�n77�����Jq�[�4Y���w{��W��upy��i�ѧc�D���KI�Jp�L�0�H�5��?���z��������+�Э+&�i�ĩ�k��6�R�g)�HM�x�zy��A���(֋,����!������륖`�Gx�`�0lj��~4
yAS�8��#�@>�����k�6_	|���:yK�lM.�R���ج�����ݦ�ݩ���4����T".�JU^_�#j �����Վ>��D���[��i�d�*r�u�L'P<8$2�Ͳ@SY{�0�Nd��ɲ�N@9p��r����/P�0)A�����"�B�餐��ٟ!M�I`��,��.��wB˙0A��b��N@	�g�VM� �4[kU��bD�6ӦlY�ߥI��|�� �k]Uj�e�N�'�3˲�>YKU�d�y�T������W\.PB'��h���9�Df�4�B���Y��إ,k]���ע�IY������(�t��J?���h���2��L\�T`x N&��@�NRܮUA<��j�uJb�4Uɪ����)���
za�'��j������{SG�)'2S)ti,MX�՚G�đT�k��m�:�j{퐭*��pR��զܐvJ��	�; k* B�|�N�ٺ g�L�(X�B��,ffHa�S6� ��#vJ <$|�*���hƩ*B����q�F���έ�e���uS�����4e�y3���J�k�))���WE���C�IZؾ,2�&�3��i$"ۥA�c���04��"�8�,�R ��@1�'5�Q���S�*��d�����C,�SU���a�G�&&�h5Jh��l�i��P����B�Ҍ���jԃ�¾,ZC�=�V��JL�Z��.P��˛X�D�$i���\���:Ψ��{\(����U�ND����|��{s����8zsL�U�l��b��l 3@̿��s��7���z����Z��e�����|U}���d� �C���'.�iZ��>%q4��)�_z��OU4-͌ P��/Ē%b)�� 0�x�)�_M���vp'�Ku�J"�
FA֒��;�~r����0�����W����H�l�<�з�=R0'��GvRZ��W.�~c�mG8�R�&E�T�}^�{#�wtn~\�7�@�>aZ~������ٳG����g���?~��g_��?������}�������\>�^ȁ��?>y�9<�mN�v�/.�/�7��O�|L��������nO��h�3ңG���G�����η�lN3g���`v��-;�b)�l4q����"fp1�0d���;7�3���U���r�~s��ѺQ-�y
M��1y�bLV��^R�Bcp�ě�v��<rjh�Ì����l�fV޽��J�E�����XP�!��#+Im�4!Rl�LU`�zu�S2�jy��C���$b
�++�cZ��`�z�D	���R��bN-�M��;�*pW"�@�X�.)hQ<�5?5�����Yv�ܻ����'k����٩O�������������/�/Ͻ�w}s�ݜ�nO�v��������|���˧'�wo}Co�-����=��=zx��~��~T������if�ٚ�������c��_��_���-�^�������������]�S�v<B�pdx~.�%�{�B�f��ҫ*���r�goi�צ|Ц��H�xTi�'0tB8��R�bF2��T�b�����́��[ҟ��͒�(��Tb�{E�Q����G��C���.����Mn)����M�WV���~F�0��d}�J�|�ᇿ����+��=�����O#,kGք�k�W�� Aй����k�^>����C�N���Ҩ�ȖŪ4E�d|������H������?��?��?��_��_���{nU�B`b�<��K�O4�ӟ�fWD��"�Yvz���DI�:4Y���n�����o��G#"@��z����  K�$����ܷ�?;"Hy���3 M�ݷRm_��� X#|Yd�C(�N)ǯvʕD��ӑB6���Ny
�˔�	�u��֖��B� �BX/q��f�\S �������i�L�ĥ�1�2~�2�y0р����*�GM650�4�����(�Gw)#覒����1B
R�}��Hy�D�&�q�����~�mw���45��]�0�$�&���!~.��E��)�I��M���1��M�bK�1xs
<�x�Pw�F���D!Y&���ю:c�"ЮC�{8�}�J�ԢI�B����H�H<��k��h���CK\�%o�ld�5��7�����`o��8}��)�$6�Ɉ�C��ඥ���OD�4�2�E���Z�@M��Cx�d��'�G E���L%�Y����T�֊1!b
���~iҡ�R@�������M�Ē�.|jR�+�.�g�Dx/I��F�Yadqa�Ⴙ�dc�!�I"h���)�(�EVHM�f�4�Dc�����IxR��d�ᥔ�D�uDp�b�b
XRķ�A|�R��췥]��r�!dyʪ����EN\����-;�� *iY�e%v�H�|�Z��&�0��������jd	����Z�SU����V��J��#fI��!���ŝ��Ѵ@k΂���˹�65{����o�D���Wܒ�o��dSEY˂�j�X�MI5�0�4Ͼ �j�2d��Q�e�VP�(>�)����Zww{��dR��Uզ��BX{O9�Y
y�����M,;U� �M���3����� НP	o!}qK�ҙ��瞥���s�x�(�S��l�q
0[�
�	�@l���@%<�4i�pA�#6a��R�4j��1��2~��q�d�Ĭ�ԲF�Y��������R�ڢ�j��, �!M�l�8�������@��T�6U��C�9��u'� 
�V��!׆w_k�H�SB�e��qҏ���\a��_K��Pv�1�9�)I�9�A_V�	�
���A!)��:
��ȣ at�A���0��l"K�
�E9}H:�ݲFx�)�	/ND���ǚB�	l)��6�e
m�^�8ʣ%U��"3��Q@�/`U��i�
!��%�O��7�J�3��-�-5m9�p"@�ډyYL���qJ�I,J�h�q�j4�((o�t���۔��(���us��4��ZU�ـ����I��v���
��͌ߐ�B@yFU8}K5CS�w��05R<`�@3*0r<Z��t�wqg:�����N&)����u��<��C�h������78���T4�dYc[�V��Qn���ɋ�F�]KU�C��1ꂠĲaL�F�7hf|�^�-�:�F�HQ.�&��W�0-yL�@U�� 8R�DֱT2�#+a�kQ\���KÇ4y���&��@�	��8�
(�Y�uQ�PS�"K�Y�tV��۵)�ݷ���7� �K9}H�����F
(GӋ�H1�bV
-��#M��
)�E˒Y"7�l��w�=[9e8f�K֛Bޓ�6�w���]KoJ���[�������{����G_;~|�ڋ/�}��o�����Dp|��=^>�{��ۓ�ƷׇWϟ}���ϝ����h�\�j��W�����7�>�p��!��@ӎd�8f_b�By�߽d8�p��G��5G�_I'O')���#(�ԋ�P��V�"�X/���5R�b`���r4' ��G���i�ыx���)4L�zu&ݻ���&Hy�
�,��l�t�oTX���B|�L��oB4���J�'�p|x1<
*)��?
�='tD�����j�f�iT�0��	 �NK��#7v}�-�{��,qxge�lл��o�g�-{�2!���k�������b�|d�C��s�~����vwq��������`�9�z��p�����ׯ}����ï�����e{������zf�7�����/_<�ϱ�ʯ���x��v�٨fxS9[�	8yY�7~�������{?yj�R�4<'�O-���	�	:=xL��K��8�a�𥪂P�m/�*	���ӗ���<� ,����@�Ԯ<*��±몙6yY�K�)��l�F��c64)NY�Z��d� ���2&�aJ�7��XI�����S�&. �iϖ��f��*�������(��D�������^����ݦ���	|y�/�ќ3���]O�@�����6���4���1�ٌv� 4'���/Z���y^]�^YJa��ϧ��"ԗ�W�_��W�W�W�}�frL��)�=w6A������?��ϕؚ1��� ���Ju�Ζ66�w\8�:^)kK�c�#��_
NL߷�z�E1O��5?�,NW9d3�4�d3����@>]TũP�Z[�p3W+�DL�ֶi�yU=��Y���k
�$ł8����!�h�e���'�
M"^��'_I`�.=�*^(\[-N�	x�h�K�%1��0@>��G��Bw2q�6�+��p`���u �n")x�ɺ�C\qO�b�D�-����<�B(/��e�F"b6]x�f�4��o��|Ddq���c͒�z�-?���G��9-��;|�i�y,e��X�C��5�!\�8ݙ��S�˩��0!f��y3���#Y�.М�e'`NqG�od�~J �%�s�K�,��y|�� 7mc���i�Dx�'�@)c�C&��Зew��!��l��в�4B���de��ؐ�i!�t�.%2<���Vi�v꫖�T��*t	��H	lj9��f�4��ۛ�b�M���;�N����U��w���z��N�@��� X��w���v*f��bY~?0�e��j�أ8~�k�ݓϾ�SVI��X,+�L�����4<��6��*)X�$�AN�'��cN��e_aj|A[H\��I)�T>��Rͩ�U0ה��@�h
1�	�ԔR��ï��<<)LK�Fd����{���T�N~f��%Ô���1�@d�axK��ƴ4*r�8���墻vA(X��w'������V��d�Wk�� ��'����e��.:���!�+���^p�$��\���0ۅ�)��q <p�@�.t����������NIU�ڣF��m�#�%���%Ȁ<f���S�V��}eH��+g)K5e`�de����FԺ�J��(�c�Y1/n �hg&��$��!�t��/r���i�2�&fS�?���zr�V�fㄔ�)?4���g8Cn/÷G�e�1[Ȝ��*6������h	'���RmR�Jp�º�k�����J�j�#��v$.H��šä21�+�fÇ���S�<Y��B��J��c�7'�d��%�t�\�&�v[�2>߽��l��,�R� �CVۜ5�� 2�h���D`��:�6� 2�t&_Jv*�ҜB�z���TQPX���Z���rx�X�AGK|Y6x��y)�@A��e��Dn�t�v�$��t���K��T#�̗�}g�N}-�
��R���q �YtW����0A�@	A��F̥�:�,����u4SÉ�җ�-��QϋY���!s��XmR���_<��f!�4��i��_(��+�em�p�l�ၚ�R���F۷�A����C���������]�<}�`��:�D��Z�8+x�W� ��J��7̦c߭�Z'@��癒��Q
�2}�,}`��mJ�yǝ��
�F_ms&�ץ�����xq��/�V�`�h��F
�41�C# �W� M`rL[��v%�[�gގ�j6ྲ����:6 _�����4X�4~:Y)��%�:Z�  �U��2��f���[W�֨����}cSU�J��y���?������˫�~s��Ƀ��ÿ|��.??�\~����ۜ����~�3<��e	��L��������ţ�>��Q���֛��㓛�Û��ó׾��o-_Q�k�e�E �-�{8N�N�I�lw�����d�d)@��3A}C(�j���e��� $���/N��.�H*Y��{�ij�~��)G�������W%h�J����Y��΁H!L�,p,���Eh�{�T�)�f3Ԛg�*/g�	����J�jKŴ�B�Js�� �U�$�����:&eY�EUy�J�7	�a����'����Ȗ�Y�B�"�bV"��֫{X։im�,	"x~��h��镲��O7G[~�����˯nw�~P���񋗷7���nNNw�~l��~���gG7����g�|��_����ۏO�=E~���U�y����b3|����4�І�W��f���^�� �Q��V�=	��R4!)�#^�g��0MC<����J�)�l9����� ��L��R�G�Ti*K�zW�x˳��fzP�9�2P�+$�Xo�)��e)=�,�j����X^;����DV95��zK�DJ��Q�#�����e�ιPƱ��U�9���B���{��
��P�$�!Cđ��1��|������/����D���.Y�@M�6�R%�HMef�yRL������Qy�A��i��R;R^���/e�R&�r�O�-���c_bf�����h������G�>���F�:v-�l�&�U���6�p����´�߹���W	RZ0KL3۔�N�Hġ�}���2}�lG���E�ߴ|(�#����c��D֨"��f�T��9D���M�B�ģ�R˨��H\ܗ>pw%,�p��AƄ����r�j��,>3\�{AS�ɻ�*"� 
yK3�󮗒Ѕ��@����DF?Y�1#��U��S�û
p�4c�Ol��#+����Y�nT��!I��H�#�=���s!0Mם-OG�B���jk&d+w!���@�ҝ ��@aÈ���2�G��d�t��QSKun����z���!�w��^�
�0$$e��w�́�����J�S����]8�X@V���<<��^�ӑb�{�������r��S��[�8#n�v��IQ@�ė5<��k.X"K�F��X�0��#��Xy�CͲvYVV���7@���2�CKܵp�ւWB|�J��#��z��*ۦl�+�啫��I�l6/^}�<yG�����S��o���l%U/|/+���/�gk
��`��L��ֺ���_,�p4&k��җ2C�|MS�/E��*��˖����@�%��!�|��ķ���x�Y
,�@m�rg.�8��3�*���Ӵ|�p��J»p�yʬ^��Y|
�@��L^_4Y�Dj�[�ʑ[�H��l6�J,���X���OD�rZ J��{f}["D��Մ���B~j��lӴ��&��/�N�GP�ϲ ���A1<q qKVS�k]	o��v&)�#�`YRS��Ѵ��Z)K��<�x6�bF�kB^w`�TTG`S.Ƅ���9��t�f�mA�l"��2H�CCf���G�/�[jG���6�<|��U��y�B1�V	_�D�rZL9KA��5o�r oiG��G������Y`#YF��8��1��J�z�WR��9��j�<>��-�Mv_���]���aڲ��N:�'5��+�W��q�!qX��ˢ�q�h�]������a�[@��8����zM����Ip،�V
"0<[�˩���@�yƴdR�C�W�d+����d�C0L4��
,"�jç)��������x
���|CV���l�,��[�xx��,D�,Τ�
R#���&����+w�    IDAT�'�ǟ�ʒ��R;̂4����)0H��+�!�QzI�?��v'�Zq�!���*)6�Է��!��m�����|n�9�4yF�IС0��˜���#�
�K1OV@�^᳋���/��RiY�z�@)A�
��%����{�tV�_�R<dBHK>eH�1�B���'�γfV�6:�� �U84�@K�� U#q��][[���T�2٥���E�+g�K������j1� ��G�q�L�3��M�}�� +W(`8@
�w�߇���֚W�l��fk]� �U��ߏ*�?�dk-�ɔ�t�,�ϐͬ�w�N�R�o`���U +k~�o�-3 >OM�?��>o��N߻�Rp���@��,AP(UA����5A1r���25){K�<C`��p�.���t\�«��[��]���Y�0n^\^n����������ɟ}���?9y���ũw��Nnln�~�{w��W(�x�	�^x���GN�'o|�rw�u��4��r%�ⶽ�>���ى7`f���4ڦ�ڠ���E1��R��1H��5`|��i)�P��:��R���8���l�)	'�3�/��f�PP�.��/\�J�#�H�mG\��Ei�Ԑ�+��'���%&�?-<A>f�E��Yz&T�c�:δn-q��׋2ޒHR&5��p-��~�U`�j�@���7mjuLDS �-_+�UI����/%����}A�%>5%���b�v��U�����P-A��Uy�8�;���~��;�>a��vrxp��J,O�>��]]�-M�`}p}��������f���kGǛG�?�k���ڟ����l�?}��������W�?V���}ϵ��=������Z�b�쟕�yvz�� ���??K�7���!2���?�.5>��T���� ��L��QFM/ŀ�7�B8�)�:��%%Fv���^��)3��e���N���г�ޖȂ���i2U4
�ڞ�T�zu���n}i��Q_S:rK�8P-h��a*�'>�� �Fs'���,�Ȕ� ��!�EN�T@�H8�����r��׹�6�+w�>tC�0���2pg��&��a�dd�3s�k��)u���<Ϊ�ڗM��3��^Z��Ph�>��0Z}�	n`4KoR7X]�Z�	��6�Ш���O۔�!3a7�,�
:[�h8:R+���Qt�p��ɛG��#`z�7��h�@��<�I�=vDF56� �E����� p3���3�0c$��&�l��u(}:!�kr�: �K;u��B��6&ok����,�p��5��4��� �'�ļ�^8�\�1!o�f���m��uI�Q)$BA %0�ڤ��rW"@k$H q�1�p�Z��Ju��cI��!��[\A%t(K�R��@U�I!��Z���d�	�:a-F�2�d�8�i:v7�*)R����@Yd��
M(P��kǔx�ׂ�I0��+�1B���~e��v�ä,� ˈ -�����#�1�8�M
G�+�k�� KDY�3��́�-8:�#������_�w[��?��=p�*�!ѼV�RN�G+�Q}�V6E��Edm�/*k�D��lWJ	�%`V[�S@M�Y&�L�y�azэ#6�.^)��@9� ���'"�+��޾�{�T����Q(4�	����<{Mq�����h�[J��}�jYg�c����H~������S�*d�%���qq ��g�#�-�8�Gd-e���R��+������h�9�<�r^��/;�m)�S���� ^6�� YY�E�����СM9f�	�e�BR�)�R�0���J�Rvt�����QK�M��!��2��L�7*�Yb�u� -���Z�ȕ �ƏE�#4��[[cj�2�%N)��<�8���".V{�r@J�bkϻ�W-梔Bo9U�$E�;�S�l`�^c�� ��b)|��R�u���r��H�^3a�f)Ր���wP�J�J �Q��Z>2q"��-�T]�1$��������ed)���O��-�h�6�R��F�e��L�I-B K�$&O\JI��(O�����Y��A�9��	�OS��B����-��L$2&K3�
�M 3%b��@-|@��`@)/j�"ĩi�>Sa|)�����I�e�ǎ@aKH�Z׷�!�d�Ԃ�{�1Ƿ#�2����a[��h >&B`]���e>��*H����h�r�2��lى�L�PIw�l�Ur9@K���LU>��p��Z�#%��GK?�F��:0��x%!|#�`�)�6a��J���T�&���ԥ%�h���Z�j�czE�x�;�Sߖ)�6��x_V�e������(G��#��u�P [�gR��8�#}��h�7O��v��F��ɔ�1-A��>G�,��i0)1�(��y��դ�LV�q-*"g�YR����h<<�l5�����z�(	��R�x8#�/c�_zd"h�1ıw�@��W>A�RJčT9��k*Y���;����"�Lu�,O�yԊͰ&�Qe}�����B1��
��J���ׅ�Nj�״ʕ�q:�!�D�AU|s� N���&�s� �T�B���\
��{��6�بm�W�@���}W����8���>!M�c �i�	�-�J��.���)^
�[Q4WY�M�	-�u�%+�#h<1D�U%��f��g����<�C3�ZH��-��[E�9��������'O�{�=[�ncLUD��M�%��������?�s}{q�ٓ��`��ÿz��o~������kg��'_|y��/�_lϼ�����㳇_m�_������~��藇�c���������\�/���Ó午��3�t,˞כ(��9@��؋i�'C��[�#�eG�W�%hS,HP`)���Fy�,��#���K5�	�?)�,�(��i2j�q �,a%��ZR��LU3W�l��<&��d��-�:����x��3���NJ�L�����kHٞjg)`��� Z��@�:3�"��/V�u���ňÁy��N^y��!�Ϭ]d�,>D�`�RbS�}��Pd眧5���J(Pk��-��Ҩ
'FV��W,x뭷<$�k��OO���>�����Ƀ�����o��/��e��Lo�o���||�����?�y|s�_�xq����c����?y��:����zws���7������p��n����ֲ��>�A�Ñ��,�G�@�-�rHwQO��R,Mp�Zx3\!ǌ�d�]|�\~�B/�� ��}��s�� �^'��F˸�A\��=����AԾ��d�`ɒ�Vs.�=�#��;5��w|pKݩU�Ĺ[�3����4�h�,y1�jz	h6���:�������������oC:=��V�&~H-M7�~>��T�r��Gu��1�g=#�6��AF��(q�Z؂@�*Y|�"@lD�	wO�BL7Z��Z%���
�SS�	GSh���]����텠Gmq����;���]z(�F��3�jǄ�:�Em�Z�}��X����r1^S�8��](L��0��<4�e{	`�6��]d@]���Q�%\73���.�l�֎��t��N�,M��1뢝r�P��l��@�� '>����J	М�~��5 Z}��{�L�.q�Z[:�RN@`kk��<�)}�����P�<�#�!�t��#}��;mKj|A�3�J�#��/&D,�1C�lG
�J.Wǲs��&��@9����i�͘|j	����+%�GSN�,Z37�����6)R#
��h>�$�܅���8M�J��^��9Z~�������r�V=�u��G6o76�(��7����T�2��Qx�B�@�&5t�����3�%�Cp�*T.V(n�Md���e�@JI{7$*�Te�XKHO8�#�K�\-o��"�S��`M5�]����~4Y����	��� v��g�;d��cZ:/����]�D�ldqO͒U^�f恍À�j��5B)�d-+I_L�gq&%`]���ÛM!D�g��>;�#�Z���Zd`�J������!���!��j������Ԋ���1I��)a	
�
���^���U"�W.H(`dYSAĥ��%�FM'��)�_���!�����~y�§����K�eGg�.�J���H��`�� �ƴ�k��O8��f����iA�U�K������v�D�sh˖#�>�=�{�@�D'+���muhīM�R�dn�T�8��JuPq�MK�N@���5���4��I��7U'�E�%���$XS6�-�Xm�RG�m����x�#9_I��|�:�;8��i�#���C<�3�A��$)�>N�+@ �=��� o�'pR�AĬ�����_�4�V��B��B��O!�10��fxq���+�a[V�B�lH�>r�fk�Fj �r�]���
��;gӶ��fR]��ENm�R�R?D�x�Ku��!<�Hp������J�GVj���G�S<�@1�����R8@���xG'%`+��Rvw?PhȤ訢�D� �}M8�f���[Rh�fϴe1�Ny��-C;��5s�X���)EM��,)�� 2[GX^z!H���!��v �IKwPb�J���$��K���h �c)��t)+o��.�a���!S^	NͲ�o)�A�oI�B�|H�b�AcR��X�v��0�R�S��d��b����l�
���B����њ\\�x��Y:[%-GV��d#%�=��>|���"?U�\S^ʄ�+�76���[4$o���/��1xW��'1r�([,G�('�y1	��٣�i�7k��0��o�2�&����3FR���:�{>��]̒U%�oY�Á����/0��0g����@q�c ����SH'�7���Vo:L�����B�c���9q�i�eyWh)HP��cT(�܁�k�Xn���nT'lkh6��R� �[:��p1M�n���wvG�T��Q�>:����}��~��k6g�ǧG[��������|�=97�n����ћo�=8��խo�u�n��:<����������i0�I�.� �/`N�~�;+q�j;1fg�C��J 8��	�����}q1>�ࠔti�G�L�3�&������7jJ�o<)K1f8�Yj'hG���+ܲ��;��@�,Y��?�k�AY�8I)t�͑�a�ŷt��Jww��h�����;j�J��o������B���&��l`�]m�B2f���X�.���T.�X",�6)�Q !h3P�l�����݉3L��'���)O��
�w�w~���]xxr����7�^���˯�/�mN_��������[�׻S�hs�-ӯΟ�<�x����O��m������s� ���ٱ�)~6(p�������	�u�<�W^��;�|�v�P�Q�w�Y��k�`)vJ�����FB�����h>`�"}p����ⴰ+�DՒ�7��تfM�)��c{p|4�g��󖪔#C�����pD3�@8���%�ZKYf;�j��z"��͖����Xδ1�J�>g%�@��O��5���q���ұ~��>{����iU�o��o���+D�!���y;�B/uԺ]���ĚJyf_y"��� �"���"U־�sPe_<#[�����q��H��!��h�O!�����qY�ε��҄�:I^��	��#�P�vԔcR�1e����Ȯ���顔�B}�e��lz�-���ˊ�TYC6*�)�/�+�[��(L�#rb8������5�Z��땦�_J���`�_9��~�I�x3�5�AY�,RP�2��-1Y�B�U�ƀ��\l6KAօ�b�2�f�����Z˔� �[Q#�9U��,� ��t7�S���r1��+��i�*Dch�ӫ�-���Vh٨4U1����$��Ӂc*�btd!:��@	0?���p1�<����L������va�8��<Q�hJd�6��CAS�e%��B�a���nNO�}��f�����n�/���57���v��SqG쮮_,?�A�1 Y����t#4���,�Te6�)�Mã�q����@ac ����=q�b�#vJ<��t��F*}RRuG�в���R�����AdX�2�L;��Qc�tx^5�rd�K��	��Γ�"�<���u_�!b"<_s)���q�N��!RcMH�ɑ� �C�QS�n�8ʇ�'�/�'RJm���wV8ʫm`L%��A�
��<j�E��IZj$n/Y󐊃DƉ,6�{F�O�;�f�3���v�q��-2q&.H-�pHY�ن [HÄ��&��YM�/ei�8dDl�'�C�U��W,�+���9q%�S��Q�,���lg�{<�Ť��i��Z`�A��>�O��.jG��fp&ݍq�ЦQ�P �R@�X��夔��������=uH�����U_:>�E����X6j|^�?2�fW(.5�,Y82<d� ױ�1-SD�#TGjb�hb�iQL4��H���b��{�&I9��h&h�9��#L� �g�t����+���Y&�x�WU��!��"R�R��4�c����~��$)�m`q3τ��j�VJ-fϙ@V
��t��#��O-�*��q�X�ʮͯ
�C"����e_�!R洤@6AU,MH�I�1�	�i���L����9�rF
��|V!� �����G 2�ZK3�����
q`�Ն��{��eM[�t�j��b �e1�μ�x?&��I����|48�恈c�suf�D D,l�	G謀�A�YF+�i��Ӕ��#��ŏcI����>L�p�0&��4Z&��x�U�D��锅SS��h=^������2�ĤX�i0%I��� �^�
��XfJ��K���Y	��	�Z� Č��Zx/I�����k�<��B`u���RI�pf�b)A�I:�
ۣ^s-ЦE�x��{���U�s򐘂�ua�'���]�B� �_M�]��{�dUŬ�Qō���&屐`-tG�/ S��eS[]�8�R�=�*�W8�׺����/�V*5�N�Z�W�f׼��h�$�S"��R�l��=:�X�d]�1���_)KJ�6�,5����ײ���a�|cC�mp�gΆ��!�N�.���@>1<D/���	��,���f*H�!x�7������w��Kn��_�m����t�٩�۫�O?����>=y��ܧ��_��]\��~x������?<8<��x
���]���==�承`�=9~�[�:����G���l�x��s������Ӈ�����Y�&�l٨�6Uw���y�9�K�Lx�((�����t����\,e9�k~)ab%���"�gR8<8��H�ҙ��T�L��(O䕠I&��'��� �GEptJ�x���|[��j�ߎ�E˺O���J��3��;3>�ƃ7����[�M%gCS.�'�ϨS�R���)o*�
hs�@�6�j��Z�l��
��/�t�D��
���e���^Sx"�Rś����6��~�������n������R�򛈻����8�+��?�p��u��m�ۣ��7�}��K}����n~������?����>�K��O�~�ͯ���>��~�ÿ�x��`�|�6��xO>n ��:�R�,�[��x��Y��k�y
���8�Ѵ� ��,hBGd���Jl�����	�gs�P����X^/r���b5J�6GS����D*�X�%�����{��i\.���G`�v�@���#�;�!�5cTMK}��<g!0XUhD�b����1���/�����e�oa���������/�����;?D�M�%��^���$���-|؄�ԝ�	O����:�R���I��ߒBK��5�����*[�p�>fdB�B-t�ܴM���o�f@v�|�k�l�l�e�;�����?�K�_1�;�&e-|��V����/9��s��w#��:��+�����9�U��e^����ѐ�a,C�m���
b��+}��N*&q)��UXJP���T%@Ï_\	�.U�zշ����]�o$Y���Uс`Rc����!��G
"f�f ;%�R�8MH\
"+�랾¤��C��q������r�!�/ւWh	W"E��r- �o��    IDAT�����i��|߂0�@���b� ��t�S��B�^��;��r%����T�2��-����R@%t U��x�ab��2���e�]!U �֒�K5 �N8�����;K-�ۓM?Ex��X�%M���fw{���+O�v'G�;������Hi�9U�z���o(P�QX�1��t���G��,YcO��4Uޖu��CGY/�Q�0C�J�ݕ���y%������������^��Sy�
1=s"{�%�'�}u���y�Fr8M"�0Y��� �Q�)&�T�q�l��tg���)�u��W�}�`-��7� ��#�AA��i9W�����k��3�~#�X[@��dv�`���4F���R9Z��z9�}��H����t0��z�j?Dy��ͯJ��jJ�� _v�3[#�2��t��Tλ�b[H�B�Laj��A0���-�2�M�o��6K_J\�vS,��yF�F^��rRpB��N��v�Q���D�[����5H8�T�&�T���
!lո����i��<r�%�,G���,�������#�� k0
M"�0�RӨa�����D*���D�\��3���{�ll�I!Ȋln�R�Y���h��u4��@�l�ӚZU��X!/2�8eMb�<	��p��*̯�2)����S@`�N@��/nN
�ƛ-G���%�Y$�h�c�	el�bq�<�G�֋~Eب8��R�^V`U���
�R�c�����&G`)D�t��8���G�L� �D�eY�*q��ʋ~�:"0�eߜ�5�M�C���)V4y�"��t��v���z��9:��S�M��a3v�f�cx�����+kH�N�GPR�td@��@R|�^-�M<�)�#�(�01��ɳqBd
�S���l�ʁq��C�2"�u�mD��˄l��f~R�k'�y?51B��9#!�����5swD-�\a����
 p%q mhk�-�m|h�J�<�p�1�L� k2M-�#��2��8٘�(���#+D�� 6T�~h`�y⫊S�%ñd-*_ớ��sC�&�8Mxgؾ��G6r{���0���̎�c��/ ���Ʒ?ޅ{�w~��_�ujB��R Qh�:�iD�#ũ�f�y_!3@�)�Z�l�ld��+5R�b4&�������8��z�_�6��N�w�:6I�|�$�����[�U	���`&��^9"8ZY�����N$e133��{m8��޲s�p ����7���l���,���^�L����F����a=��^��f���}�r6?e�@H���b�f$��w���w}�?�Xd{߀�o�}�n�Lw����G����yy�y�}��3ol}�����O���7~���W�����~��W�����?�ʣ�ϼ�p�/�<|����ó�p&��mǨ��*@�,���
l�q�D���TY`%dh�<��
J��d-C��$��T-�!L����� K@��Ӳ����"����ի�Rpq4>B��V�i�xd���R��$��8?C��;�^�f_ŖsJ��O�Q�rD���/��
�;޶����u��i<YS�Y��@1Y"�Tk6�����f@� �g�X���R�6���{C`��kQ_M}��G:X盙&0����'}�����)ȇD>�x�U^]=��k.����;���������g��<9}t}uq����G�^����n/������x���_������Ň����~��ɓ/n}�y����O��?�\�Y�?~�������w�5g��_�y��x��<y����v���;�v>�+<A�A���tP-��E*K��V'&��T��@�x���#\��4��F@"��^>>T�ƚ��t��7A�e�[}��Ra���A�A�����9�����4h��z���#i*O����{q��&�T
��y��aj�i*��d�RV����7W�{���G�4�r��ܝpw��W�]�I�������ħn>�����=���ӷ_1����o�JLe6ʦ��L��΃��f��3&�O��z��忺kQ_S>��	)3 &�*K�;�b�@\>Y%�:7�1�1�_��l��-P�O�v_A�Ϝ��5E��@:.3 ��3Q%�����	��)-7�z�1�81:0d�e{��Mn0|�]-�^)�����J`:�y���+�\-��*D���Ɠ� �Ԣ��kZ�v�)�R�
qt�I�ɪ�I
b�qfZA����,����	l���_�:pUhL��(LG����RZ[���t�.nc��r����&[S�8�
S�w�鋙jy8Y�S�؝� %�T��}ɲ��ْ'���[T�Hs"�����B�Mh��
���� lk3�H
�i�n?���A	�C@5 �����B��OV�r�����ڟ�?�].�o�l������W�
�}���������Z�7W�/�O��o��&����X�Z����];�e��v��L�x�+6�:��X�K�t"�m�}Y��i0��v�-�/^^�<?���^_zx�W�l��F��=����w`��.�M/C�����q���[t�e7a[��-����1X���@��mxgn���9XRA�pϥ��� ݷm�k��︴�Qiv�K�G�9|:Z�&�����uo=��ǹ糪���d� �-˔,�se`�>��/0�6�H���A�$EQ<HM��u>�o�:�CO\D���O����YU��U�m$q"�v�n-K]��l����JBҩKqU�f`�y����ץ@,K$�J�SF+��n��rJ�_	���m?�pK��!N��8��BY��唆����/%6��ZH��Fɀ��
�RS��ä�R�P<�3��w>����*:U��̒��5Pa���3-�M)L`Hؾ��B-Y`8�o���ƳJl��Ia�j����<*�c�H	x )%5MY,X�6�A`�"�=����Ue)��S�Q)4)kS�-�i���J!?��b�L�R܄3��e^P�|��p�8~YL���F�~$+�`�,�m����̤�V�6�ZK�-�Dk�۸85��`�V O*|t�,���w�N�g����Y���5ٮH�bU�Z [���e�j����1�bA)��[� �N��H��f�%��#�Tȗm�)��:+K��$�TU8��d�"�G	U@٦
OSM�ZA�!��������yt�}�C�v�b*�G�^��4FK�TA���
-uiw�4g�Z�!���MAn��D g1[��4�r˙!qK%�|Uu2U�n*d
��JǴ8��Z$�>\�2��"Z
J��>�T��PvE�F�+53���8��,���)�M���R`�V��L�)�9�&LsJ:��,�j�$+��,N_L�	 ��D-�{H� �0�� ��]8[|��MB�W:>\	KMв��#�9Uu2��u�Y��\�|�mJ�`~jhuA�E���`{w�u����2��Y��F���FL� 8Y��[6�8~W!��&o$xA���'[_�t�h!	V��A��T���,Y�bR̟��
N���H�h��,�4��H\`��y8����j���w���l�8�nQV�I��S֨�\R�bht��[y���NGw/��^]l<:p�4�S���/1����:�)0-e)%bӊ�X
������^��U�]W���0-����~:R��+�}"�K�^a�rP���'5����eq���m��,�&��<�
b?��2S+�cY l�ClGL�^�U�.^�w˫��jm��x��?�e[�F���r}��[�;zW������9�������������!/7О�H�{����ws��F^_�3�7g���������j��f�^�{����W�G�N�=|���7o	�Jдf�7s�l_L
h0�egRl9������|G-XD7�y��Q��7�IR˧�Y��i�?P�`.�HU��r�WI
!<�a6@A�����v�C��j5�֒U�R*�P,^��R�R����RRfN�5ۯVn��a����+ن�Df�:AGdY�*�Y̧�k��´R�<�K�́��·�D�D�0�cV��H�=�0f
��X�� h���fP�f8Mo�:�Iߒ���S����q������^-��|u���7�O�}���՗_=��/|$��|���ww�|d����qwp�s}w����8��=:_�<yt�����љy}]��ڻ}z�ꛯ>z��G�wOϯ�?x����ͻ�kN���i�C�[K&���sb�"�	�ɥ�d�����yC�����0Y��fU��K��;U1I9Ob���1" ������zqҨb�
)���{J<mI���c�W�/�[*��h`o�锴jO����a��F���3���Z�*�	RТ[D�#�u�PR��e�#0��� +�l*�D*�iک��0�T
�t|ǀl��.�@g���������|���7_�h�r�4>;�m6f�k�&p����;�n&we�����f�Y�rKQ3�Pp�9.�~��/�����Q��$��5B�R�2�bI�.pz4�r睼Z����1B%D���2� �C��ʖ��$e�O>�Đ�+�@Ќ����s�@c Bٜ��f��	�	:�M�c:���?��;�&Q�))�N��!
�m6ߜ<5Min:,O�-��9�8�Rl�
�VL!M�ژ@[~�j7z˝,� 3!)�l�C�ج!��d)��AH��r4��p:R)A|��Dc��o��eb)��0��4	]tA�Y����N٨�F�ߤjW	B#)�����) )4/�N$ç2M�JE��RXڔ���@�n��hLnl'�� ��$E��D��{H����L0��_��	�X�x�iB�r}ƣ��,)��Á4�Z%th���Gd�D숦-�a�/�\�O��w��;��X�9\���n���w�;�w�~S�;דߋ��s�%;7��c�^��~E���Xb�Z���^taڵ}�)L�,�<��j��l�@�)Q��	K��|�;�zq����嫽�ۃ��������ɮ�8\�؈����W7�G{�.����r���<n���KS���Bkg:��X[3�y��<��m�2����|���q�m�ӵZ|3w�Q3|���&)�X
�Tg�R9���2�t�j��"�e��O�q�s!�4�&[,`u\$6"���r�,��p^	\�W��2��t��xj�C*A+��,;M�8���ʻ@@�J���e���ᥴNR�M�2ڔ�;`�~�kS��yV,���XJ�`&��f�<>��J,�'8˶���pH��+�B)V
(N0�6^�hd-�l#s��(.��h�r�mӶ�b�<�tD]����dg�8�����!KřZL�i�����*��Gj��l����!��jѲ��p�x��Պ!�틸e�<�bB�S2���:2:U�<�G
GSV�2j�@Hن�$� `�W�C�H���p���Q XFK����B�pqKH A-H�e���ņ���S@�cɻ��J�h�ć|�R�D*�`.t��]2)�mGU��B��bo��;��!�$���@X"�b�F��M�f�O�d���{���xiD���-�5��X�����������3���Kj��fZFd@x�zt�$�<@U8p�����ӻ`�8�@��'�T4)�Z�IE�����͜T��2Ē	ҏ��Ԫ����"� �] $�K*���l}GD�iHm3ɦб$��;�%�&o;�T�Rh�KYک&�0:�5��)%�ҁ3RJ�8e
٨	0�������oj��8�79�������,k�l��_*�<`}���n:/_}I�~T�$u�+O_�/�!��X���8�,N�R��4�B�3L�٢)�4Cc��>q���j�N\�M~�QY����
G��6	���SB�Ä`�&�C�'���K���������� �&�yfB�i(k������O?���A�q*G`4Y���d�a��~����hz�[J��ٰe�dU��_w�R�k�Ǵ�KĲ�JŤ� )08�O��i��Mثs����3����IM/K
����7UM+�i��uS�*A`�L!Y?iⷬ��8+��� ���*V��)�r��z���yŵF�T��l�Bb�	����߮+��^T�cN8��	�Ev��KYvvT�,��Jښ��A��%�ӎ�]݋c��h���Wm����w�W���xû�>��|�r���{g7w'G'G;�W7/ϟ��z����^�_\./�_���Wgw{�������������g`KSI���1���S��xH��|������c2�c-q���_m�xGfR�A��r,�XV���-���T,-
���]!�$n�����C�&(�n����<���e�R�ƶ4 �8h�@����@�l��&�6+�L�Rخ+��SL�3���6q��L�TNG\��H�D��ZR!h���Sp9�D��������� ��m�R��1�6�����8��f�/A8"�$G�B���/�'1|�7S,W7�_}����?~������d}�|ry��f��K�8}��փ�/��?�[����o����������c/�ޜzBy��[/9��q݋��ÿ�����!c{��[0�R�U�#2�7�<�[��f@�(6�3����I@��&��ΓW'+�3��|1A��@��2�]�'��@_me}Q7?�W5�?�я����X�W�X�Ɩ��X�i $���"Btf/�gs��Ȋ�y��s��ihR�R��/�D9�Y�VH���u�C�42}qRhl�Ԋ�.F2m_TT�#�7�7~�l
�����/��/�����;e���v�+��dC��W�u�^�q���m��Ο7D2�,�YJ�k���̀�7o���NRh�O�؆��.�ji���
�����Z�����nG�}���\k��>����nюG�����[��ϤjjTf4=bu7d��d�J�{7��ڙ�l��v�7G���;��w�R4����4��"봕��X֨������Ay`x�<e{Dc���Hh�j�	4 S��!�����2�p`��# ��4����� )���uo8�7�V8&O$M��I�H1K���"��,U��?#�Ϊ�C��7)d �B`� �q�fCp�(׫ Ç�����+�v�n8���j�a���G@
���R`��Ѕ���K� �,�� ���i-�r�DL.��,����;�f�b-�m&o��3C{�T�$@�!���t�S ��@A��|M^��G˅w}�L�o�<�����wK����73��>Z�#Γ��#ɛ����w�'�g׾�X���zy��Np}�<�Qv���&/�3���S�µc���H[�t�ێF�B�oS�=����Ýۓ�ݓ����Չ�������r�������_����9���5.n��q�w�����rg�?�4��7�L]��gi;j�ؠi���l�w�TbrwAU�p�3Q�˹�-�* �)FӴ8�����deK)@,A41oɧ_U)��"d�q�T��2�&Q�B�U�<^�R��@`u�G_-��0C����\$^�Z�q����'2��+�
L�9y��5��U"k�p
5�}Y�jT%�=M��Ƙ���lR`�vȖ��#�����-2"8b��GK\�M�Ҏ!�6�~�j��d�����T-���rS!�� ��e�D�G�~��5��<<�T8'�������uTh�ʣ�x�t�La:)DK0�I��۠.�]@��(��zb����Ոo�ƶ,5�GTۃ���`����Y�]�"�e~��A��ʖ���<=���ɒqR��`�P9~x"
�l��ȁ�4�e�&��Y��4du�ܲF���0�R�VǑM!)�ԊN�M)w{�L�~��u����_6Z���G
n�v��`���I�.�Zq�8�� J(4�xC���-3��0�쾝��dє4�r�|����ntЪE�]����j����G��6"3�t�)F��0��)e����u/;^y�y�`;���Ԛ�Q�g��G��2�,Cx��y�(NM�l�)��4�Y�%�rd)#��.�6G�ER�h~Z�5��$20H�Y���,sJ,�\�h&$G�\�&H���8bx��:��G��m_���r��,|�BC:dY��75"%��-�7"4�e{QX/�7���    IDAT��[R���*>�<f#�	��ᝪ@m]�D�ŗ�TUP��֨�a2�Z�)�i0�����!$��b#%���Ej#R��Δdb��x����kg��|�jT���Ѵ�GGM.��.A���gow����o���e1A�|SՂ8�j��H���NV%% [U)��5\��%K�����R~�����H�RGȈwt�0�Y���²�L��/�}Q��/���* M"�*+���J�O�Tc�:�vA�fem�E���0�R��J�K?sY2YRK<�}hNO�-�1���_/�z	a��ՔDI6};Y}�,��m�m��a΁�!Gv�ttȂ4łzQ�M���m��^������ ����q�AU�������v=�x������������o�v��ホ��e�O���3�j�v�/�ۻ�ӎV7������;�~��N���n�n�*Zݕ�0��$K}�Lq[.ab��
��K���&�A��x���ө$>&+�����FA!o8ٖ�	F'^�,��w&�)P%��lbYq>�!����vS�8� ސ���׋GHP��UG<}e�|3���Y�7
:��e���~�f��L*���-����x��㗪P�Jv�[N���|��J�(I�2�G *�9���r��fKg�]�q�Z��i��b�&��/��SU!o^��Ǚ��7@}�<7����T�����x�������/��i���Z�__�]�\��v�v��׷g�>�w�Vxus}r��K|s��r�r��������~���o}e|�|����['�{���~�o�x��3> �#��]���[B��>��8��}�g��G�&�t�P���b�s,��l�R��pZ
f��yOǿ����;r��zztĆq�j{
E�Rkx���f]��������7��U��.]�T2Ժڌ�z7�lWAV<�E�NAa:8�y&eP8~�@{���d���8�jjQ�[��K٭ؗ�q% <5�.�`j'e��9�D�4�ʛ���O���G�������=!F��.����%A#�F྘�]HA���Z���g?s!�]6��P��&R�H�,5UZ�2������������L���E\y�����D��@PN��a�&��;�>j)�.�-�u�#1w?ߗdd��!�λ��``R��S�v6��t��FlA���7C��bz���?nw�E�M��I��kG��S�fI���K��e/u�M
� ��@1����5L��y��B��Yd�T5j��� [�q� ���) (��$� �V���L���A���*~�^�UŜ$�G�66A
�g�J�
�PV-����,�f��"��e�B:���a��i˚j�CaC���K�L�#�*M�@�f�+l솄�i ��?M:]���&��1�X�f����d{	O��C�#�2��|Su���Gͦ�ҎH��
m��n0�q�����(�cZ���)��TmT� ���ww��w��y����R�����.��/�g���.��:׽��z�/�W�Z�j�K��E룞{�����4�_�0������HM5�	0[���^��S �����W�뫣���jϗ��[� �������?���ͩ���ݳ� ��������{�����������h�w�v�����_�x������A~��k�\x�j�rW4ܐR����~�瞣<v�
1e��ss���f���*d���e�x�Y�aBbj!�I�+o3uo�|$Q�OB���c	l�)��#��@f�̄�k�U+F��[E�B�l:����K���j��jQyU@�Z��vz����orY��*���mAUCHa�ΐ���7R�����
gY-P�^|�Z6�BFl(���X�T��/���@� ���,*K'��b��,�-n���I��rDJ�U��sHVm6��84L
��5���c���&�RV����K����i�p��K���������Zq"�rU�H)Y{���c81�����0�;"1�� �I�Z��xC�sH�a�+�T����?p[�y�Tŗ����p����AǪ�����l���*?Y'@vj�L�lU����v���L�T�ގ�X�v�8���%"HJ�y��l`��S
�"�G�"����n�شCP��R�DU�����-���:��RkK۬�Rm��lR����os��C��S/��fqM�W�¦�}���Sj�(O�K��h� �F�t3�冣�D�S����D�Պ#�]5:8&n��F�^�?͐,�&&�/[�gtFj4�@���pX�&�O�B��0[n�Q�����3U���w)KA���CFܒG�b�
�&�!�M�С��R��������U'�Z�8��1��M-|K�Z8���C�Z6'�/�C��H��%��yHF�g�d�v�ɦl/��b�L册/��8O�	)O�jC�æ�d�*�<�E 
�K Z�##D�j7:&+�� R�=�G�xLG�R�p�B��
;vj^�lH��*� I��:%�	"���Vҋ9�����O|��3�a���o1�)�Q�e��Sw^j.
<H�J���(4�Fv�r�<DV�����%P�H!3K�W�h��-�uR-��iA��Js9�͜~n�S6���t!✽��5@�Aj���ۄ�M�e�N	Aܦ�V���a1�I ��֔#�e��@(�T����R%��ݩ�US�©V�XJ Ŕ�����	f�/�WGo�<��ë�Ͼ~��_�9��G����������͝_[u}��w������o������7�.�Ο>yq~��[��^���R�/��z��ӗ��.�/���i�� B;�ڵ��lT�8�w�AVU%U��O�.|�8�ѥ�7��� Pᩩ*����p� A�uM!������a(Ђ>k#8⤔�2�d���+ǩ\J ��*������J���#K�����=Z/;���&�6��C����r�hVH�UY_�DHDUGķ�K�#��b8-�c��
�ihNqdHx���pΤa�\���� 3
M[w�E�,;#YvzL�8��x�7}2�|8�vw��/�~s���������ov��{��^��x���Z���w�]�;<8y�����'O>���?|����˗��_]����۝�w���/�����ө�o�y�kѳ��i��h����Rܖ����N'P�]�:���:�Jjg��B0�3x��˛��=��]#���ZFVh#��z��x��'5����9_,k��V�'������DyF+/��ND!f2��6R�M����	6��.'OA�'1C��<�d�w�D��Y�o�)���^�bR�Ʀ�L��R�]*�$�p���Ē�]rL����c���@���?���v����~x3;�>郏sz��x���w����4�^=(S������2L�۠����8D҇�N�m7�{�ۊb��o��0o[�O�&q����Aم7��51�,�7��əw+}��� ��ƤC���R��9y��Ɩ�MUN�ز|�)-�Dӹ�����^'k<s�\js��Cੑ5F>� ���<����X�QbB~i��IA�����8�W���/��ێ���p��*��l�/��e�� b4F��/3�2%R�
 ���᪀e�K�Jf�`M��maT�xqYKd��Bʒ���0�
H��C�8
�M<�ZMg >2e8�X�ډY3;m
�CR�Wޕ�!��LN�^�-�ʺ��qO�8�|L
@H����_�E ht�W�ДP���0#
��m�FE`RD��ǰ�߷�g\ַ��w���{ؾ*�./�����ӗ���ۯ�^��ݗ
?��?�qΣ���G�Զ�=��
�?�y��NX��պQ7.���'�p*�2��c���b_N���Z�w�/�W��g��koo����~ы_sr��{�j����/�_�^�8;��d<S�}
N~����]޳�IӃ�;'��Z�U2WwWm};OM�u�-T_�]hK)fބ�$���J-S��y��"���,JPn������֦#!���"˻Q3_
}}iR�E/$>A}���XaH
�2%|
�
-���Pʨv:��#Sf�0#$KD����� �)�р\3�FSdj_W,d�
��r���i0x;��h�i�t��)�����m~��H|C���&�Ϊ-�M,`�B30��f�bYKAY^�d-�,#�S,P+`S� �~�_�8m�T�
q#r4R�l�������S"�f;=4�l���L9rgRm%���*1��ĒN�dx�}���Qi��:e
L�D0-6��,x[�ΒT��?Y��i�L��6�	�Ex�i#�E}�I�g�9�u��D�y�	�#��P�V#���b%��|�j
�]���f*)f�q��xR��h8l�D
_,H����.pU��H+���M'r�|������Z�)�D*ҙFq� <��[�b��h�J*�q]r��Ϗ�,e#(,phl�0�Z��l#�-�L�fu��C��`H���9�h�m��Ԍ=|Y������L-<��e-#�,E-�1K�,���JhF3�]W�� k)� ���R�4��ѴH��RS��6E��q�V�Pa�4�jYL{��c�@^�|�1M�,p��w�e���.h�J��] Uu��w,��@�&�F5��jQ�>_��j$HgKq�u��*�0�LSUuO�{�]�єI6f"��D��j������<��b8�4 Z7s;x̼%S��'�f�b��RH��ŜiC6EK�9!�֖����S/4���¶7	B���#"��oAI_6e˦"!�W5��e�s�#�1b�Ë�������{3^��#�sY�>��K1�%�`��� �Vy��Ф<�\Pf�5+j�
�Y@s��r?H*��<f}x�|�l$)1�F@LHC�Iծ,g#�WtD~N46^�Tjbf�,��I�.�4�n���l/p�u#�� �r���OR����ѥS_�Dd�ϳz��奌TvN�%�Kd�W#�
� _��I0C���od��\t�S�:�N����ꋣJ9k`)�������;�����>����o�^�u���x���7@Ͻ��?z_^���<8���'��~�����|v��WO���.w|���˕}���������|�]�iTS�hgH[���6n6��|Ƿ���@�u��YNIU4��e��Tu_�ecD6��JF\aR���3};pH���Ͼ*ob��˲����Xv�'hY�
�@U�t�	dm��f�����B6���8!����ٴ��_��>Q�M�i^j�J�@��ѥچ#4���Oh�TKC�f����U��/�6C
�%o]�z�U
XwK'���ZC��g]ZFnf�
I1B6���p�{�KsOv����;_@�nWϾ9�����v�}�/=�._|s��˗/_�no��3{���7u/v߹��ͣ�o��zt���>���?���@��o�{���&nW�_~��z�EB/zE���;)�&4�y��9�SVo?y_���bڋ舌�S\��IV��*g�xG��n$���Ձ�G`�^�&�ˁr_)���L��<��?���?�gk/J� ���u�]��G�Ye��s�{BG�W�A1r��C�J|}E6 ��j�ZwR��FD:V�jq�J�`�T�Zc���F��(�������M���iH"d���F�w3�U9n������j]!Y�<&����6��_����6w�y#��%t�^�k���&�4-`6ǅ��H����|��=�& �}�a� ��[�w�݅R�ѱ��[��YCڎOL����b3@0�&h~�P����nk^�n���9O|=n;7��,;��0���I0��lnV]|�� �#7�y�Qh��D���ω:F��lA�Tb���M�M`���
BR�Q���@��qxs
��F ���<�)��L�x�)وkgYmU�8~q|M.k�8�p��b�����4s�C�
)&n��ix�XK�گ@�ךor1Z1�@`�h,�%_�����0� �4"��x����i�N�|%�xL&��.�wDb���(��T�Z����;Ӵ*ލDJ�̓���@X/1>MK����v�F>�C�$��	�\Vy }�_���K�ͥ�9KL�n������>ܿ><��y�O���z��W�_�|zz}�.��E���;�;8|�{����o��p�X�������ړ���W>u�/X�X��]�*��oj�Vk��F
6�z�`l�m���w���~�7�r�{k�{y����g.�A�]��_���;ٹ޻�����W����ɫ�/.���:���=����e荇'�z�7�����3��r�|���j}���b�v�����3����2�ScFZJ6�
G�A�} �l��=���,�,;�b|K�J�N���T|���g'f�T��ä�VU<� � fp��� YШрM[/'���9C|��2@��NkK���b�V)V<�����mZ48�HUȋY�`NU%@Hjb
p&�]H����#��]��~�pҜ9����0�`So�ሧ�`��@�-��ZA� ������1~RS��m�fˑB����	����l��Y�\ϐ�0Z6U-I��[
��$�œ�P��r>)�&��B)��y ��bbKfY_��d����M��#;Umd[
�yj�oU͖>�l��~�Y�+L�2>0\�T1�e��@:���NL
� �vT�����Z��4��<< R"u_��J�4a7@K����UK��x���)��;ߙ��L�=�1>�^Sb*��(���l̒���L�f"Z�i�J�� ��0�,_g�|g���\д���h-�,ۮ59�����LI�ږ�v��^��q�L�v��_Gd|j�.��bc��3H�?KA�q�Ւ�4s��9=R����¶l:)GD��,\�r ��W�����g��#�0c6@�LDa� ���ɶ�N޲��`9G������FfB��i!� sԉ��8|��%�ݩ�?U!((�j�Gk;�h���p�4��C���/�_P����y�!��I)ɶ��L��C�7D���,[)K&ؖ�bY�blTA[�YR3s�A*,�М<C0'P�XS`&W�C��M.�$���xHcT��ʆ�5���j1G�{r#�\)��r>e�d��j���yzY��T^k�Pq'��0�qR������x/p����p�$E���ģ��5mwLK��IڲeH�4���<#��8&��G/�)�A��+�"U�<�h�Q)fwbߓ�/��!bAR�(7���-C�a����RK��H?c��نI���a��k�L�oi�za�m�Q���7F��0��@Y�� �X��+������M����7m%b ��-�/�C�/���Ȳ�wȝ�@���jo�ss}�CYx~����t���wC�Y���W�muu��=V��f��#��ͥ#|[�=>}��W�o��~���������ޕ�4~��ln� ����g�vm9N��_��#��la����#�͙eG-U�Ө�����8iN����ђ�m��BR<�s�NǙ�P;~1)�M	fjCnl�L(�w�p��Zq�l3�(o�,g����j'��<r_w[.
��'MY8�Q��`��#��R��sȕv��YU�f)�:���bp�i�� �Ӳ�qD Vdi@�9�Z��[���#�b
�Z�)�^*f�l�z��W���|���񞷗-�퓯w|Hb����݋�ӫ�W�ήnw���.��������#���?~��7��嫋_����7����`u��h�ȯ��;y�c"��V���<�x��ἁ"6�'dO>&1?�{+G֨�م�F�2��)�2�3)K�bA
@ǂS��@�<�cz��l>�cN�W@�-ioϗ{��ԉy�R����i�^MR�7�H#y������[�$0ŌD*6�Ӗ��!&��	����q�)��B���0�lȫ��j�33)"�&��DǶ��2�T~�T����L���E0\����y�"+զ�B4^S��P����0��}�6)8���ו3� �Ks�    IDAT`�PV"��A��75]A䎫�D
_w)U�=u�ݬ@��6�2X%��˽k�N\�� �C�P�fu�:���7)f#���I�mTUt~�ӟ�;;u�*tG��M�8�|BT�
������Wَ"��X�!h$�o,dm�kd$L�U����XJ��L!>_\9e���@X1�~�)q�Z ��*�i6Ϥ�Ac��Μ'�BD�_�H���F�͐x�fF���٨�8�By���Y�zu�����J:��4�Qܮ)��91�x&��F�9;x��b G�62���y������!���mv] �pK�/������M��.ڗ�ΤF&�Lvq���4��y���Z�0�d�)<��.�����u79M)�j�+�#+E����o�Sk)6�{\SB����[';��W������~��>����ݟ��<���������lv��?�×Ϟ�����G�|��O~���޵� ��nO���[�ӯ�S�=Wæڗ�����l��v��̎�Qy1�)q;u�,�8�s����ގS;��{p�r|�s{�޹ܿ���W������/�>��ju��B�`�u�׫ã�7�~���_���|�/ݿ���=Rl���z�򿖖�7�.Z3q�j6'	��L�d1M.0���`w�b��	a=��)��@������t�B�Q1�V����X��D�`��BfR�RP_��F�
��P Gk;�9�6g��m��8� S+��T�o�KdK��[�Ɇ��_�G�i���H�q,gS��*���R�M���EK��"���ydMg�NI<�)a�U�y��KmX�"�im$j������c�K����d+�Y��u� ^�Fbct�j*��!.�	�����̉��dUQ�
آ���&`�G�!����:�|L�����U��q"�Z�G�R�BSͲ�Z"��&��l�ʥ,�ب����ZX��p��y�,2��� d��q xVw�h���"&�!���;Uw`~pA��Ys#�b~4h(;[��5@�JzK�M�B��Sw�ٯ@Us�/F`
-���v'&�/�W�Ԧ��u3L�/�p
�Ŗ8K���U%�rA|�}�U�ἥ�^��e×D0U�i�R��TŲ�,}�6(6�r'�Ҝbj�2T�m@Yd�C���Eˀ���Rh���VVIG:���Ȉ+t��
(G�mׁ�j��!D�C�,kx�@f��CK���Z�t
��@*f�B�h�8D�����!ɊS�Sh��X�Ո�T��KEN6�<���l6)|3����](Ip�3y��6&2&Y֜��R���H��f����UV(E_��R���R��M���X���r����Z��N���1jͬ.ȶ�S�rc4m���YY
i����Ok�څt���l/�h�Έ#LG1��qĲ)W��eϨ-!b�� r~D��B��ȉWb_�K����)W�>�� ��q���R�B�*��t ��R�75��ǐ9̲֟/�e:��;b"�����J-p/U�>f?$�1%lY 5�D >@��p�%N|�b{����dd �k)HS�hm���Y:#�f���w��,��"ח�X�y��iӤ ���~u'��w @B� (��ږ^��E���Ў>�l��J�K�fS��+|��(��6��$��} ���ĉ/�?Y/ȸT��^м�*�5��,��DF\��]_�s��{�wWϿ~��7����;Z>�y�{p}��֫?;��ݣ������ս�����Я�:��_*]45�8��߽��=�[�]]/�5�.��m�7o�v�rfk��C(/�^?��#+�,�$�_IU���R�x[�R-)��ĩmbH��"�I� [���,<�w ��8,��`f���U�9�{��j#��ր���F.HD�@���� �7��)�њ!�O0jq4�l����E�#L�Ԫm��B��
S0X�SsN&&�!��TU��v�振��r���^�c�S�Ŏ��.�MDLAJ �t��E�T��& �4���|�b�g� ��xy��N6S�<{y�ǯ��������nuy�ź���÷�_�����[�>|������{/�8����������7O��N��c{��������ztқ}���F�'��x�+~K��ٯڲ7�l�Ͷk%�����5z�l�R���H{�)P��!�).E������w�=����C������i:CL8���>�m5�m��_N>f��R}ϼhO�X{6sP���X=?B�*&5��pL#���%��QP�b��L�>IQF`� ��{#v"���Ȳ|cPӎWi�,�]�;o�y��wKbdc��hL���Cٴֹŗ��i�M�^�p���z�9q|�B��5@-��4D����#�B�c7�^̄�ۧ���[Gy�R��{U/:Ⱥ�j/�@ϴ6�s���կ:�z|�ͺ��F�]H|Rd�u��lh�����XS)1$�F���G�vD��3�b*�툩rb@"8,Y^,�fYM�#�7��5���Dfs��X*�G�DSsv�6_U�F���4-�ĝLS/C*de@jLw��)@+1�r���FR!I��uz��EƗ�|dY`��$<�5Ij��H�� ��aJ��="c���&ơ�3�K�Mk�#E���!���������3��N�l�кM!g��!��5ӓ�Td�p��p�&�3���=���php^U�C B\wU�|���~��U_���olD��kJ�� #��Jّ�xY8�����)D���vN����Ͼ�ß������}�^_��e
w��{�ˇ0�G����[����o��/�zrq�~���z5�g:�a�ó�������ʯ\YF]�ZG���5|�%k�|3�����M
Rfv\��Iy3r�`��~�=zp|s�ju������/���7_|��������Ƈ1}L�U\��Oʛ���������ۻ�g���'�{'G�.7�������zo�/�8�_6o���.�.�!� `�#-Fk��g�3sOS���-�&G`.�y�+)&%@��Ж�ߌt�����{�$��p搉4d�b|j��i"����)(T�#fhI�4jw])����яY���8e��ר�d�oHq�i�Tk�x۬WLUM��TU�o�C�������S��b(Hpz)L���"Ĭ��LS6#�l�QK��j)�.J:
��F��r���`Q&��gp~�FM�Tc�����[2��[��E�m��&|�f���<f>�����%����e�P�p6�v�=����r�;� �tfGM��<�����R���l%�=��#0��Ӕf���UI1L�B��/��R��/@�,ْ�[�m+�e�Z�r)KUMR�pd�
!Rs&����SCC�ǘu�G,�"V�T���T�X2����A
!Y~�.�v���&5˥��F�,RjKsv�O'r'.do<wѤ�u�hj��Պ��ͨ��}a��rʇ����t�(d�4~jpK��+����V���-�~��t�qJ�"���Ų^��v��-r�Qd��) �u8)[����1U�������C�irH�H	� �ϲ�e�H�L�Re� �,g�:�]*7�x`�b�l�u����<���,���
jѲx��5R�V�S^6dp4�w�^�Z��;)]Ĳ��T�>���L��рF�- ��gJ,���B"0�Z��B4Ä�D(�Fj4jSe;�J >f7����)��f�ьg9U��Ԋ[�#�b�jj��#X"Ӵ}d�N�J��>�ZH����ĒO�TŌ#U	"�ƀ������W�#���w����ۚqO����C:�&�'����j�������&���4����+ш���jI�O�1-R@�L�x�i⌦�.��k���l������Z:�
-��R��Qs@���E����Z�2��x��]GP�֎0��ʥ�֏����:��1���R�������'\��PV�Z�N����+������'�x������fPh�0���ZXk�`�F�&��&Mk-��Z�v ^m�pz!�+�����ݻ]~-��˽7>�77O/o?~���l�����������Ά��{���6�V�uYv�{�\���^��:{v����|5��ns�t7�8o�R:�6�4}}� [���A��66�E PRSqH%IR����)�*>�,C�gb�!��7�e����u�D�d� P��Z����l�+�o_�R���5�����zt��V���f *�}�$�)��q�����H������W(`M�<-R�J��x�����b��M��K�Vk3[V�2����*N�+� ���7O�Y�4qtTe9�q,�x��'�9C���w��swy{yz��ū?}�?q��������W:w����yws�w��7��;���}����=��:�����b�^^��_��o�Nx��^~%��o��F�^��M�yF5O�}��JrO����+�n?K&hxD� l��b	�d8D�SV�R0�,���@P��7(�/��#tl����������)�>��^��5	)�n[��&k�h���Ve����T|2�Dl	�k��Ԡ����L,jTw�
M���I%�#��H�)�Ë�)]\6�IXPcbD��oޢ��1��6��Ȓ"�	��;˲�ʵ��҄�`�0S�7?N���pĤ\f>)
�7���T��K�d�����W�^��⋙\g�R�i"��u���|���Gy_�B��q��Ԙ�����/�KcԷ����GS�j�3�sc��oS\5
8��r�͟���鋵�E����l��dc�SY��,�r�k�}(�CV���u����x�`N���F`��D!P`6�5q1�*Y ��d8��
��N
�
���U�)NM�)�v�;
m_ք��W�cJ�@�"5K��,�i`������/��eT%�8����cAfZ��Q�麨�KI>��6�,>+K�9X֨9�p�� J��S����X9S������-�,E'>���Xj��&C�/;��4�h�tjA��v]��<�����j����c�G'�>�x��{x�~�~y��O���ه�~�������j�'.��n����ݛ]��ݭL�;���1�ݞ={�o�}�x����/�wNo_�a�s�ܜ��|�ry��������j�rs�ڣI��]{�Xw��0�l��=�\���Ϋ��vV�;{/^�z���򻗿�ʏ!�"]�����t�R�}���Ϋ���œow^��5����N�}뭣��j�]_�]������=��3�j��_�3���4Ob�T]���Y���h⫆,�u���e���mS���2A������z#s�]��*�/讐mG��if��v4s�*ѝ!0L �(�#He�8mmd�F�5���
�oY)1���mr�(`:�z�FJ#��r��-�!��`]��MR9Z�E���I�� Vk)�7����w�=�IY��y���H8"Zxy6[�"�p%�$�j�M(��W�:�
˦�`��� D�)Q�WUib�#@����	��9�^��y�i.�_�7O.V�&/��R�Y	7*/Ukx-�}7XJ���qT���e�q 1#��&�cpj��Nju*�t>&t,��c��v/q��F�����5:lN)�x���-�b�l��hm�v�XG���
��|�O
�Q%��->��I�W�	�ᑋ�E��!MX��(������9�̯5Z;�|�+���'pz�mS^kN�e{L0���"�dӱ��������f��4���b�9�:�m3MYH:�M��]�UޞV,;}�ˎ� D��b6v�.�j��!�7g�4��`{��8p�RVa~�l8�g��e�q��r�2�h���nx��sZF(@�N,@`�ʥ y�^5�Z@�5F8DIj�R+���^!<��<Y>&)L��x��;�^�������`R���pRsY*�튈)�eu��S� �*���J�u�'I��	S�S�8�#3�WK���;�^b"3~��^jeS�1q�,���R�{��Z��v��`9�1�삊;���h��lBL���X�%�V-�>?��04Y�\��l�$�e�jBLK�-B��׎/5"%��o�vAc�d��$����@��{Y|�� �b��zt���#�;fU�F,�ϊ�G�$\��Ɔ3?����,���x1?���������gr ��ëE�T<Uui`%��F ZVM0�M5c�'N����f�4w8�X�x?k�#�������Mp� �msF�\	S�S��,Y&�we�t)+�RZJ�kԫ+��X1k���^��펦���9>�v-vM+�L�W^/z��GA�*>r��F �x)A��ta��-d���^��B�m��RQ"�_a6�չ.��7)Ww�{�n|���[����O���׿xt����_�使�ُv������Y�-}o�r�j��`�]O��xu~~�z�^��
�wt|us��>�j���;����55��m���cF'� p2��W%`p;�i��-!st
-��)���$Adx��lwr�,pZg*�ff)�m3@{��ͪ�J	��q�J?В��H0{�A�?�7E�ϥ��Ri���e��4���BU�7?��e�Ζ$;�+��9Ԁ�D�H
Ŧ�-u�1ӥ���yA���u#�LC���� 
C�
U9O�����.k'��o����}{GdeDF�D�9'�`���`ZJu�#;��0ţlY�5�(�`A��l���ZV���S.�.lk���J"nH� �������x��3����~�d����V��C&bNbR^�\����G7�^��_>N�\����o�~�٣O���ݷ�~�?x�����e�o���b��۫��ۗ�^\���z-��~�O_�<}y�sus烜7�N�����︻<�<���G$�L�aN���<��u�[l�Z��7m4��1^flA�QP{�hG�m��펗�U�;:Ȝs)]�rjsD�"K1dfZwH�k
���V�_>�g�g��L�S��5��BҵԆ�!l��b)L�J)S"6���S
hqഀTE�@�Y;�.8�u�͍ 
)K�.	��oY�2�k��}�5Z��I���Q{1��~���?���R^v����?�|i�_�M��U@�� h*oH��RF�p �m�0!L���*YFع�K93����ɟ�	�?�j;nk|L��lD�b�N�.� ��"@��W_��R%[I;m�3�*:f�Ӥ���,��&����%oB"8��c;�My|��xd�
���b��A`|A3W�)��<~c��ĪX��Q�:ORR�6!�<��9km8e%�D�k�e<�%�3��ì5�gR"b"�H��s�g]p�DМZ�TΛ�Z�S_MS�wD
5�T� qjam����[��<��`�h�@%8�hN_�#'������ES%+ձHU� �.��#d
����ԋg8NFֲ�N'�I���X-��)h� d1�AM���o^_`���Y�����&d� F�-�a6��_��'�p��2�빳�������û���O?���|�ų����-��ޭ��{����94����C�z�H|���<z����u�;><�5�vs�������ey7���֦o֯c&ir�QMk�n.��R�l�3*����x_��W�Ʒ?��[?�q}sz{q{�����/��=�ۜ�����Y~�������]L��������ܽ�>���˛��~��;�>xt|�wz{f���u��>����}�13��gt��sx2�}����r����g��ա�(G�d�,���,�1���R~b���Dc�p� (O�f�5"3�:b��U��J��!�l��f�]֩M�g��̒�3�	��)t,%s���g{x1�JR#k�|��t\�2�:aq��#�`p�L��R �2�πD�FJ'L'�6$D��^�D�J�-D���Yd�G�6�����)5Q!K�g��.�%2�0��8<p�f��@>\� n�7� >[�#~��茂�L�KKU�P��!�R�!�Bx��J��i�!&(�g�
+�wwT�@��l7��LTH�R�Q B,��;�� w\d��-y���}�X�H{��E4K�8���)	�V��,+�Щ�i+ԫ�Rqd��� ��    IDATMv{�f�¬W�p0�`1?ݧ��I'�b�d��0��Z�jCT��堔0˙0$M�BL�����x�X7|1M6���DЁ��KQV��I�"�-�����O�8���r�x�ȭ��FI	:����J\.�,�,.;�e�#%�Q�f3*r�q�I\��[��\ڿ���B�ډCV�劄��7����Fk�/e>~(�.4��Ly� �D��EL��f	.�u�RU|� [*���JΘ��o$�g�WXmݑ�d�34N9�Z�~%m�*V�㤠D [P_G�w�k�3�4�!�Ck�ZSKJa�<�v8���4�ѩ(`z���ֲf}���:�*A��ZҔZl��+<5��w����V�����ͨ�▪� R� :Z6Cc/[�V_��*�A����pH�jd��H��Z\�x����-��LJ�R�Ϝs�p��vM�F�G�K~�i
A��v
�.`8ȼX�f@(���lB����gJj���,�#�f��s� 7L:R�}c��ܜѤ
�)D�K�w�v��,���(����20�tL�B���,Ş��jm�jW\	��������m��|-��b�}U����o�-)�ߨ��,�����ej�DU�h���xM�OD���	4ā{��}�l`���
���W�+�\��<�U"�"�8��S+�r\;r8�R���~JA�]���:��^<�����w�����~��o<z��?z��������7m.^xS��?��G�����w����������^��Yn	����H�l6�,�NK��dȖ�T��	 ���D�
t��?��?怘f�����7�4�9(�|��G(!��!�l��4j�M�i�^<�1�͆&UI��`~)7����X%pgM�y�f��0�����{�Bp�����j۔v��S�<b�
X�LA��%qKq��eU��M*�7Ϥ�
�0q �	�Z��i
!��Zfx�R͏Ю�eyF!YYK��!3�eY�H��/A\	>�f�r�w�q�&�\�oSy��Wk#''/>��#����g?�����WO�~����'w����_����꓏����/�>�&�竍Opzc�n�u���N�;�y��F��3�.�p�`0OO����nc�ɗ������Gfb�'f���|�t�$U���Z��۬� jTy)K�Dl��``��y]������������}��<K�_B4�����|���I��ڌ%żNޞqf�6f���UA��B`��]�����_�C����rU]d!}i��8���f�2t������M}uє>Zw ���M"R@��E�o�,����]����i6T"�#`h����T�x�}����r�5��_�⋥U[9_��֪u�0dU<){tQdiˍ��*"d��0-<ΐIue]�
������q�25x) �aL�Uu{�S��$�Jf1BH�����-�*�(�DGK`:f��hn`|Ad]�$��o������Ҧ���,�a�pd|&E!DV	2Y1/k���P�!��5EP���F��*-�W�۩T�8�MٶC'AЅK����*�,KAP*� �H��d+�T#hT�F5kＪb�L,��Ґ��,�R�Z"R=R�Y
��cqWH�헒ESY
��T�r' a���`]M�H�3#@�K���L�Rh��ٕ��`6� �5)8�� N�@�ٖSh$�71m���3����������_�<���;>�ۿu��.�_��M��姐|'�9�i�o�������žٿ���/no�?�އ�@=8>�>�~y����������W_e^�f�j����p��e�"����ZƼ����m�˧H�;��*�=_}��g������ԧK���V�v�U����[���ҋ��mn����廏7�s|�o7�6r}�{�w|q)~uqysx䫳��I���l�v],��/�� ��_����y�8�y��	�O�ӵ>Sȓ��B�?���*L�.�n�Lk��I14)� �<�pq�x��
�_yU�"��p���X��!82قi';MY;�9L�a�&�N˘����2� '�,�z�4�6G��xU�'�`ͣog�N�|34�<D*�Ų��Vy����)NJ0�a�EHv�p"��{�q"�-N��M`
8�q���ҙ��}Y�^w^^�Hb�BO�ɷ4��x�<d���HT��St��f��c�@hTڐĥ�G�-ү���FӺ���Zq��
��Ȃ<d��K&�ehⲖ	��rYc`��Z��rM�P [�����<�%�5�$�0��M����#��e?R+�O!���C����")x6�nI��k�[��Ӎ$�(�Sֲy��}�0L��8��j����*��,0N��G$B-�n�pK���o�@q�*�m�m8���?���[2���A�ǲZUe��8�1�8Z�Ri�J��p^��($�O��	��0�v�gG��� ��l!��c��F���Վ�
�r�f�t���$%�0�v��(S�Vv���0�Dt1�XI���:q���L@S!� I��%�L�y��iH`�+,�Snk�
�6�ƛ�ln���,6C�
il���xA��U���)e%�$q3V�<�� hR�R�
�%�%h*Zk��q�߉!dyAvb�dSn��<dh�`"���1��p��2�Q�ӱD��Ѷ�D�X׷�� H	�',�[�}��Qm{;��<`���C�%%۾Z�<��_��7�� G0V��3Yx:�G�g�y�h�u����/�KFn�j�@�UxfxV_ۙr�EK-qHG$KG��Q��]�����뮤*�	��F�P/|W�J�w�(�Sh�f)6�*���N���q�L���U��,�N��8q��;�!7��xNɅ����<eՖ��i��^Y]����>���
����^�;YʞR~��V�O��S	5^ֲ�3�I�T�μ��@d�Z,�צj��ņa�6��p;�Z�w��`��T�!>`���i��Dt~�WV^]�����'O�z���k�� ���;?8�?���l�'�����������ur���j�������������������#�3t��S��Mn�x8o|>p��)A�8M�Zʘ�q�Ө����0c0R��2�/�M�#+Χ�SI䲁��X��;�^R�rx1&�ir�~:�c׶�� 6%�~^=�K"����T����<����K��A��I�O��J$~R�5@���y���Y��YdcXFPh	�'eixYM +F�p�B��ȧ�����-y�A]bZ214���%h~%.C�$^�����!+���2Z"@?�p||�������W� �O���ųӗO��??�߳o�Ο_��=�����>;߹9|�h���O|�uv;�-?3a6O2������]��,�v���+��x
��C��w/u���HJxϊnڎN���Ѵ�w�|)%s��0���PЎ���0ZU@O�<Ώ~�#���㏟<y�Oڋ^�X.�2��4�� ue��!PT�׉oy)� �*�ĔjY�!d�@7ʴ�.��F�U�D|�q���M��WK�)�e1� 5B�>��|~ei�fSХ' ��?�_iL��_����<]	-�zXL
�X��C#Մ�/�r�bC�u���/[���r�Z@l��.n�Ɠ��fx�2��/�A#oT���?��A���7W��B"��#�A�-��ӟ����� �� ���QY�%�u�R#�Ⱥ�ٲ�C�<���+�ߒO��B�2���g���l�զ�i�cб�D�Zǈ��eK:
�Ě� �rYq��×bIa��&�(��ė� ��T"t�l��1�ǡPSG�C�,v#��h�C Ay��1��
�G�Lk)+n�BjD�N�S��#��Ԣ�)�1��cU����] ���mǖ���j3#��]�-��	��
���L���)��J9v�W"nG|��d"M�rU��ȵ�x�ͧ ��0�Rmd-]..�؄F�(@KYKq �T���o � r"�ݓ�ZfU��������]��_ۺws~��ۧ�NOμ�p���>b���|̑�w#vo��<��l�mM�-������ˋ�����w��x����ӽ]_��E���}E{����������Ռ�nZ�i�E`�fv�Zڬ�M�7���ӌ��������^qyv����=�ڿ�A�v6��;77���/"�\AF��QO��v����>�I��f���7'_�u���������A�^��y�֦���k*O��0v���l�i!]�w�m]�|�Ds7v�֢�;��[,ŕ�5��*4X'�BL������Aĥd�2:��
ӯňx*s6�Q�J���
���H�����1e��l1�R�ʐY�]2#�,?�B���o3���v �Ȧ ����x�|82�^G�,gl��-@�.D.@`��!�:��L��R�[E�Z`��3} P��YH�RL<3K�Bp��|�i -� ����]��n~��-h�!X�+�}�D
��J�?������ 2����跄'k�6Rk~������13������?}['+vb=L&A���$��5�,D��^�v$k�G�@��'�i�'/ߓ�4�uݧֲ����L!P0^�i*��d�?���,�-c�Yyۦxhe�Y���<f��eY�r)���@S�<}%��*>�
܃�D�o���R�XY~���]�f䛡���� ��i��"ĩ�� d�8�,үB:e�&_�\���p��ѨE�������O�N���o��BYAݓ�Y�ͼ%�*&�K=:,�,U�ě�$Re#+�f�2�%i�+�D��+�B�R�@U��mh��9	�,�2����D2Kۏ�Ȑ�l��4M�6"po�Γ>N�	��2�T%!1۬x�p�`�jg��k'E�����#(`t�%6�b���8<�8��XVk%��8AK�a��#���%5�Zx�y�H�8+n����Na&�e��!bA;�8�3��R�k-�
NMi��B�dh�9�@×M�6�HyUT(n���Z%��M�"<��P�]UG�����u,Iũ\	p4��q�\�>��\p�<)��U�Ŗ�ͧI��!�e�,U�����L?&$e�t�R(N����S
rwc����'K6�-��esD��";Y�љ�y&B:�1��] F�>��LvZX��d@�L���#���X�q�Z(agB���^���e�6�/ߌ�C�t��!t0C�;�?��?�#�^�E	�,ܹ!ęj�"�Ǔ��7���[� ��	3��0�59O����|3'e<c ������p����k���<~����/��Ǘ����(���������g���ٹ�?��'�7�����7g;'W��gW�;�{��?\����5vc�e�}���g] Ch�-e<�ٮ�qV$���;�n�)_6��}(�%�f��0\�S�������S�&D�T�e�-�pX1��XJk�7pd������d)ˌ�S�; B�P:"����:CS�8�����vh�)�qY̖
D�JH%O�@��XUg��l��j��G	�P�$>�p��fc#4� $$��,G���חoTL�\��;�̑��;�	���ޗ�3:���do�<"|�n��Һ�|��_�\��^�ޞ_,��8zv�����������ݳ�~G����ƣۻ#�ѣ��G�{@Gϟ�s��%&�����ڛ�����l�^�k�j�w`���Ŝ0�����96O�&TY��?\��q��ie�%b/Bpl��������GyΐJ��`�m����M�9���@��1og�c>޹�B�g-վ�t�:�����#�0�<MUR�}I��8�*���	|�k�{��m$&�Bc�IM�,eYW�<�88'�ﰅ�D�cN�����;FN�1�K�c:+׃�{��J��9[��MK�[��fNK)�FZ��	b�Tw�N��jZ����tQ"��f�WBMe$���KD�O��;
�z����>����N bk���&^����O>�ľ,1��5�s ��6!BY�\�	�G`������Tg��ҡy׹�5f�G����B�� ^G��*sJA�4��m3㤆c�[��aż���l�%�jyDP��6���ZҤ����+G�e@�<�|�],���`�#��$�NO�Q�:�@U��Rn*YK��� GKg�p�6^[�\�����u�����s�|�hb&ƌ\�4���R�3��r�͍�s����J��F�.�s��� ��8%�ɚ�Ԝ�e4A#����P!��x�˺*�IP��w��Fy��"��Ko��b��6.��kg9�D;�� @E��~#����7_<��ߟ~{���g}���`��v��p�z��y��ջ����N����;�>�y�{�9�����ý��pq|�y�დۋ�ib���uw����1�9�D�`|��9m_����(e~V�77��
oT��h�����Ͽ|�'/w�	���]I�v��/��/"������7/}��ߴ�_�N�NOn�6��v���xC����G~�D���ef�Hy�����鹺�Ad���}�2������bk����;
�&ň�� m��@�'adw��^���W�*|Hx�	j�-�.�@�8m� N��z�J�J���&����� �6Hg�\�l��<�����/KY�,��0�����t���T.�6_�̐�E���^�q��M�IQ~ʪ�����"��R:��	V��tA�JA���_�]X#�j1!�Ty̐��F+�f�GS�3)�ݜ1�R�L�&Ʃ�R�ٲ�F�V*��1-�f+!$OS\�����Y�R4��\��S!0�ZL#x����M�%k3�9�p6�%|�j�)ڨ�ul���{2��K��;��ʊi6C����]#%�)�N1\PU�p�A�UE�U!��y,Y��P�<�-�+�lq*YZn=$ţS<Y�ZW�� e>�l)Y1��)D(�r_}�"ͬ���Y��#���X\SUFj��#+�0�H�ח�QGs�H��L$�z��n��� ��Y×*�鳖�X
 U�)0��L�eÌ�yFDJ��Ʒ��o�@��ۜ^�ek1R���z v	"O�,Y��!����3��a�J��e�@Z&abO����
��<H�,U���sC�ս��#�)n0��<&D�_�Th�Ϊ��S.;�@m)
ۓ �!X�k!Ff��u3��u�F�u�L���p�vTy1ϖf[���k)�@%ԲN�3��S��FR�N'�Tc�M*�Ł��(Imb`xj��S>)%�mĲ�ʻW��cN �9�%��	��s{oϓ�/&5��F ��ͫ�ȡ��Zō�Txʍ�O�� ]���ډ�0�<k�ZXV�f�8�@�<�&�ֲ��� ������}�����G��P>�4�0[�d
�I�R���xuVη��y���4���i�}���Ia�̑!�Ȫ" IU%f�l6M!�+��k)�4Z���t��0eC�Z�����ھv�[o��oZK)K�	6a��Z��or=�o�6ai��4SN�w�^�մ�t79A��A����)��J�"+fj��[�A���˼�a
	vًKb���}]�4;�j�1�����?����ꋯO�����7������y���˫�7�y�'����<�λ^8x�����o�z����ot�������ϣ���y�^ڝI�c��N���J�[�;.1�t�O�r��1��m�H���ZP
�A��B
�RV*�H1��hȍ���l~�FRUS^<��g��"��U��O���p�im_��g�q�X6@�@���ΎWf("��t�Y��x�`��C� S D�AAU��C��,o6�,[�^w�+�W"��.k���p�4� >�3�%2�X`;Ɋ�m�UM!�i���gZ8-BSUR!��5CY��T_��D ����<���<�{��N��մ!��/M��������������ٞ�E�F�c�#��~ja���Fh/�iDA���Ӛ��?�����l�XkO;��կ��C���{F�,��1�	{�
HD��W+�:�R�pM��	@    IDATښ�wݥL�����٬O
��\� �dњ��)��Ȇ��﫥�������Yy8��D�ĀY3Y��j�	2�J�ȂU��Q�X���fx��/����¥�����sA��f�k�X��*�	i<����I)�p�� Mⶠ�����yu؄΁�eM�uaG�������ľn9w���߼�MH-Ud��t�5d�D��^��5�����§nu״�%����i+��7���72-ݝ��neoj��KQ��X�1�/��!��k)�Ż�?]�i8
����xpRN�%���[�,O?B'��9t5�lS)Th~GY�^U7�Z84YK�U)����p�1Ę�Q�dJ����[�(WhZ&V�ׂח�����v��ďL��eK��D�'H�$��B) �<��J�oɦ���<��lG�n	�I�5
T.`]G4)&`3��ј%C��bLYC��b��Yjv��`���d)�kT�;�ʧdh��/�Q��f���	F����'o��W�v[��y:I�D(  GSb��A\�,h�
���O!8j4U,�4k4-��1d��q����6� )ԥ��,���Ko�bH"�#�#-[X� ����/�~��o/v/w7�\'qE�����������K�����_̼���/?�t{}u~�����xg���ѣko�x/��_8��)��ǉ?,�ɪ!ۈ�����l�nH)CF0L�i��\jW?Dy{��Z�����<����듳�+ͼ�y��i:��D�����0��_.�1�z)�t�ߵ��2���.�n�|����͵߮���N̨f�%�VdY6�eO 8bK���V�V"����K$kS��k�+��/p9���:"�TJ�x]|U��>MUY�-_�b�x"���^@&�)ᷳ$\)�MH:j��ז��8�#�,^j�D`RY3@R���W0)��FR�J�u�S(��8?O�tb*/^�[�8���sŶ��94dY:<��R<�.�G9�UU�6���� �A�	�~)�pw��L�x��F��|L	�,�uR��F�1FʲZ��X��0����z l��V�+Q8��:�4X�����g��'�Ԣ���K5m1YA��|�a�J�����Z@ڠ1�T��{~pu�)�eY�b �8�Rb�d��x�C �D��	\$�v����K
9��� �I����:����@�����CxS/AK-p,c��e�jō-([����雎%�$$M�T�[����g�/��<� Χ̳�
X,@�{���'���-,Z������Z�7�X�!��tiZP�mZ����<�jQy�0+�a����TY�%�˂b��k�����%��E�f�%+&+��HGa[�y���+�X��D*��ƴLM��mY-Ĝ�S��%�3%�J�#ӄ0o���5�8��b"��l~�z�@ͤ�nlAY
ey}��uU
�Q8�v�jO�K� XG~v�}
�,f��)'�R`x�XP-_l�����X�� ��ls5!3�.l���Q�,�E�|���s� W��}��3�4^-rcT��h��U<d"(!R�.�Q�ЌoY��O��l�2DV-o� ,@ӿ�6��lז�EI�[�K�1�E� RV!ĒMmq]xF��J:��%U9D�4�Rsmd���U)��$�v,ӝF'~
����^R@��$��B�2`je!�T�Á���e�F�&A� �6�2�
�=[���o���8��UЌ,�a)�M���x�v$+0�#�7vC�5�K�����ć'��*c0R�1��Kmˊ�D�a�1��)8����ʦ/K��#�(�wj{����^N�e=����
!���x��妣�e3P�꠪2�2�:���0�}�&�b��Ȗ��W�r���k���Q�F�J��Y
��1,��K���i���3C�kRl��?d�x�n�X��<]{o���v���+{G�ܿ<��'����|wsp���y�;?���8�Y���gWO_��`���_����G����sV-;F�=�J ���X��S���`I_6�%��B�%��ѫ��c�I1
�� p��}G�O��hy�[J\)�
�KA_%|�	&��8MShd��%N4�{�q!����`���ɷS��BS"���d��[KP�p�Y�;d- ���	�܈7������|&˔��mp� B24���|Y�� N*B�!<p�)���
���t��v8�G6}>�)��e_��B��t�4_��]�^|{��u¾�yk���>�K��on�=����S�Χ���w�w��qx�{R~�6�ú�޿����ӆt�u!nO>&�$`~���l$�j�|�bz[�UVh�J<�z���h<Q.+�&h�FP#��H�T�\!>D#���+O���d�R&��@'q�Dx˞����Mϭ����*Vfo& ���k��"���2���W�V��Uh��WK��啐� ��G6�u@����A��ԗ�X�0J�������8�R<3	�j���r��0���xS��A;��0{k���>K�o4�#�s�tV`9U�:y���������^�N��9�����QG ��Ҩ�Ӷ�ι�Ǵ��q���?�����5�~���)D3�wR?��ö��ɓ������;�
�$%�Z`�@'@��h��Ev�ȎQ#�!�b�-�4���ǰ\A:��5݁��aR�
�P�.G��+W"�%G0@A]xK�$+�SJ<�ډq(�Lh�+�3���,�Țf��j�SS�Zv���@���}�bē�,��7mL) S�T4��@���G��r�i��P�FjBYU�q4c�a,����&|�,�f�e#Cp����R��T�Ѝ$fR�t�`<%�n��T�pK� NAJI}-k:�vP�3YY�������,�eHq4q֒f�,�%;�R5���
��Y%�v����� ��eR�)Ȫ������+����_���=ǝ���|�=8\��v6�~~������+^o��.�/n/�u�;��m��	|�����G$w���w��t�^�ɭ��oT�E�~U��P>C�8���f�_{�iG{��Ӊue=1� ��.��� ����?�{簯�Ww�pw/�Z��$����{����|��[��o��������^_\_�����Gw{��\������uO����gf��]����M�x�؞��@LK�H}9�D�_�C�߭U
S��v�����I�Ui��b��7����oj�\���'X�
��H*/�fL�F�c�jm*D�6�J������8۱��E\@�r4;(
ÑZK�lL��RN�5�43���tT1Y>e��᷅��kG��]�9)
D��k��*����G(���D�W�wWy8�m�F��K#����T�G��.�Z�I�2��$��W'PR03[6C�bZ�l�n_R�! 	��F,�l|c�ٴ8�k˲u��l8q��ngӏ	�����CK"s�5��,~�@��F��y�b)�D���X0"��9�)kiM�G��g��^��0���01S�6�}^��ֲ,�H���NK��"�68�S�Fj�p`;��M��p䂥���G��.ȧ��3ؗ�j�l�Eh�a��5�d�T#qW�r旍�#0��!Ͳ����Q��s7F�D���^u��ը]�pH��� �MGIHY)U��L�TU<�!# ���+���CҗU���HA�SH��j��&��h�|��$&֨�t $��Zv;5�\̺��U��5	���v�F�x�l���XMǑJ�]�ʍW ǲX��31N��F����a4D�P� ���z�w�)����B"�ó�֎p0Y~K_����_���$�_��-�?^�*��YVPӥ�ʄ'b)�µb)ٮB0	f��\2��8��aj���vT;8��8<�y�G�S�ߙ4�}����9>B�:G l���CT5�{�H"p�[B�ej��� T"@`	���AUK{{�W��¥~����Iav��׷�t)�7db�T�~sNI�gܹ���FH���r] �ҽqe��^�=�,$2_��Քo;c#4|�U~i�Y����X�t�H�g��/�`�HA�!�xl8h@����<���)`啠)шG��!��8�����������z���.��AaLI�k�Z��Ǧ�4*�"�e�-P-�7���r
����v�4���(�#2����ډ�����;���ZG!n0�@|�u���Q���J(���bR�@�|jm�낳}�Y"/Y/�l_���/�5�"-YH/�h�;w����{=��r�W��~��l��ݛ��˯��z9����������#�N��z��~�����7/����q����|������N��ٌ�C&pK�Hvd�3U�Ρc�<x):)Um�����Bj��#���<Z� b�p��)C�
�YUR����(�)�Z>��5Z���2�e4޵6m7���Vq���.�K�{Ns���n�@�F�k*v���6��d��:5� �i<)4��j0�)�A�=L����C�[�eAՒ��q�h�[��&f)kԒW� ��l�·c
 8D�>�� �%�<���%�%"��L. v�5���G���U�ٻ��V��}}R�kh�J4�ʫ�ȶ����a6����w��{�O��y��x���co�>|�;��W���o�z�5���{;gW�;�+okz��X� Yf�Ƴ�ğ���x��_��_���ʝ��g����5)���`B�,;��؁,�YMG
v]VɈ4	D
��iН� )ә+��`������p�,�/>o�C��y)V�tTl'�Dko&�P-fY���	p���T�R6���V9����TA�#3Kj��-52���&f
�ui���r9���en#�PK�7��(�8�@j�W&?
����}�"��i0�އ`���u��.(���Iz�YJq%.��M1��zl��$�zq�]��N"1uG�;��A:�vaIV�$�mkt|���!G�	؅/�j���i��'������@[#���&�i��j�vJ�j55���}[�� G��m��ܬ�h��"��ܩR�d�)�)P\�l��,��7XL1�t"8_@�,��HH:fN_�d��,�HY��	�o���Ĳl�JJ�FN�F���-�)� ���;m B��rt�0��+��2��b8d��)������3�DR�Hl��4�nKU�sJ@6�d�ɺ�^ʣ�)����ܴ�ax��	�J@�moY|��oT~�6-2$���㧟���Yg��#|��A�_	2��c �ᘉϜ�B�7^Rpqh!�9��.��g1�x��x�_����ػ��윟�<�������w��`�G���f��������{�����3��y�:?9�f�����ў�̲�7�n�����9�|~z��<��2}p���e/�oo���˺�����i;7�e��n���x���z�s����/��.�o(��_n���\���Ӗ�G>\z���$nw�'���c���f��6�����ŹЯзu?��J.���ڑ��z����o�?6�s�_e�x���G��xb�!�6�a�R��-˵Y�ܮ��$~���`�lL��<�S0X��p����&BG	��M6�RⲪB��!d�!̓�d�״��Z�L!MI�M
$"��Ħj��xlfPXyj��m�Q��Q����o٨y卄)V�V�t�21�1��j!��R�p,g�m\!$�lS-�������L� l#|�h��4R�}�ݨ�J�.����ůĖ�,��m�,P
-pZ[-�a�Rp^J��%��#0`�kg_b�b�)F�<~ݧ(���h�v�oB]��D���T�#.�\>Y��&�j�J���
)Dn<���L��64�!��
,��da���u��_���4̪�ĒYF�-�"x4Y8B'9U�S%@F��ǌ�,˲RK)�e�	�n_�)�ׅ!���Sk)f��{�*�,/�G�6�8~���}�൬P���e���yY6WJL��off>���DcR&l$�T%�)׷��%`1�u�Q`��Li��$P�y.r��b"@�4k�C��q�WhY!23�AL�RL�FR�đb�$<�	�RSY ���j	��N,%���� ���|�Z�8��t���J�i��D
�[lȥ�Ձ�+��o`~jj�Cb&TH��G����y��D�@�e��B4gRu�e⌲������N^�9��Ɋ�j�fL�l�@>�]��UեR@(�ϖ#x� B�pv(DNS6fj)o3�Y2AR|
�-�ꎖl3��JMPI�|�fP[�FK�W�	ç3�r!�d7^��[2�3���YJE Ju�v�؅ɛ
�I��XP̏r����r 4���@�-�J����2)4�v]S^
��񵨩y��L�Ti���UJ�'(�jw��t52´ F�ǁ�P�yx�Ȧ�P�b%'�34��A��0&P�0i��,�����T�K���� �*>0�8�n$3��r>�Ul�g,�ٶ A�'��%B���D�8~R���T���:2&e�A,���o�e!��7���#�kz)�k���K�f�-���;ۼl�� �9�F�h'��Tb{���l�)(kN)�F���L�~����6ɀ�
1q�AA�� &������^��}!0�r��7���瞗�s�>���뻛�k/*x�q'��jy�G�/wn/�o�y�лe�n��|����?��'~u�#9><��{�?�8������_��;F���e�H�Ɠ�k9��ؼi��t!��xK)��|g�/�aۣeJ�����R��u�@���&+54 N��)����_��mg�H��@�35)4�0D9ĭ��3Q��{���o�R��_����*,5�v�_��l7�v@���:F���������yˀy�h��Q�u<�rMy���ȋ�t��e��CD�M8e �n���J(�E��Y �0ܞ!~
�-��6��A���������JВI��$)���5L�Xʩ�BY/�!x��W���4�W�qi��y/����s������7�~�-���!�ϟ�����?��??y���,O�~��f��\�K�.����FW˛�˓�Ѳ������Po�c#�u;�76q�B�d�ڠ.�j@�AI:���D����7�[�=ir3��1�Zd%��!k^�[�#��l��G?H�i�R���ee�ڒ��Al&�huU�&U��ى�-�뵝��%.��ng��H��K!�)TXI��_�@L:3@|�8�����t�@)���^�e��)��T�iH!�;�
uw2��>���xn�e�<�R������p��P�3F{�>�P@��b�@�a�	�۲^�<<dU]�SbT���To�b���t�;�'�D_c !�A����(�����8�MU`�D�@�e1uIm΍V��)'�ijN��8e�N��*��K�@����Q �!� N�.��Ǚ��2��4eL� niw|�e�!�h�����<ZU�S#ݻ[ҧ�J
�\@��;M�lM^�>��IKYv,mS\�%�#N1��R���!��kS��eU�׷Xf�L�$
�%Y�xŖy�+gʁ��"����o)��T��K�Z��#�0!��m���/�z�B�T:n!�Gk�3pR��W�xPH)t5CL�9���p�)�"�P&RG ���X&��J"��\������g��#_������;?[t�9~����Os�?<x���������|���o\9��>��:9�v�op�u�{WG>�yxsz�w��6�m��w|)wW�Q_��u�N[`���tP���oY��+�&uw��K~����G�Ӯvvݟ7{W�����R��=k3=�Kp}۲��z'v�ȉz���z��~�oN�o�����wjw��Ы�ۋ��뻋[۾]~��S��#~����G��eN�o����NX�vfj�̿��~��z�n'-��-]S�d���Xz��)C㫭E:*ap~��xHx�	db�/Xv�^2Y���;�B%�R�8�R��i*D��W�>�	p�#�)�0�)��Z�EG@?�e�D�j�p�h<k����<�F���𶠪.���c3����5˩�Y�Z�)�,>�ƳD�6�l�hFm���=S�bp��@*2_�l�q�����9�� �SЯ��"����˖���:    IDAT�皿�o�!~����%�`J��k�iB^�rpA`�:AU�|̖��i6!φ &�J�wE�h��� 5�-���l�h@�ED�w�B�H�l4A����� ���lAIWV	N�L�N��1y�l&���הC��j9���Ke�)�H��J�B���TbH]���9���ײI���-@Č,|
[T�� �j�H��Cx%�@R�tJͦ�7��څ ���L�-T^Y�mBH�����������L�V��x+w�Zl,鰡5-³tp*�,6��5��+��
�MUlI-B�xK�-� 3�>`�4)X�� ��#~4�fH����& e�T�gc��Ȏ�	�]��)�wV�bcPed���H	J5�x���,�E��!��f;��<!T�?�L�ĝ�r��0�|�kG!C�HP0K�1U��q�����@��Rs�@�N������{o�<>2�eUo�����x"��iJ�M"3P��Xǂ���.	R�D{��\߹hq�Y(D6Ӯ�T�z�ل5-;�]�ݞ��eegN�S���Um?N�[�d�Dxq�^.����J�l���g��<	Z�Yv�DԮ� 6�c)�7瀪���{��T�j_v��ש�z�_�QPEm��K&�P�Bs�T͝ ������d����(L��B���eɇ�X�#�|���)�9�YH�8�b��xU�8Iav8�m�i��o��̶�rK��)#Է�I���e�h<6ҧi�8��������fߧ4ݐ�������_�����.�}�������}|����o��'����r����`�v�Oc�D�;V|C6v���3xLYc�"��"0'���T;I]T����wK�.^��@���Ջ��g����gh>��c"^��-�Ow���C���_//���7>˺�
�\�����b����y����/��'�=4��`�y�Go<����������w���G�;����C�؅�/&���aⲂe���l"Um� Hmg!��L�e
�Z6)��K�<g.`�ZS�15K�&M燯c)��qꢝx���Ҩ�#����|^�q��r@���kMS��l��u��{@1:w�5)�f�@�k�&[�̽���[���|�_7Y��r�.گ���hz�5a�y�T�l8���TA8>�<��׈gt��8�B�]+���}fh����Cm[<B-0��Z+2A ��FPଚ�8A[�d^��aM��eZ����w���yi�w4~��_��_�N��ȕ:���s	���<�����u�l��J��{U7�7>���n���8_ܽ8�?��r	z�q����o�
G�����aJ��lYZL�Bx)U��
_Onyڴ$����QI�s�;�'�#2B�9iB�!.��s3��W�)���b�P5�]���ẍ@�� ���4pU�<rӫj�Ų����(�9�}ʵ���
��hv^4-��������J�W+A�bT�r4��DY��I9�.$ߙ��)�zґŧ�;pcI;�Dh�!j) d�����Rf ���������h��MjRԀmG�K3�T�<�!����,�~^�z_VЉ�ez�� S���&���GT�c����!�(�+�V9��d�T
�Ց5���5j��k��5����Ł�V�Q;����vj�(�d������4��&ˀ)�i<ʶ`�8y���3L%��*��K��T��[*����*K�b:l�iڡEv�tWՙ��,��O�A	0�-Y�(@:�eo��U|���K)�GH�iF�A
��ݙ�R��J�)W��F���&���t�lS�^8,e"��u��W�N�B�@�Z"41����FO��}���+�����#�B��LJG��"�:�6�L(`�C�є�u�,�ܨy)�Rd&Q�jr�U������9��;~7����ó����ۛ����G�=<|����#�<�ݽ��o./�	l�=�%���w�����G�7����qo��+B�������e
�2�𝕠
��L˺@3# K�:1	�]��ʗ��]ϣ�ѱ��p�g[6G��Ý�͙���{�>:>8�/�wI��1>	��z�u�FsP�2{Ǿ����o|'gF������Ǿ�::�=���`F2дf��A,�x1&P֍�Ir����g�0��u#��<��R�H���8}�Yct\<&AA1߲^�H	dG_�2����ښ�V<���D�1;i�e��W-C*g�7ΐ�ˁw���(@���Բ��p�0}˥�j�^i�3͘�����D���[b��J�l`�](�������l�`)�7�@!�}�����9[��Hj�n+�"�&��,_#�h!-Ū�:b�����n�J q�T�EP	��F�Z:ɲ��R���	(��c� ~��%�L��! uq�-qXU3��<:�0N픠Y�ˋ��-��O����jũU�	��[
DC:�@>�"��`J�i�N����� 
����舕�a�O�R@��Z�GN�9Y���,�y ���-�;vHGT-\��L-�^���B�|�GcV�tZ�UeY,;cOG3�4� 3��S9pteU��$oY/��RM�ݴ8���<��Ҭ�!y�8�ĩ��vL�/s�z��+q�㧼�]��d�KVo��5\-��u�M�]W�ǳ�n��ݲ$��,ٖ%��x�	���o�&�/�;xC��%YV0�l�/uϬ���w-%�Y��Z�Y�z��{�<Uy��*Y���p������R�6f ����L��
6���ի��iN�WƊ���J[A�M0BL��ȇ���~IqJ/�PE�,��ĜUOKm�~i��%��Ȕ2��A��9�d1s���zMY[ġ��=�P?�j��(:⥘��%I�Ŗ���ԭ�JN]��Df�}>M%�g������h�(�C�,�0�J ���E�����s�9r��~�=�!��U)��ESÁ<C++�D"T�(_:�§3?�P%�C�5I'?��|�?�U7rѺE(�PV�J��(�/*T�ۆ�V�7v��_4����� �,B��Cv��3ƙ�L�3�1Ւi���f�p	�AIw�Nx��*F�rF�VaԌ�{�A�z(Z��e�o�j��dU���I1E�dM+���Me+8�ҍ5���_���>�d�We���,�j�fj�ea8t�Q.ߘ��n��:e#s�Es:1!���~�y�^y
}��%���gu����L���ң#����p�_mѸ�2��|yqq�:������~��?�o��Yq2Z�X~Nدl��x����N�9����R�Y�=sp����!�X�o+�Ȕ��)%��$|�����	�/��ѻ{?�L�F)dz��p�^ѣ������ﾸ~�r{��wo��ޥ��γ~|�5���g��6Ah�R]E�A Z{+��n�!��t�(���M�p��N.2��#J�� �t�\H����6" ��yE����*S�ϒ5�T_j��¡�e�PK9ӏ)LQ%����ò->�(S���v���ѿ�s�N-Ofz��h+�� )�t�̕��6���P�S��%'�`R ~]�>�+����z���T	�2�Ɣ&զ�!���ߪ�m��ed1K�X`#&d_ц��H�̏� �UGC���
a⧜Ԩ����E�֤y�����y���pTW�g����5�yo���~��?�������{�Gݟ~���|�'��9�N����L���k�ý�B9q:�kSۚq�($�F�����O
���չ,"R�|R��<��C�0���#�cl� �(!�t[�=�t�
���\�a�����=Y�*�U�P�2[���-��(-���
��T�4�u`[�w��ؚS.PhK��m+Յ�KA�ՅG��,dʩ蒶��6�զ��"KāP�u�.�V�!0����̯�D�
��e$��m&�/E�+[��t4)�}G"��a��R R3�N�B�ZE:��!e�K^c�hjI'pgD�j���&��q:PmhXV=w�t��U�*J�Jִ�FS�(Q�p���J������4SֶH�OzR����FPEc"`vp�!S����i��m�p!464�����w���c�F� 2É�ђ�9D
Y�RigBΥ�i�L3�������)\.����\��$�o
g���>MY�V.�z���S �)��%�r]��U�S?�e��ǔ�E(�r�DuE"R�]�s�8�L4)� ��ɑ��df��%�C(ԃ}V���C~*�VG_b���)H��2���E�r8!�
M-�
a��h��Ь7�+M��d�p:@�.��pD��� ?�kb���yusx��O><{y{st��� .�
�O_�Nx��#����O���������pu�w��yL�r�:<}�h�ڼ������oQ�w?`�-���_��m��M[)Do��//��7���h�k_bk���8�_x�R:<�>����C�������6�/W�+�������/S���8:{��;�qo�_�m<�0���?��_�b��>�������U�s��?O�󇾿up�t��S'�����ۚi��P֥ۘU8&��c���W_�;�v�!:d �H��]��V�2����0ő�"�I\K���EM9]�����uH?2�VM�V:rj)q �!Yp`�i�F
�-M�=l3kc9u2�Ԁ#�?)���lڊBZ�,`xӢ��qGYV��˺���I�ф�D.��(�@F�-��ÄWN�oǄlȬB�h�d�4%�Rch4�p��4L�Jq�cU����ME1�S�E����2e��0�S�rS�Ҳ"�����XL�E}oo��� �,=�_!�Ս|�6�b���E1��Ѹ��{�7��G6�h�_-��z]�����Ad����i�TO^(\:5Lx�Ư�Rlg����6��9K��ș5��&G#ƁwX�.����$�?0��i�pK�/-Ŕ��lo�9p��%��m���D� ������$�}�T
��_:�1�tB��ގ��D�1�!0N�,Խ�|�Fki�5?��� DN��zK��p�Dp��R���S@��BU��w��N-�TG.|�§+���d	epS��h9�l_����R�ˍP����9}~�I$�ωl�o1�D�h�`�� mH��D���k:��IG�+��O3��s�"0>D'�������,�N8��)��(1~%"Ԁ����%��X�DR+ň��Y[g|d�Ԉ� �#�2H4��a{YI���#KM�X:Mʦ��L�R����K��XS�*�D3��LY�h
g�%�/G�R��Bf@�42#|Rd-�;�/��5ɀ(�� �]��8�h�@>���4��wl'g���%@��Tb�85!N'kY.r����A�J�	DcVía�K�����+�h��ֈC*���/Q
O��ɻ��m����������F��ʭ��@
���	oa�����)B�)ZE!D�(RW�#���hR�0`ݚ
uj��)s��we_1��p�����i
�b���h�C�Aڬ+����n�*�rX��)�8��]}��1K��z�B�����`urp�V�\�k����ۓ�������/T�v�Zn�/�_�\�u���ڷ�|���!h�Űt������h��޻�9�=-����<nj&����?^w��GIht:hxdY��F�����&�yP#���O��X��ˏ�u%I�gN�L=h�*��f�gQ���f�2��B�B�G��U�o��o}:�2R�'�g�}���
��F=(M!ߨU�	1�DC�od�K3�_���g�R�H�[f/��'��1��T����\��r8�tD9M����/T?�5�ݴe��f7J�gݟE���YHqd>������?���H��tH1Y����@��V���˲W~�*��#�o�Z8�sj��ѕft������cB�) {�Dև�U��o����T7BJ�
��ġ Z���#��1�����I<<f��R�hJ�š�o�Aj�O�I��پ�`���@!�Z�|��ql�/a?�����p���?����|��R����{W�Gv>�sȮ+��Ө�*�.d"|!�C$"*��W�`l����w�����(�9��g��pdQ�o�҉Q�%�r�T�M0�Gìm��������S4N:.H_j��'�A���F�Y��ˇ��!$�o�R7�[�P������gr�1q�FRz�(��r��b2)l����e	��#���:�_9d_�:�7��4'��,!�]���]^�����2Y�e��:Fc�����&����_?F����5� �@R�b�v��ᠺ�Y#Y�d[�Ѵ�Ev�;�C�ĭW�uE�c�DS-��rb��:��>�E����ՙ�U��Y>��hF'����WN�>��pX�B�������h,e�q�D���Oc� I�]��=#�W{��֒�jL�b�[����d)ͩV= kYQ���^}%�<<}%�&~FJ(ݏ�j!
p���M>��	4��z:dw��Dk���LH!P�]9j����ANG���� S����V�HJ	4!�Bi�[HՍ�T:��S���u�O�F�r!#��:� ���M4��-�����4)_�,S��eY��ŕ�kS�,�#��դ�Ϻ��=miS����=�K1R��+#��[5m��u��2|V!�p���oO����\�������7�n�O�|�������x�=������㛣��Ǐ�ݨ����˛՝��z�X�%3G~���nuv�����v�9�:�[Y�׷������ܼzy�?�n��W��m�Q̽��
Yl���4ӮM����:w���C����f�}t�=q|�����ѡ�ևޞ�#;�@���=��2o}#�k�?�|q|pzu��:��W�e�Y/,o��w+�l�z{�]�<ӿ�:�[�w[��v|uh-��v�7=/������b0z�cyw$�ޞ����ʄpL��V*˵�����31�(��v���1
p�)>3e]�1CgZ�Q��K��n0�.oId�Yl��I�n'�9D��R+b�_iR����h��:�Q�L�XB��bSD��d19�_Q���B��ÕhiFֹ���(c`�p�B�SQW���A��%cm��]]��d���)䗅�yY8��,�+]�äDCȑZTvV����»����8rq��m�#��7�
╘}0� *����8��|L&���@H��唘��8Br�N��� ��M�K��@>�X9�K��=�bʲʕ����$�7��g��6RH��K��W��tڱ����RҜ�ڐ.���|x�i���p�V�|����T�_��۟�p���!l��ȅD�;����*�z:����Xj� 2��?�%p����Y|�J��)�+�BC��VM�D��)'�H�A|����ST��҄�1�I�"G�/a�('AӚ�s���aHY1��l�1�3Qƙ�#a2S%
E�gp#D�/%��
�=4�UT�B	�.M�Vaıi@���Ur�~�I�˪�FQM�S�X(�Q�d�-��iR65j,͔�4��g�-�Z�v?A���8RZ8'p����X� 8���N�}ő~����6 5Y�Eh�H��G��%j2�h�pS���ӡl(�9Pbc��L.2d�M-x�8�^V��@�N���5Mٔ�����L���։���8�:��d���p���EK���J�#s��Ym�8|�En��]u-p4��i�����I
�W�rD�о�X�ꦪ�r����09J4� 9��]Z	R����7�Y�t'����O��'�|♃w�p��+�WBue���v�s�h��
���BtR�^�2�#�O�rƖA��)˯��VJ��{/�% ��{kQv���II�b�уi�qLS��HA
�.u�j�÷��hI5��
��=>NU�I�V�(��ez<z��2���zs���������x{�|��甏���g��7��no.���������{su���v�~�����Ɵ�;=����c�KW~	�݁�uU]V�f[�����Va���e��>�����2ܷ̊h��iM'�l���G��O�����MOo8�F���ޡ�!��0:�6Ӆ�٦��g>��GDُ    IDAT����)T�Swي�cv����=;YE���h-�F
j��p��^A�hE�vfh4�,N"��Z	
Eȑ2N��J��_�^)%"d�k*4V��)��t���T>�Ӂ�R�� ɩ�q����^8�C8���GP����}��S!4�Э��]Wᶂyx�!m���!�L����_
���:�sͺ5Jt����u�t]�x z��:��|���)&ӃZ���6ESoK�;�����������r�
��]����s�e�2���1�'�op����Fvڃ㷐8�]fq�'�T��P��~���I�(ב����y��?�ܕ�t0}P��M0C��o����ޜZO�!�E�w'�$A��C�C�ZB9�p|�s��}���N�KbL8}'�at�,��b9]�m��X����4�@E��M�����w��V�8_'|�tL���H�vW��"�4LH�_�����ύ��T/���%Д�1��k4iS�iNc=)ܪlnMK���($��)�Y�t��5�B��9�F���8p�۲�=~�E�Z,�S�|�7+�,����BT1�ү=c�9�)��\�΢�C�G�95d`[at���ի��^3�UQ|U���E�կC`E咥C��F�+����f��А�c�`rԅ̦��3v��d��4Y����(d�ihL	��D��.�+d��-
��e$RJD�)q$�2�tl/�,G�JX��y�:A�F���K�i�Дn��D|�i&K��l�6_���^Q�LHux+E�C��N���;wc�qtb�L:�,Q'�W��Bhr�.���ClB�RD�g� |V������OV�����v�������@�+M]�Z��F�pth��=��DfhL�D��/�Vo� �G6m��eY`�@h�!L��9�@Ӥ��@f[p� �Pc퍾\]��9^AF�����wi2���z�v��=�����g5@��`K�p�R���))��p�L�u�e� Ǭg+J�������=<9�^�~��\�|���w����o�ȿ��^o�o�>߮�g������͛�c?�y����^n/��~���jy��������������N�f�#GwgՔ���zs��|O�b���V����&��A�u��ۻ��O�ػ;���[��GW۫���{���ַ�?��|ux��ɕ)}��'�]l��=xͿ��\�3�L����g�~a������{����f}}��s?q)՟�����<_nD�W��D��:��W�}��6߹�vA�ˏv��N(�������� �����X5&�xQ��m}!%�VCj�n��X�r�Ԥ�M�P:�b�A2�U �w�e	����9�)�$�����)qD�+a��ed��?)��jCv������X<eY!����A���)Teҗ��j�o���[��Vp�|��t$������UWW�FL`4c�4�O:��
�f$�C;	�UX���,f�#��I�A.���L�8����C.�P�BU	I^�����
ݥ�b��i�+�����+KTJ{[�hj��ւ\u�M[��0���0�|��L��z���@r�`�T�z�)є/Z���n�/����$�课�(�HP4fu��R C@��R���Oo%�O�J�)w���������-r|R)çD;D%�uBdA�E9�E�U�i�āsy�㳖�?S�����|?�'�)�VˍV��ݵ,�pY�����"!�5bVg�/�H�#�1��(k�n�����!?�G���G��*2��S��4"$kLph�z�ԡ]r�|&4�
�r"��4�I����ei�A(���L��hr����zk�πF�#�)|�9�1��P̮v�dᜐ��о&���k�ȧ�a��(������[~S���6Y4�E9�F3v�c���'Aj����o��.��7J��T:���4����lm��+o/+L&D?�� ,���1��IUH��Q�|�8�tдğ=Y:�� ��8��l� �3���M'�h�|��.+�h�"���Rf��?��0ܔYT"��M*~�������@7�8r���v�&Eb�g�Ò�J@�T%ڎ��֎��J�b�O�8�Pf×R�C���*�H��қ�UXQ�jq,S����)�_�d
�C%��%!��-��'���+L�w��E��9����H1e�B�� g�Ǒ���M�����6��{U!~R�� ���C,��juVY��;�� ���s��r�DR|:u�g�ĩ�Uq{�99\�/���G��jsw�¿�8]ݞ����_d��>��<��(�,����_K::8]~Ӭ��Ͽ<����S���+�����py��M��-���r�̺�`;��i�v^���n-!���S��+�����7
���S;�I�ry'$� �j��=�BV�S��E�պ�X9>��{n�|��\�R�r�aj���\-���I����SY��:���V�W:�tF�f�0~!�Yͤ�ß�| U �t�rLۍ� �YY���.���!D p�Y�)K*B��+>B�1��m,�D�cWm�s���O4}b�w^Bh��'���YSc�N���}�SM���5�h�;;�	��mѳ�2�k�����T�ԒO��f|���cN�ׅL�+�G�.�>F���tq��t1(*�>ĒMg�9�?�4�>�O�~Y�H!�,�h�օ_�)��Ö(+���Z|Q���h�[�bѦ�J��\S�fڊ���qHt.�/��/��Ǚ?���*�����9gT����b�q�9�J�ta@r�ƚ��������L*���i8���(�%G��qt��/��mY�e��_�,}B8�hU�X%�B�rdY��t$�Z�'��J�-�d�?�?�Q]����P�5W1�ȢSԋM����uf��.'*����X� �KM�R�Ŝ�r��b] Ȭ�1հ1;GTA"<QN��M�پ��$��_��P��B`*�G���*:B#A�5�O�srh=}�tM����Z�ViQQ���E��N{@7Ϳ�˿�F�-u9�����\�ܣG��+�`���X�4Ɯ�W�����EkϏ����Ŵ�.$���h���ɂ�i�>m%����O?�TK��b�*��^��==��ˤ�)�u���1�R-1?�$�_!8D?zp��/38d�|�
čbu�B�HAK��S�д���4K����2D�2�ǱKZ�~�����ہ6S'�L�u�sd��r!^��Y���H���b~ Dԗ1{��_�JiSms�'bEh?�я(;�ƨ[�����$bJl�zƴ�R��t�u:�_�t��5��mc�F%�Ȏ1|�uI�HPԨK�Lj�L!��M��	r�$��rF����>�R-)�(D�;��2q��s#Y�L{��L�a�Ju[>��ڨ~�ZE�2���#�Fj�����4�)�#�,%���%��X���b5LMn��^i�BU�b�s)���t)Fߩ;)ת��>a���"��.������|��������}��q1_]�<Y�^�����_��psr��K����9;�9������ŋ��ksc�����|���G�T���w�����bsp��������o>�D�rm��9�ԘUX`W�6�h+�Ț.�s���A��m��no��V'Wǯ�=�굷}���˛��ۃ�������g�ך�9��Ur�:��z�����+Nt�ڷ������Ώ����7zq�P�~���v�3Q����������M��]����w::�jMZ�� X8�W��1�t�������	��t�|H:9p��t��z�,�o�����3�Z����V�)ZS
��3`�z�A��2BF*P�5 ��P.�|QMÍ��E%8��n�#�+!�d���
�+e:�$�����Ma��t�D��*6v���8JH�d�Sغ��k�ęr 5/}8��D9�7E2 Kߴ~ʝQ{�~
}VΈ�HD-���N9�*��B�|#)˧����"S@��f��b��8�K���K�푪b�`vJ(K��zck��(T����>�k?qL�}_">���/}dK�O��H���g!@⦪0N��}���hEKT�;�.����j�U��JD 2S����h>�4���2��?�DH�ZF $��rB�����v�J�Y�^|�%��+*wڐR	#�*r�P9%�0S~�Á���"�>뇣��DL�"�VH(�(�%;cNE�B&=ܘ#4}Ҝ�җ���.���59����'��P�,��B����R:���E��������?���wFJ@L���Y%�̔A�1M[��9�#$[�@~R���(�84#�
�w)T���h-VnH2N:%b��>�D�F�a��/WKn:pS�)f"SV
�>>`�ƶ���.�tlZ�_�p8*F�o^H	�ZR��1d
��'�)��hBFSV�@�ow�-�1���4�9#�&#$�2|�����h��Vn�t"}�O"�7���	D3�'�_�U�MF�[QN��:�^}��H| �:�*� �6�@�JsD��ū�"ر	�,BY!�+׹��L�S�|��G��k^(5�9Ü�@f����_����S�`�m������Z{��bßtM!#>靠�{�㡐g;.]VKhR�6�_�DHUη:3�U��F�z@�#�M:P�*f�D�g�a��D�@�پ�`�DK���V�BSx;���j��O*�k�,���C)$���N_����S&%��7P�#dd�߮�G�co��7�w>�|�oɸ�lo�67���#?�_p�9g�����_����|�>�l�nw�C>X��-��z{y��ϟ>y��[o,�a�������' ޏ���J��05�[��}`�Q�L�	��#�f-��6�v%Y�HM���(����S�=�؊�'$Ȟ��zW.�i���������t���n%Le����=�R�l�)f�THKFo�IY�gA.Z
~9-�DQ|jt -������$"`C8�U�\�8���(�)�,���FYM�c9|�1�L	���,#�����I1�ce��K7�X9�Ԃ�ı�FOW<�uk��QjOä���<
���߁q
N��?��9����Ѥ�7�� 9ҵgg(�����]T6Nǅ'j*��B�V.2�CZO�="f����`kҳesZ��Sc���B.mۊ��0]�r�8�j&D(P�1L�1�(� � Z�\�Q�\�,jс�����Qh�>�*Fg���)kZ�\酌�	�7:-
n=m��������8)�\?�%Rӡ�J�(�P�єl���"�=D(���85G�'B]�)�R�hjtQ�ϸ8��cz���QE�l-!sL�**�YH
�R��Q6N��*J�����[�A&�X���v�e��J�ӕiO%7�S�T�
�&�V�45�@��'wz"�S���׍�(\:K�5ۣi��ˁ0|RkQ.k����r�>�\d�Z���:]c�+�-r�. ��̸G�\�n(@!��/5�P�'�qI�ES�M�f�C�&�FYVO�kF�*���#�d>�K�0|��t�:Bf!mBuUј�*�	ז�)�oC
i��~�iM��@/Hk�Կr�V�V�K��J��*z1�N�gi��4�FJ��>ת���|�P�·�E���E��;��*$�e�J�k�O���&nj	�(A���G��6�}�si�|��O�C�� J7�(
��Ǻ�Ǣ,A?8dmM���מ{y��9�EM��Q�
:徳��E�T�/K��uѴF&j+��R���Ǿ������O7��������7�4u(���UTi���TWǧ#t|��>��o��9�����w��&�WdѨ���*�,�2�e�N��i���O�*a�;e[jj	]3�Y{���eC4���RK��ѵ-�yA�kIch�����N��Qo��L�)#ܗ%��{bj�J��n��Ƿv%�;/L��V�r�W�r0-�y�u��ŶuĽ�zeuQ٫�k�5m0"��7Z2#kJS'髈�5YuN���wv��u
�Z�z@`-A��o������_'{��|�ų�]��������o>^o�>����`���������͙w=WG�����`�ެ�=9����������G��f{|��������/��CF��ֵ>:��i�-D�z �P�[m�{�U#j�D!:�,�M�0?w��Es�^.3p~������˛�o�����Go����7�����v�gR�s{��>����ϟy{�~p�/s�'���������ӻ�.#-y���������SE��Ѹ�5�unE�鴊��8���l+���/JJ�RM4gԅ-d�f0E�5�ikL��D>�1�OS!YF:U�p���`L3>$���G�O_Keዲ���1��s���[����fu�M�EHٔ��*d̏��a9����ݯQ�4[B!�C�OoMQm�N��ҟ��j�T���&�i��t�O֏,�v�!)W;D���hY�����d8t��k��LL`
��VT������$��L5���aV�ܾ)����,�>[�X��DH��8���O����9>&��B�Z9��"�#Ĝr�-����+dԉD�,H�oD0J	��o�ANd���SQ~�*:\/��E��QKWӀh~wQG���)75d�|�hE��rBEMK�tU+A�iQ��4��Z	��0�_+�6p҇C�����2^}i Zr!+~#)�BL�C�ʙ�MYN�9Fcm'[{����.����h�ȩ�BA�fQ�1M�E�u��i	�GH3NSQ�X��@28���'~OY>F�p��43]M|'��Z�Be�[B�� 5-ע���z���8&��Ƒ�P]�IarT1��J���:e���?2�\��)��i���)�D�h��xj�CT��R�H�O �!K�[iј)c�6r\�"q/,�HsZBB&^{��B&1DKY]I��q*Q���!��w�B������D�Q�����$Z��Ʈ�B֛8����m:���P��lV�Ԉ�8gJC����?�8%
q��©��
NR|�����KO0��K�������YQ�b���'&�,�\�:7�\L1�Rh!B)�T��0�D�7��HI�o����r%⏈(�˂�2YN��]��+��O�����ԥ#�i����6���\��z�M�e B�S�%��}DJ}�є۟�N8����d�r &�hH~8$f���e�+��I)e�r�	G0�F`R�h�H�K��h�I
�Á��o(�6�b�>�<=��b����c�{x��g�~D�h{�VW��������w�׷��c?�,�O��Q�e��V��������f{�|u��c�_;{����o~���n�R�������Ó��W�#+қ�HcmK��9t!��Z]`67�c2�)fw�.!���s��ZUȃ�ҍ.3y�r{��Y
G���q:����B�=����	�Qz���8|���"{��m�gY�<��jO���r*�ؒsT�7#>0ܨ\K�S�j�!*$�o*�q�2Sj��g� SH6B�|�h|E;_�d�85S�#�T�+i$�K���t�uL�yB�o��o���m����6
���|��O&�F'��<T1�������5Zud��@�n{��q�6����n��oN�8�)KT�?"���ٺe��x����-��L��v��%zP�.�v���ƶ�ӆ�oBh�o�ںR4f�L��	���J�%@F7∖�_E�14���%4�����TV/�)�F�R��)�E#UI�Ȩ�OO�]�����=v���킈,%���R� һ���NR<���]]�奄kC.}�=��OM�����r.?U�1\9�D�RT�7%a��g:ԕ)Gb�/iQ�Ȕ�̌�����&M�d�2��x���W��/̼f�L�^���5'�c�	Q��V���)q�]L�Y���L9B�d���Z��A�̋Y3q����t�ЉV��V����a��)���?M����Jg����+��@v�g3�AD��Y�JԤQi���X�~�UrX]5�4r)FYuΡ��Rrc�r|�t'�:Q��	%��f�G��xh8�,���A�%��u�����Rť_-�J�yH
hYƇ�	r�X����H�B�0�{�����K���F��c��^-dRtT7�0k1"��2}�`�^�����5���T�K�:e�Qm,    IDAT#�&��Z_ �B^�vF.�D������_'��Eo�唟>}j�|��D��D&K:�D�̖"8#=���C�-B���m�6�ͽ��{����i�Ҁ,���t%��֛%�(�!7_!!�Rr�6n��:D�)YU�!\-ˡ��U'zӧ(Z�a��#���-���Y���)Ñe!���i�C��l�����?��_*�+[�6��%��L9D,�J��O�H�e*�>��,�1��/�K���F���/�������\�	�]BP�J��};�U�Rpr��G�˲K�M��-�����±:R|4S)��n��7�6V�������α3��8yy���������//������㳓��gnɇ�̦�A�g��Ճ�ӓ���Nܲ���}pq�]������o�ɷ��䫋�Ս/����=ֶ_Q{}����5����}���o,4�4�IB��X�KNhGyuo��"#�"�=�'?���k��]^ܬ7����N������W�����g�'�~�����O�����Ng������v{ywx���O��O�}�S���~���?H}y#��u/^�=zl
���Z��ueW�=g|4Q�VM�s��s�8qѤ��7��ܪ��Ο%crpL/S��E�)�����NHt���(�*
�b��@#D�1'0�L��P&�#�,jz���h�������8�R�"�
�EM�~z�h�B��jM]
�@D�s�~JO�nԏ��PMNV�R�DeS��}Չ���h�F��h�M�*��o�O<)cYi� 2�U:Ajp|�jI6eY9�R.Ǫ�S�C�l�4�ۦp��7�i����H��VQ"dQ�!��v8�E����r+=�h��DY5��Q� ��G�L��#O�(_�J-�}�p=�!h5�T ���z� A�BάZs:�t�pd��X���hV�ޅ�n���n4�?�T��J��?|��� ������D3�װiYE�j�oD��NuK���/�<�rM�J7����Y)��oɉ��.L�,�8�1]�zHS�է48�fc�o�B��U�s=�J�H�1g�J�*��" ӯ%�x�)���e�9)Y���#)�Hj�1�p�
��d���Z�".�)�/7���*%��#5
�v^��Y�y�Tژ�-���)�u?)u}���9N4~:��J������s�����,*�4�`���IYԔ�n�	���3�,S`GRE�VU�(����B@���)@�t�ʘ&g����6�߿���_=�d�T��B��&1�#�P"\W��1�fO�ߴ�k24�ߏ��Ʃ.��M+-2�*Ŵt�Y)�D*(��P�9JH�38���)��M��>(:��BN�A�y!UL�9%&X�| ���B��|SR����$�_H
B,��4PK�Me������j�ɑ�#
����_�ڮ+����T-��2M�qB;���Iy�x��g�=��K$[�hl�!j�8BL�F�q����J��bp4+ɇk�h[� )����!U)DД���Z
7�L{�ȪW�od�t�L���Cd4�!;��M���nJ4c�kl�@l�������T�������^Qf}��������~��x��&�������ǰ�'��?��pm�����[o�)��y�-G���ѩ��?�����:~�{�����~���g���7�1�' ���~v�����5�<�*X)�S��r�Nb+v� (�+`|#�)�g#�)s��O��q��En{�+�!�Д�HP�;z��<��s!j�,�Q�m�nQYay ����/y XuY�4�Y� �U���ꪋ�� !M)�F��hɢ	�!C?pj+���SB�A��:����U��iN��t�FD�B���*>�q�'x|����>��Bd�x��#�#�g$@F��4��Q�K�%��j��Q�A)�U4�f�F6j�y�����'�RЈS�KS:)�����z�+�s=�l.�1�|��ǘ&�	�g�.�=S"K0)uU�����Q]9'�(T��E�<?��s��
f�F�O�tNH|")�jD3���{����5�0S��Ԧʤ�����Ji)^�FY�)�����O���jc!�Q
�ѕ��C����o��&JY!����OSȔ��UH���@�s׃Cw��Ѕ*�UhXK*րܖ�r�HR��/��Z�#P	"����ߞ�.���i-.��>����-�KuMׇ�u�#-�T��fHe��@#�('~�5�g�M�SE!��q�S��!��6Y�!%�{��a���O�O
�3U�	.��]V��1ux��x�u5 D&������������!WLK�c\��ol!#�l�e��s�C0u�"��%2���	�Pkr�h�2;��,�h���#�ۊ�^�D�׎ �4���zY6�+�=�g?�N}v"p��X��@�mo�I�§�L_��45�V���W����S�����p�Q45>���c�}֮�BL�$��K$C��0��#�i��._��t���(Y#5:�8)��qL��yux�k���� ����*v����&�m����i۹(�WBi���T������eѴ�Q�5Z�W�D"u��r�1)Q�Z��Kw����j pg��l6
�&����S�y�%��hC���ً��\�B 4��8D?�8�Q��r��S])t���1IT��rj��EHD�(��;��6D9����ڽ���_�B�)}׀�f��P�����D�+�k�ӧO�Mf�jR�����Nom}ʭ(�k�������sgO^?=x��w���� yvxz�������?~���?��g>xtrt�`�/�����k����yx�~�'�|�v�;����ͷ����y[-_�5����5�;��fiK��{؞�{ՙr�ߘi���� �,��+�xosuyu|��[mN=~�'?��[_y����ѧ���g��jܻ�����j�]y#w�O�lV����~������?z�ɣ�������_�s�=�;�E�w���Ǣ���׸:וf|G`�n[n���%a]~��(��:8����Ǌ2L�(e����Fx;�z�؍L�J�N D"M>~9Y	4fF02���	��H#�R�)�)�J�sX��!��ő(ķ	ӉM�a�) TK."y��k.Uw=tVKh����r�i
��1��J)�T�*q����hʢ�J�X�1r�u[�H��Q��� F�F��G㏙�Υ����4�"�a)p��B�^?�j��F�VW:�S���duK���MT
K*�9��:A�.��K]:4�"Z馽*I!�ǁp�S�s��qZ���áC�qT�q81g��bd��G�R7�hd��b탧G�t����g�K��y値J1Bl� ��3Ȭ��M�4��/�Y|HQ�)���G6��)�A揎h8��Y�F6�bd��2�K��R_9�D�
Aˉ�ů[�EQ=�6�D�M1�z���Á��R%ͦ����ȲDk���>��GG�#��8������l����� �)�2ME�Gc�Ȍ_t�
$�Y���vG�U(����3���?:B��hKO;����?��YBYm#�i�S4!j�$��L*p�tYdѐMK�m�{T����#�1fi)����,�F�>��6DnR��{�B�*��7��W�=}�J+�)wpS�bJ� �d;}�Z���($.*w|�)T�8||�V�3!La9q�J�Bgͩ+��K/1~K�t��4�� 	�p�8��]2��a��?mx��98�D�o��CH�3��X����`�ȵg�R#�����)� O"��C�x5��KOY3�)�u�%����F�ǅ4�H#ޔS���cZn��cS�����)�4S	������:)�X�B� ����!�>�UB��q�%񍵭O47�A锅X��J�I��yos�JٛDui�2��B|�5>eQ����H*Д#�=�������2D��]��)�1���f�f�E}�� }?W�B[�o�s �eE�<ǻu��V�,C�Գ�m�f�M���h����"���m�AS���M����|�y�2_���31��<��-~?�zus}�4�͍OG�V뻕mv��'4��O?d�]o�WI��g�oί��>��޺|����ϯ���>����{o�W�N�mCu���w[�|d�r�9�>4Z��5f�]�@j�@��Ng��p�=Cs���M}o֥eħ�k��w��M)$%A�}������pL��JT���1\z��g/���C8O�E���S���9�Eіu�_���h�Ȍ�\Qp�*7Yp��qtv����5馅b&2%,��	��֊��+Ԕch���):k�w.M�r���s�h�Pд�ҳ:��6߃MOc|@�<����y��h�l�ǡ�u���SV�:�	l4,�[��
y�2�z4'B\ۊ:w�M-Y���<&�O;<��<��C���O>����e���ܯ��Qր��8�XQ>\�@>�+��V$�ZRRf]|���|L;�JmD��%��P:���$�qi�����!)��VA֔�̉f�C�J�"�t�SW���Y��R���"����md�.�օ�I�G�M��Zc���a�к��p��՞~#LU(@v����)���Nd��6��E��L�̆ �Z��x�i�d�JA��Uc�D]Ϟ�����3_O~=�w�S����Ҩ�j-wp���"���|�E8�#X6��P%����1��<NM�F�ŗ�K�i��$hE�8&��~.	���8u�p�;
p�B�����\�^�p-U�"�)�8ڦɯ���B�>vێ g!Ȳ�i����GcE�Jh��$�Z�ҩ�MvF|F�HJJ׆k�&��B����i�i)�r���ȁs�	�Ic&��	�`=i�'���s�6�����J��gD��hC$V�M0u���Kg��u�&d����j�q�rqd���d�������t��BZ҉i�u�� T��!��L�/ٴ�E��L�LQj���L��&����fc������A@6�#�t|�s䊚�������D 8�&v(��B�dB�A�/�tJr�3�Ɲ��/."�A��� �Eг���j��@��i�v��ٿ��0�z�z��J!+���3e�/�5�9�qLEk�����R�PS�sWH��+D��;������;�B|��q|��o���֤#뭱eZ�fl���困��㳇O6W�ӳoyt�]����_�<y���n��Ko������������h���K_NV�g������������������/����cղ���%��D{Y'��
q�'��h��w+�jZ~�h��|1����D�V7q�W�?��?}�ճ�_��^l?��緇g7�cm�>
%�m�����?>����~�o�y�셟:�xyx��j�3,w�W/�9_�T]?�����6.��=��:��s9��# �H�Dh-V���JWHޅ���]���n^}-C��B���'�T�z��P�Ԍe�Ԇi�������)}h��C�3�>-0����N��B������1M"`V1�5"�L��0N%�G ��LP�h4���5����Hq%�C&k8ҁ�%���`��䴊��a����3��B!Ʀ�Rc�X��NB�5��
�ӈV2��Yx�@����@2�=�+���pL�˛�U�� ':^���S��@���qZ�0d�c���餩B�8ɪ^�)t���D�j�t��,��j)�k:�#�^I1eh8�1S֌)k�?�R�H�CaǇ����yS���3���Y���R�B ^w����"����iHc��Q"�J[�prFj�s���'��U}���4�����¸�2��(�N�t��-B�D>m'�h�E���������4��O����k2��N�19���8������CQ�)���$d�D@6e��R��	qb��$�3m4E��8���������6��i����rpX��r�P�t�|��g�U7�:f`L��� �qr�E�!����=j����3�WB��+׹������`�\���"���;�N��Ě�T�]���q_���!�^!:)8�\��4�����9~����G"���u�,���K1դ�� ��˚� ��PU�D�Z��Ѵ��^n#Z|Ѳ�k�)�����]9��A�7��gRD����l���@ dh����m��9Q
�J��t�Kڮ% e�i�fD�2:qi�W��(<�
ѯ�@�8�q85�����oÁB�,]	�,)�C[��_>��:��U8��b�W��=�3�B�r�5b�-�#�,\.�|Q"&�r֣&�~p�tL��d�r�� �M���Sh��F8�Ȓ��� �?�Ȑ�E�m��g|HY�L	N���#�&pz(�ɏo�Y@}�jEw�6��\�������s�w�>�<�&��غ��_R{��^\^_�g�oo����2��A�du�Y���$�������Ͼ���у�뛓�ώ��7����~�<B�c�>H�O=-����fk��g�+}ܭ�������´L��祍�ɱLfo-�	�XS�Vm�����Ko�<3�ڜ��y׌�O�T3�������(�D�C������]���~���f�W�i!>T�+�1�Fj�����k� F`M����ju_DW!BL�غ8	�%©nd�H�h"���I�i��1M���r����Q�;S��8!��<N�裏��?�4L�#�/�﹢���������X�,�;�=���	h�3�V�F�_c��3�
#����{SKci�z�փ�� �+�B<�%+J_��?pQ=x��a�d�Z)�g����T��>׆��Vѕ���@�|�ζ���,�*���br!�q�Mr�*҅���(9H}B��0��u�G�!N�]2%"�T�JMJ"G(f�p��9����/~�R��DL#Z]��d�QB{L:�Z)8&��)'e�Щ��c���R{��N�����5 k����b�P r�8t��5"Il�����4�d	
Y,A����9�_^f�g��,6�8�XB���"���{��:�<^���R�f���jY<0�6/��z�a�@�`�#���K"�dw�s~���B)z�C ��+b�s�ʓ�Y+�d��5�zg9_�����h�?�6�b��X5��e�(+$�r��M�-��v�p��|
,��D }����ni��a+'w��t�Q��
A��O
gdȥ@��8���a�P�)!d�Cj�3'�N���d�B,}L�Mй�-�6wdYN
�>�r����.�m ùSZ"?��p̤Xg�!�Å�s@.�A��%�hR������wb�F�)a���B��4�M�3��Y
×���VԠ_3pU�������J�Q���X
r�U(�Lf���@�Q�7�ȶ.��m
h�֢1E�D� �+��]�{�p�)�p���Q�,!���No�$��C�*j��	B�m����/E-"�Z
��p�+��L��Ko���
��S�.�zV��!0��A܊�l�V�_tLuY�3�������9�84U�$����r���¤C��)��Q�"��k.Ż��V�oW�Uק��x�"�&�rR��G}�-v�H?M��"��րh��!��>�ꃏ��������ޟf���N|��?#�����ƻ�w7��n��?�������ć=wG�ó#_G�o7�;:<�;>����/iJ��`�Q�Vؖ~}�R=4p���Kd;@�-D�ҁ6��`+�J�v��pɮ�Won���k��|�����/>�ч�������|�����\������#o���g�_�ϟ�����{������w����W�_���<8�����a�޼�y����ų���5�1-)��\KV��0+��u���e	��^���t4�~�"����f�?��ɲF�8��!Bmf�,���WE�,��L������+�@�p�QQ��R�n�u��+���N΁���Y�ajQ�S���(<p� �DM"L�h�a�Su����b��Z
\V��8Q:4��e�ONjp���|�@Τ�9B))w6F�j� ����z������`aMq�cq��Ǒ����_�� '�ȩ�Е�MQj�s���:��U+��lZ{�К�'+�?#������"���D�V    IDAT����+�ZL;@��z�H�t=�U�.���#�վ��~�=�Y�����MmT�!HI0��['ٮ���.$W�� ������H騵W@Y8p�)AN�1�t����)HAV���6L9�פ���J�#R:pN-���c��)w�+�� 7��M�t"��$�T�H	فh5I0�BVDJs�0r�4�鴫ql�U�4��	�r
���_n�B��F~�e���(� #dG�r
l~� S1_:���h&��h��cM��VJ����D���a��'����h�qX`N�Ps8���.KK��á�8!����S�oL:e8BM�wnԏ��`��#}���rDe"RL�9lRE�B��[�e�z�J��c� 2�o���5O��DH�BI�EP��j 8馲ʅ#���B�ZJ�p`8�T���4�%w?+?�2�b��"Ȫ�VYUX|L~���N��uP���ʤf[�Д��Ҭ�t��@���A�-�b*B��UC�)��P�w�Q0�K���CR�3�rj[��Ӓ�̢e�Հdk�hS)�[����uUQ`�������i�Yn|��#؊�Kr�ֶ���, '�Z=˚���NC�ՒE���x�ȗ�߀s5�'}"�6h¡�6Əٔ-%e�����U�&+�E�h5>ߐ���
����XQ�t�Y|����u������!s
B�2-˧-�����͇2��xc�8���uz��9}0�vw{����|����c���>�����W���]L�����;��k_k�����/{���ۯ����������w>8;yztq~��7���^���x�ܺ�Wb]���ܸ\�v���� �8vl�� ��L��������{��SӖ�m�j��=�%�cP3��\Q �Q-S�5�-s���>���T�^����X��8Cގ��?�����g�*l���l��
Vq���7z���U�9Q#D� ޴Pv��׸����(���sp*gQ����D#w@M+���`+l >G�=��w��y�������:������Gu1:�}u6M��3s�R({�&ѝG��<��������j��!Á�dY��י��e56���B= �5<=[�������>�����l��_�Փ4q�@�B�>���-��{H�����du�����*��t:R��5ř��B�j�@�'.ц@���Ӈ� ���1��	�N4Y��HݚbӼhus�L˪.ٹ�ҳ���ױ�]��� SH?_�ҭ4e�8MHm8s zV��=�C��&�Cfլ'��s���Q�!
M�3Z�C����t��+)��8����
u>S6��Ǵ4'-����Z�g�D����q�)2�eRQ�2uY@�B�PD�FQ�|"��:cBjI*M(��=V��~���J�RQ�A9��U)�δ�ٴ�:�8�,S8A+�w��eDI!Û��g��pLE�d����6��ue-!e⥏��
�꼬+�	A���G���DKP�3���5��$�`p�U�O�wls��P���0���l�i~v&��EYm(�7D�X�fm�(�90NY�G#ņ�˦#���!��6�IL�(Д����g��.ʁ�p�,~H���69r�aNo/�z��;I~2���m�h� '@ؿ�j�5u���c�H�,:�U��&�#��X!4�[�N(P.�f+�b�i�B:w��B�X������"�U��I�V3����ą#�eр,�lӺ�"������)���f�2eEW�4�B����eU�� K3>�A���n���'��"p�P "P��Q ��A?΁N"�K߀��F:�Z~hu�wp�$ �c	�vBܒ���3������ �#e]��7�R�C�O=!hU! >߇K������������_h�z����*�'�·�.D=?9?{����fV�d��xQsswzv�*:8��'�>��<��+�!�O�Qo�-�_�Z�תPZm�vz��c��m�֢�?ݾ��Կ��>���;��绫��'����|�����^]�{��_>���o���[�0�����\\�N����/>�ݻ�/��ͷ�N.���g����w��������i�Ԓ��	ў�yY�s����u~��-�q�g�,k1�R�B�(�e�b��f>|;�K��R��`�\��Nu1g �e�[�>MGMnjY4Q~S�I�[
�lg��9rq8]t%��9m&�i�XS���ȚVsj;�h�p'e�Z[�Fh��+���t�P����!��n����97�8�pL�s$b�s�8�g�+��L���@6�Ӝ���q��a��V����>;m�6m��0�����頌NU� �n7&q�A
C㘶]���$�HG0��RXLx�JoZ��@p���Y���������mJ�cp�����앨Ќ�¬%���ǔ�	?�T'�)d��78ӀC�M�(Z�����*���������x�@���%NE8�4N%!�Z�%�:0�U1�a��[,΢>�H�/�TLx�#2:㣕��Ǵ��C��5�p��J�bi|L�i>%��T��d�E1YS�����}}̢�2�z3�U�g�����᳄V�ڎP�#�T(���jnPp�A��a���=
l�C䦐���E�QC��Jz~U�1i�d!�F���7M���:�R��x"�� S^9"u�Y�Uë��%�����o@�ٮ�l�%�^"��L�" A#G.���K��V��'�ڀ������"
	,���&����LEgZ�E��96*?���Zi|��o)?fU⌟�G���&k�pRP����J�P�3�ғ��5L��9�����J��`ZJ
�<3Z��G�T�����83d*BD�q>�j���1:]em0)���L�	���"d`�"ÛN�A V��� DV�D�LW�m�@N�Ӽ�No�ֻ�$��P�-)��V���c�y"_	YuN��sj�k(8��@]���'S���%Fˇd�S{4��ѯ�I/�i�e�Ų8��0���B9��3��~{��Z�L�;�A3 ��h��Y���z.7���U��ܟ�;쮭Y��<����ӑ��lk?�6�,��\ڼ?��N&�z��l�S�~?�n��+�d�*[�|i��}N��0�ۣ�/�o�ۣ��y��o?��8�xv��_]ys��}�}G���;��_���k_���^@��ϱj���Ęeۖ��rv�0NgQ���۽pG�׉3��>^b���@Hd����m�-���ԶN8h��k���l=��*5�L�x4 �~ʵAD
8SU������Z�%���#�c�O%��Ԅ8Uq
�,J!&e�)d*��(�&"�(������CF葋�j��������s��h�K�֡�>Q���O~���J�1 ��;F�bZ�]b|w6��gҩ���U�g�ᓒ�)]�Y2ӓ��k�5(9CD��tX4I�=8�.���[���կ4����P�4��&�[�`s܍�g��C9��s�j���juZ�����$��o�7����P�t�MYQ�BM-D��-���m���IjȺr�;�+$7��n�X�v{�<�up�%��=�c��԰�6�V:}`u���ׯ_��C�`�AQʎ�Χ�RJgf[!E���6L�h��\թI,W�J w��Q��������tҗѰ���O
>��3�6�z����������S��{��FkE���2ܗI#��Z�a�N��!��̑���0-�Ł�N>DM��`����$��XY���Pb�}MxR���xK!Ţ�|���%ZW�s��K4f	|d�Spx�⻿��eH�6��Ǜ"�\���*}�S�-��ԃ~�$��OYh��l&2�u��;��Fn�g�Znys�:#���*W	�.��A �.U�o-8���AKFM�!�O��ij8ӆ)�!द_�&)�)�c�ҍ)�)K�4qN���dф:|�Rhʂ�	�~m�B�B��C/��&N�IqN���)�Ԋ�%���Hu��g�u�6�F?ÔhO��@~�mP�!�9n�ʩb9�h�K�IgH=�[��B�ګO"�~(�>��8ǐE��Fmh�6
�C B�
���,����'�oժ��H1Ⱥ
�8D( �-ʀ��0�,8��{ �6V�ހ-Ѕ�7߇n3�X��plH�4ݥ�@��s���>��v�~���.�8�	���C�KT���%4���2��W��)Kik1:�D�X%�G�|�Z��"j]B�.Xz�7^~�"�ӳ�#�c\�w�g�'��'BG^�����\�tn�]ݭ�q�^!����l�]���/�}���6��H��r����>��S�.?���7�d[�~֪�:d��Z��;C�PNsw/{���a����@n����������7_=yz��ًCߏ����w����_�=;�9����/�~��n��۫������ˣ��o�����o�s*�{ٳ'^�����z��{n9�:
��XBX ��p,P��'k�aYp=��q�Z����;j�)�j��7�"k��i>+N�5����f�M#KG�|�j�v|�)2k���P�3�81�!��#S�龦�1�[͇[qd��rj���B˪n9-ZBk�9l�8R�;4]q�FgB��X��"t
d�2;P�c�%�FR8��,ǔ_�93�I_ԺTg����`�9��m�/o�L��N'S4~�;C�)��N>}W�݋og �Sbėo�B�T�h �L'|`�e!���V7�Y�&�-�ү4�i�Il��@�_iʵ�Տc�la�RY�D:���Ɋ��v�R�$Y>Ć�L�\8g�}hi��ժP���V�I�%j ��B]�V�(X'×��R8��vc4�."�|VoB)����A�(�|��g!��������
ٖ|�F:���}����~9�PU���J/Q��>�����NzR���u����׳PS��Vǟ��J��B$V�Q�凤���I?_�d#pp�\c�J�#q��֔-�'��I9�,�����S4Y��"Y�M
2
�)��BKJ����
�Z���50S|-i�;X-�p3�p>��ң	���4��h�B��6$Z�U]�(��I1 h�(q"��P͔+�1�1%�&�7jƔ[�h�'Lm��3�[xjj%���ޔYYz��uH��	�o���4᭔,��b�t8��$)�4-q���LG�ȘU���օV����%%Hv|�kC(��Mt���d������EJN{>�R"%��,xC��KwS6��1�A�s����ْM�%'>�ᜊ�^Y)d�-Z�DDx:m ����C $����U���h8e�L-~!�m|Q����+�O�$�����t�t�
!hԒ;�����Z��%��ν����ߟi&��
��$�m��7�fj�K*
G�鬅?L}6%8�s$^�h�iqj�~ؚ�6�N��¥@j)oaj�t�Ps�;��	�ޤ������z���5��������4i�2w�7w�gG'��'޵�i�����&�������^T����]�L��b���۝���з7�|��������o�]<}�����o�xzrp��ӳ7���as�{�ptp�%�z�����ewX�O��[]ll��eځ��ZնK��o��b�Şo��HA�Og�2����uRW�rQ��F�K�㕾f<tuzC���zb���_��R���z^��F�%N��! �F��<���SL!A"%�mZt@x)�u�����f�!�iM��	���W,rL�H��^9.�=�J��;��'���?��w�<MZ�����!�ն�#8oYy�d�=x���>{X���Au�=Ǔn�J��&S����mg�.�)��N�Yj�8��S�Ӓ`u����^�q�����(@�nx��Y��`8�<���D�1鈺�-Y�t�|R��f�:>��Zy����OQNL���ഊ��"�%�)�2��PQ~Y Y�ҵT�Z�[]�C�}��X[���b:9��GpO��fK9�:�Bu�1:���%�a)�N?��BͶ�R�#P�~R4�S�HAv�X��#8u�)�Y]�C�i�H4� �U�(BQ4�)&�8�!�UN?���2ԀK����u`]S@�9��WUϻ���ATTR�"�kLy�E+�f���I�R�:|X-�)N��I����ȡ6CWG�]�7eI����P��!k:~�)v�L�:��55j�2_�B��t��9B4�OEC�
�Z�n���d:;��g.!��,��dj��N����8���t�;WK�X{8���c�g�79�N��@C���;��͕�N�m�n�R���Bh��@SE-Y��>�.cQ��֫�~H��d��fn*Wh�n����)X�\4�J�)[���[+TTu�b��T=X�Z���hڄȊjI��X�j�uE�n��Q։aJ����(M��cjU1����Dd>��$��-c�u�*8[o]�<)L�'*�t�����@��?qGMi{k��y���#��l�X��hU�d�o�p�BC �`�h��v~�ZE>���B�pR�'Ro���BR��6����aMkG��#Da�mɵ���r]�.U����IU(�Q������6q\b{���僸�߱p:�HI��X�jֱӧ{����ʅԀr�jc+MYTn��i����BS:5U��j�ڦ�ǭ�,�w��y�.:�/����o�qj����U�[/^�{�tw���[�?��9�Vܟ�|����/m+����6j������m��k!8ehF�Vu��8jOM�t��բn?�e{.$�����]�x{r�)���/O���ˋ�soΞ��;�l������f��y�4>�=�Ǩ�������[q�l��;���+Gٶ�����4�q\X�D�+kԧ#�4s~*iu6��a��C(� ��TY��UG�sF32Z���H)B(q���1�DxN
�+Gbpp��������X��)������]��VBȬ�n� p:�:�,�&_(?�}4 [bc�49Q)�sZ� NbtTδ9h�YRj�J
���8!冏��E}tr+�B�Ajp�l��Ԑ���Ф��BccvPKE���8�,BH���,� ��Y}��6FٴZ�5���+!�1��WT���z+��C�9��B�UNh4[�n)����/đb��S�"�3-��䊦 ̏к"H�z2��31ME�ĩJ���}C9�S���c���1�DK�����h!�05F�_u�蔋9j�|YEN��}&��#T%��T�e����q�EL�fW���~Ud��my��Z��Y-m�� [2� �G��� �ӉY
2�~"��_�K2����*a,?�R��V���o
����N�J�s�Y!:RFm:�ub�0)@�:'2:1M1X����OD:�0e뼔t �����)��-�Z���ԭC����UO��`E�GҴ���~Pr�@09t 5	�������)$��O��6��q�!�Z|4"��@�8��x2@F?!߆w&�ED��8��D�d%N�|�H��t��
4������L|�}�t?W�8����IY4~HRx��������Z��M9U*����1M�J�D#>�)4
)K�q�8�k;|�D���%�ԨD�h��M��C5h�[B�tRE��Sb��.OY8��9�8�(��K!H�|x�l��U��lL�4r���p�#��O�*��EΚR��뜕�������'@m���te%[4���_�(���D���e��K?��O�rW�^�!�xuK�HGK�E#>���v��9^()4*AӉ6��5�����#�� իo/�HyY�t>�)��Tщ��P_S:[�! ��V����^�*���2qV��-��f��=A����.���Wήּ����[������[5oRZ����]Y��#osz3�����pw}w�9���--u��~ٷў��ه_��ٹ]52���g������������� ��g����ݳ��ݻ��������t�#��T�ц��)5��O�}������%[�5��6��i{��.
V����C�j�)8��8�L�Z{��&Ǆ8�/5~�h*�'�JMܛL�{_�s	� /�]/�/���1��Du:F�r�'��&!�YH4���jR:��0����v� *_d��A��    IDATlG?���9��)đh��{k]����[��m�Z혐7���_����{�E�I��@��/n����G}�p�<}j "qn2hJ�h�ub@b�	�E�ǁ`k=��N���>��EY��q2�<�'�p��r�]�)AÉd]YJ�.��$�xUlбz������s�C�+m��@XC�|L���tј�05
����6eѲ8��9���6�_��1ukZ�N	xm�B����8��"�����SS�D��^��۽�=L:l��(=b��\���!:�x��,S�,�P݃�Nfd�QT"\��E=q :d���Z����tKC3���rX8)|Rl>���$X֥��+K���Q�w>�[��ѳl�	�v0-iuF�29��6��j|M-}�e��+��Ef-���T:���"_hK}H���F�*��R�Q���f�B��X>&k�5(`�d+��<�p.���DXG��mگ"jZ'r9��HNz7�Z�ơ���Q�Bd����i~�,�f=8�1!N�ngR(�YKw�|�,Y�D�����_"Y4���IY}��]K��֩O��2�����O�����4���w%��Y���X��*l��U����@qʐ6�r޼�:���*�ߛ-�.I�(��3_��	�C�ѥ7�xiukH$���
K�~���X } �L�!*='Kǀ+j�j[��T"�V�	U����ߡ%��9���Z5G?4!��n�|"��\"̔k�n��B��zc!���\)��I|��%�D)�5)]���i{��0g�(��J?�eA����b�:!%�9p�c��Yaj��u��@����RT�9|d��K�#Kì����y?{\S:�d)G��v�0�)�/U��~I	��򫭭�.RD�T���@�\S�BF�oەv"iL�u�q��*g���S]����Kz物\j;��6����� ���}�ɳ�vC
���5_{!tz�o7�J��<���u����ǜ��^#]_��L�O�er}�Ӟ�kE��ׅ��*�.k��T�o��!��m�:v��9�٦Dm]M�J����h�E�����{ź(�ߋ��п9>�:��������wQ/o���ź��ݼ��yε
��5�X��r�u|-Q���f�ͶC��V
�����e!�m��/d�[�x���?���[u�[�SRk�۫;�������u[�!��bjL!62?<~LY#1𵔟 -)Q���LJq�w��D��6�µ�a�\Vv�nt�pY�*��Ӊ�F�c�_(G��t
�M�EhE�Kʦh҅8�����ʊ��i�Y�ZL>�j��	�V��B#(��.��D��-K!��-�*�A��E3�b�Rؑ��@�����yN��̮�p�j�9��Ñ哂����wVP�B��ɲ�R�v�4&���9E����h
)�.S�H�b�2�!3��ݨb���r�(����4�:y ���v N�h�-�Ģ�?Zu+Y�o��B!Ӝhjʅ!G�N�4����F~�SK�?K5�î�9Lh?)T͐�&��Z!L`m��l��,��2C"��18h���G`Q|���Yk᳢��Zd8�@�3���='��D!80N%,M�ꀍRy�Wo�pH�B8�ìg�6U"�c
��qN�p��*S1f�l:��%f�����9�he�0+đ���f ��MCb�)V�C�s������-�-P�(�!M��*�ݨ�h�W�5qdY-d�G0��Ȣ� ș����8����KLS�>MTJ�Ղ��L̚�i]٘%� �� EYx��@��/W�(�6��j|⤌B�)N!���%h� �St���L)�a��m�9�%����?QS��h��B�kC���jE��D���rE�f�ũ���u�S�:�t�*N]�(M�o�L]�4���6�9s�Jd�Q[ҏ?piIwѹ��R���h#UQ!���-�D4�t����U��Ɂh�/�h��AL�S�L�cD���5�ٺ�,�D�y}�8Y���#��@���A�~�R�<>eN�U��g������PEk:Fr9Iq(�Y��#@�z�Ł�B�8sr�
U��2��ƩS}0�RX��Պ���nwu�B#�׾KĊ-˛�룖G���Q��\_2k߽ih�m˃S�g�.&��OO�c�}Q�I��N�B���q��gn*ۅ~r|�S�HxT�;����������_���s4o��7�n���jw�����g�O}����7�~q�����:�>�}� ��d��>�8�YGu]>�M��;4�m������9���h��t'dL�dm���<ͳ�bJ,Ab%�k��E��^'-5C�Ѐ�G�^�z�WUQ��9��	�~��z��=a&�g�Vh|U�kSQ �Z1��6��� ȍL*�p�}`u�(4��M�5�1(b�>1�V��e8��^Ps����)�oFS�Dʣ0�{���n;B���'6ܓ�>E`�?��C�����J�a7�u!;
��!Ќ�1bǱ�Db�g����)�DN�9�q0��D���J(j�n8Bz(QV��}�p	�k'�i�N����>����|k��9!k���궥��yv�hC)w�UEѭ�?2@���,<�Q�(2Bd�)���Q��3j����Ⱦ��cL����g?ė�:N���U��YS��;g<���8QG��3�����CL�oL"��@��?��cG�P�8�!ź	8�i'*�n�S�����ʂ�
���%Db�qQ�(ʗ��#;���5��m��pSd��[A������f�?�m��P[Lg�����|
i12�{ز��YCH+�8ѬN
��VH���q�еQ
>A�N(�įO>���Oyu���F�4Ł�,X˗�zF����X�`���_�r���7��J;Ϻ�U��+��8a�;~n"Jۺ���AY4��lԞۮ� ���fꇜ�hk�8:���Z�� z���`�Z޴����_�z�˸ʹ:���r�_4�v*v��X|�ÑҢ���ӝxk�D4F͊(����=ֹ*��׾o��rX�M�`cY�,B6���r-G����X"r�X��pN�̻G��B�@��N!���;.�#%(T��tQ8>0[�p��3�!��j�rm�i��p����%��0���v�H9�޴j!jZb5�%T�B�5�E��*��4C�� �㈌I�Z;�E�P{�j�A�N��R�2����`�R�p���,�2=@L]}����\�R!�l�!tR KG��A���N@�4д�[+�?��RD���*D�`)��BF��#��'���ne�]�U��������kP3|͠�$�z7N�5��ۿ����bYS"R�	_-�8V-�pkd�
ٟ:����6���D'�ۅW)�^�������w�.�����:�׷�8m|_���'O��^�R��/>���/�;圃4��y|�>v�������vC`)�4;��O��HV�^�)'�8�7�vH���o/����]߬O�Z�� qdvOζ����9=�Ǭ��������~q~���������w��\߯W���|Q��G=�Q뽯Ĺ��HNi�Zw���=�;yt�UBW8��s!C�Z��y·�-���!���Z�v�L���R.ע9���M֏\�MJ{%
1�<
�I׀�h�G�r�ȶ�ɂ�b�9��E�I��*���E�������wNV4�>y� �%`�&��J�����Gn��m���R3�B���">g����Gv��]�(-�Łh �l�F�3�9����$%�/kR"�qLE�O�ʪ?�T	�n�O�B��|�E���P���)���!�vbuPF��L�"s��R���O��"N[�騅'�́s��ߔ."�h�ڔ��L`��z�&�� �d?k�{�PF�̦���JQ�8mZ�)!�Y-��S��XN����F $��Y2���r�ǆ�����!�Bz�ĖC-f;��40)H�F�%�Gk�&#8��Y!�-�BUX��k	����8V�m!i�kC.J!V����۔m�k���V-x��v����Y�t�[�Ȣ�$?A�D`U�m���J1!��(�!��1�ǋ
q"��?�b&�Ģ� ��U�Ҙ)f̈́C�Jsp0�h[�a
�Z5�Q
�o���)=��@L>k�\M������ j*:�W�r�m-�sL���T���
�n�s��}��i@'��L�H
����'f�9�)�ф&1�5��a�����EӁ�@�h�N�|�+d��as�J�f[�t��JP�ǩ���Y4�@,�~L1󑍙�2�4ж�CKM��R�: 5�9!�d�S3M\���� F+�����!����*T��
rK�������`É'�4-8G�����!�(G9d*��LE1��1$F���>o��ь�S
�r�� ^�R.Ostj&M��Lǔm��FL:��N��r����l�8���xu��p28F|SY|X�L��p�^y}�2k��Q�ʥ�'�_���:«B��@��Zl�w�4e1������S��Eᦃ���)�v�k�p�jI�C��UV��8U�.QVu�SH_:�ogL��k/��1�Y�A0�+��@/�]�dV���5��f}~r��Z��W�w�u֭�V�6����G'�}�r�����{z~�I��zs|��F�x��V��|r�ٵ�=�L�Q�_/
G>���>���ͷ>����֕�s�'g�ώO����o==�����y�{w�_]�������S��\�j�sM�MGA��p��~�;u�d;����wD�mc.�5DYv<��T���6pd�w����98B5�Aև~�����}�{��jY��c�{��(��!W�k��
�|��T�}���	�<r�D�7�[?f
,�D�,�8q�".Ħ�bj��
�#����	�8v&eV-Ӷ��c.7������g=��A[�W�W���yr�?��;�:���ķ�8^�q�z�����Q�6�X�Z��4`�C]~UШI�#(D�����Y]k]�
 B; ק�{p��\�M��`����s飏>�j�Oy���kC�LE�Dc����dE�p����FII-�PS=W�@�Q�\tJ��#���rr!,>�PuK� d�2�4�Z���H�,܎w:�d�-�n�f����l{��[0��pM泎�(���:@=�$�i 8FЁf��œX���zx͎��V��J
:*"HD�Y�LuK'k��q8!��SUD��O�c�3
���ҝ���?��?�V���UCaH���{�m��:T����(�h%��z�0}��2p���lq�q�R藫S���mrT*��h��8!mAR�F&eڎ��F(a�kLԘt8Y`4��Q�HD�frm�v
&����U�K����m�'�����k������ܲj�:уQE�DYp���+Ӷ�_���?��?׿�2�y|O����4��A��oiȤ�<� ӹw;j^ioh�z1�C
z�>#�\�U��4f��n��u�ҘE�
��{l���S�@d��-����j�ڳ
"�@����w}R0�0M;0�=&PE���,��i�8L���G3e���;r�u�z[#_�\�kXiN�Y�ǟʘ��~�"��r��+Z	�gLL���Z�,~Mj��j�u.�1�lE�F�.>��\|4����|�E�NȆ\��>;]u��U4���C�,�������6ik;S{�X�&Y!v*�	Z�)�f8z6t�z�tv����5��h^�� ��<���$B��_��}K�Qs5�s��8�;O_K��s�1pT�K��]v�E���Џ�Y'*���^g�,"��V3t(��ܶo�_m�?��r�\���/]4�,D��dvh	�t���z�+�MH�����u���F�Q��������z�������/v�/|���37+�hO���^�|~�p��Uj�z��I�,RJ[�С��;��V����!1�F��
�2�<:9�8^pԌ���~8�ѝ^^��)k��һ��g��!�nD4�OX�+�r}	\�d}U�vg^��,+Ŋr���t�Z�+�Ҁ��LA4>_o6JE��T��1��t���H4u�Xl�������JTq	=�du�ޚ�a	Bp����a u(�G:����Kt��Zm?!߈ƙަ��V��0+���1�h�]ek�&�J��}|�Bbi����!�)S���o�"5i�)���N�PV�B��}����pJ�K'U�|4|�W(���b�o�Cx|Q��V����XW���,>e6B
B���g��a��4����JL�����5�E�S9�hJ�.DT.��'�Lq�F��v�z��Gb����+}><�Sې)��S�|U��M�/��˚��ׇ�
���7�Mk���z���������	Uq��G���Y�ⷄ���A3�-�3uM�q(��lY@4��+:h�9��u�3��?=��B|�T��p`��A4~�@�I���I��*Ѥ�Nw�Ԫ��㷺��V1LU�JԭiY��p�ָ�.$���ֶ*�f��m!駹�)X����@�J3d��pu9�ʶE���jk)���̯�IWˠ9d:|�r��mۘ�0�S��7ń��1�p��?nR(�o�H%�����K�?r�Wͯ%p��Φ����٪q� Y`��lʪ>��LGYT	��V]Ԕ���o-�Ŭ�|Sf�#���J9DJ��_z ��lK�|"�4A��:Ǡ�V��9�
�S��ȂP`���J��z�p�O���B�4�y~���RnV(��O�e*�CPc�Q�(_4$YxN{�Ri �1]+��d�Y>'�*9>��|��B@CHv�>�-|48�t8���E�����p E%��ijT:�(�\Μ���S�_��3B�~��OǆTT4e�,����U��S��hx�izy�%��-NgK�(�!b!l%Z\o`���q����IS�49~oO�UT(��?�ܚ��`������ڀp�,E#��P/c���^_#c�g�qj��]��B8i��4q�I�� W�G4�w�f�7Ğ��|�½����K��K��<؝0�]ok9�Y��Ŀ��c��������70���n|E���b[Ѽ<98����x������ݭw�nv����������1���"���q���n�����z�S7��'�M���g��/�=@��'�~��Ց�R�?z�;=���+��o-A{�Kt�Fw��o۪׵i�������y�a��0)�,���R'g�ܙc�=A%�_0��{��������Y�#��1��cPc�}���'��xiOЗ3{��ɀ*SQ��L'NoA������C��s����Ŗ��,���d`�κΫ,P
�ê���HGT����FQQ��`R��e���M�Vc�!8dX��)+��y��6ӳ����v l���	����ɡ�g{#�����"t�rp��R�b��OSVJ�(���c�ѧ���\{��,����tp�d[����	�h	��`ф�Q	� �����ASgT�4��\cV�!�SW��~���>���]������?�	��rL;4���*T4�#����,?�E�؀R�#k*
Q�?���a�^�r�8,P������T:ۦ�h�����DӢ�L�|����vҾ9(6�۷F�4���!�:X��p��r��>�6g�Z���W��U���~�5G��5��P	YM�۟����!���)�(R�i�[���Y>�,S��X����NV
����Fy#I�|O���c��Z�O~��tH�$�a�HZ7���B�ƄԟJ��m��!�;�҅ �� ��[b4��(d�ŏ��Jl`�5Tj�2 )�!��gY|V'�XRnL|;hg�+]	8���q'���y7�d�}t�����#˱p�Ȋ��=��d7�-͛�%7��V-�8����f�D��[ќ
�(蓸ꬨ�PT���Ch��KΏ[�jz?)5��s��?A�qY��Ӊ�gM��*���yk�6ĴE�6��	7�@�pl�A�"'M�ט��z�i�mW�8���l;Ɨ�c8�@�s �>�B��RM���>�=��8ᆅT��
�()
�k�V�@:Fk4��ph�k&A~[�X�h�l�I�L��hmt�L5��LM	|:8S��!��u+
�X|��N�    IDAT?�D��O�4�t�h.
�@�&GϜ�"�7�c�nc��ls(�u(�rL]_޹��@��E��Kܿ6�2�����>ե��`9����#�io}�% G-�P������ҏ&��-��Ǘ�vE�SK�b`��M�@���ʹ!p�ǔ�T�o������:MK��p�}�������aj�D�|)�p�� �)���wh�1�9���`u�-�� 
N	�WQ{-����͊��,�c`V���1���GАkj-���#7�(�*����1�-qݠ���,�4����l[��!�v�q1�tN��)*�uh	b @�9M�?��?���O!��u"/ю�u����Q{��1%��T�)�p�FD�W�(1������
��q��%�(����O2��&P�5��rcNi��Y�5�E�M�,$Zj@���Z��:vށ�Iah�M�a]|Ⱦ`��,�q�}QxN
*VKQ�A*ZE;O�W؀L���s0�$Un;Y)P�U�>�8�{hI�EY">g_���2 h.�����Д̗نP6EvK麋	IV
�)�-��7�au)������ũ���-�l�&Kb>)w��]Ő�,�]��67�&�}�|
FӘ�t��Ii�'ma��94�t���L9�DD��4Ǧ3]5�)&�M9|V(��Ъ���o������Z��m���(B�Jb��FS�iN~4~�o�UD''D�Ԡ6��GC0��k�"��V
��#xݲh��R�����||���MG
nJ$G�h�f���6������e�$�1xvpY5L�Zl�F�3�R�4���o�pLg{���
�m�gQ:��FY���p�YK�Bb"�#K(��6�1�c� D3m�l�"�*i�,|^��O�5	����S.ܔ�t�B9c!/�֬h��Y	�ɚV�S�h�K��[�+;��GP��ύ���b��ԚE�V�Sb�z��(���=� R����)Aٙ��CbZH{X�r��P{��
a�\�@�j�D��7�ZDuQ��V�d���2��hSV
r��))�8����	�n+I��Q�7R��a����~�ƜҦ�H��Tn
�χ�ki~�l7Rh�L��Z�^n;�VT�k�6�l�����B����85"ʑ�<+�����!���V��1K)�?Y�,�S���K�|��X)|8>�i�2��^�[4�R����!v��!c�;c+��U3�U�#�mZ�q���W�R8g:�w^i,��k Y�~��E��"Xrgl�4���\֪�x|9�k��\Q�P�V�;�k�E�b>;W����C�ۛ�Kp]�2�V8ާ�B|l+|��Ʒ�R9����]������o�ܮ�/�n=���}Mխbw�~K��¿���;���VGG��	]߅�*��z{Ն���/j�>;��ݜ�n�wW���q|����w_>�[��N/�\�|O鋯.O��<��=�=9����G'�o��w�]^_)�t#���P�6�O�7<��{> )���)��ꙒD���t�j��g����BG��#�J�����՛g@S�;>��c!�E�x�͓ｱ�����=����hL�3��U�#��Һ�Ƒ�[���%�9B�p�A:��I�9���O74C�D����u"T��\�/ 9@ƿQ3��-�q�թ�����;"u��g�?��ϼ��%_�*����G?RB!H�{�b�_�n/.j��K�e��E��p>Ӗ�`�:��ҀiOx���f)��G���R��)}x'f!��Br�m���rr���ɖ������zp�#�y���}a��c�Y�
i�P�B��#�2��4?��k
�Q�L�(YN�?�Q�G��d�DK����*4`�ۍ8,>)��v��\H����&xg�m�|�N?��(+J����pL��dSu���up�+�=�\���S�az��[
})��S�a�Xue�?�.k�Jio�7U]]N�N � �ئ1�!�N�Va��LΡ�|��V���9�:Y���|���]��§�{T�h�Z|�vA~k��J"��镣6)5"����-Ac[�h���6��Ɛ�1L�����p�s:`u%�4����mZN��T���&�\;ϐ����fs�*$$�T-C��~���gղ!����K�8l=�'�&�QEV���f������қƈt�T7�\05 ��猪�؛*���M�4�G�)Ρ�U�e-yKU�lh̛����*eC3�8�[��{�SKj	�i�Qn�*m@����*����N���(�q8�XŶ�l�l�0�4��Úa�`	���:���Q U���/��j����J1��^�)G�f1��i=[��h{Y�-���APT�����[�ҭ���`aJђ��,�u%(��(�����p��G�,S:������������l�s(�B����D����N3�@"l�]��n�!W���Z@MU'bgE�KtY��c�%S�v��5U�w�j��5�c��p��E���r�i�>�3���O��	)KC3eM�Sd[ćS.�U���+�0��.8)��	�=�D�]�I�'(�rd�է����)('�PW��)�ZM��hZ�7
�3��}���ݔEn�~6�'A
5Utȱ	|��B:�DN�n\|���)��Id��ijh:G���Ƿ]Q�`�͈/ʧ/�}��K�^m��+K�>9e)j���\�Y�s@�r�@�_K8�pR���/L�\���4���]E.C�DX+�����u�QQ���mH�7YR� ��Ê�I��1�s��� %�mݺ�p�+�T��)
NS����2M�C�Q!~�W�#g:
�$W׀+ѡ4�R�Q����i�l]	.K(<��:�mN�h�/�M�1�Bͨ�ڐ++&'�Mܩ�Q�X�:��V	`�4E���H�Cfu�PP+�pVJ+��D����5Y��|N"�Z��+���{1��K�$�"Z�OW-*��5 w\�7Mh�Ň�	�H�m�K��bZ��m�D��-?��(n���4����7֢E)[˴� ��)L]��C*���4eô��g��
7��Sˆ�0!N��dcHm������������IG:��	A "��E���a�r#�9@!~�ZE5�O�c-�('_������r��p���sz��t�($"J�-} ||���at"�J�u6�A�.�l�[���8��S�=�����(-Z���ZTN��Fo�.��B�50�NC�H�,�;�jq��hmdv�����*����6��Y f:@��T�1�-�Չ"���l��~�V]���8=p" sX�l�zPȴ���|�p�F"@#�MqL�r"���2�S���.��h
�<"����@�ͪ���8t�QB!۝�mAK9�k$�U�t7Ch8-.wJL?6���l�Ϡ��׽�Xv[�{����V���>������@ � ^��`��uԧ�����ܙ���^*����1G�s��Wf�];S����x퍲V�5,1>&��W�&\
�%�q����Ȇ��&E�Z8BR����7�U���7�8I��S��em�ZZ4���U�1Fp���N���F�muKh�j!hM9����K�s��G���T��-S����aq�r�o�o�^iQô(G��㆟�y3��R�9\uʝ�t �=j躘����>��Ġ�)|���V  !3�j��¶��E>�:J�Tt O���g�6͞T�8����~fd��,7�l՛�A᠅��A��cϦNN��s�ÐKv��������8U���&�#��#$v�-N�f-���0�ۻ��ǧ���K,��<��7,�!L��I�xpy|yz������wAO��DO��uf�`����]O�������2os�����>������W��?���g����W߼�/ޞ~��~v�_�����R=C<>�8=�ˣ���kgK�v������Q�����<�}�[��k�]��8Hҩ�a��h�1=��i-QG�K_�R��<�� �[�~5�믿N�g1�	�Q���W|"|��A�Λ���F~g@���tժ��5�C������j�#�G&T6b�E��M�Z��G�"p*��mԞ}�l�L�r��Eub�G���7��ˍ!����������ZO*�~�����r9(�u�c *��wX�Ƶ�x���K��R���1j=N¬m�$�ѕ6��f����4j��KA�SÉV��$}��miz�:ãW�8�R<U3��q�衮��|h�׿��D�ID'��m�+�*(l	qD� ��j�AϺ�6��-�%"d�M�l���Q`)�÷���#*��Dk $�T{ɡ�s�K'+O�~�3�箬��L�{��>�����!83�Z�3�h�PQȠ���߶��1�륐��>��E֥���]��Mv3� ���j(BPBl�ק�j;"�#'�g�ZB�R�U���@L��1�cir��+��:�޸E����<)�����	����Be}� Nڑ�T����t`��!�@V
2Dj���b{a�/+\2`x�z� 
�7Ճ�H� Ek&YH��Fh-�8�qD솋��Y8���	�L�)�Q�f�'�A�1RQ]{�`uP��1�����I��uS���T��&�p;�
!�r]�n@8��(j���K�r-DHQ|L��D\��e95A�Ȋ���^6�QݿZrǱ.4)ʭ�B��k���lP+]�ƈH"�R�s)!�!8����Y�>+*�1��N�vCuL�p�Բ?��
7k:�!��Q����҇���7S�.J[!�Z�Հ�)�>��@�m���y�C���]D�� P�r����,GE��aW����V)X�ۙv��Y���`�'�j�WQW|�Z.5N<�)����2r�h
����o�ֿ��@�
֢==�|hUTQ�ڐ^J֎��C5H�U�+�φ���4I!T�5�񭥶1���,�)>�t�%���ҧ�H��,��UjZu�pB|��<y�(5��D+5u̪(������ �80�^צ4������Y�i����h-:Z��k5��Xj���7�t�J�.K��t���qu��)a��jY
$5)ĕv� .��@���!(�_��wۿ{���������w��sS�T`j�-V�qd�|�����	�%(�C��!UcȆi�|+���l��$� �)�A��c�:ҁC+�8S�@�O�������/�F
G(k��n̪�e鍲��|�������{뭷t�ίI�A���N[]!h����]^|��k��SJ'}����Z4͔�N���r���KoTn@D!�к��9��*ؓ���\"h|N5�4�b�*�U�@SxULk?ͪ�)ji�޽�NH�g���B��#�Bm�oR�r�Z/b��2?ALSQEi�9��*��Nt������:�ф$��SȠ� ۾ڗH62)S����Z ��8l�����le�O,����q����ξ��^S1d!G�m�D��FI��R]ϐb9l�SQ�,GV+
L�t֔5����D��U���\"p��l���IO���Z�Ш�Yޅ(K:d�8
�AMV.��9�Ȣ�X'��BF%ʚi�,r�5��\|�+˯
B�Xh�͊:%~���l��Q������-9߱Wq�r|����SV�,?B� ��^wp���V.ߺ�����?��嚶|����!e
q�FDV]Uδ��Fn�ҥp Ώ�|�pN!���FQ)u�̯����T�\QS�I�T��W�%�!��r^bN�0+mʇ(�0�$N2�q�槆��ڤ�DcMu�(��D�;%d����,>Ψ%8�7����(}Vѧ�DhrD�釷X~G�/�_V)@C�iͰ��E�RTl��ƟrD��M�Em:�&!�B�IP�~ 6�a�!)@�!�p��I���*�A�%ݿ"�(�*�4|�}b
BL9�9e�W����d�/���t�넚��
!Y���'U!>>���vd^�����T�� BFSu9@�_K	�� ���t�b��4��*T-�t�
qJ�(�6E���t�iBF�P0br�8� �����^'3�	,��c���'P��y��!��T�t��H}�Bf�i�E�	�)�����o ��~�Z��dq Bچ��W:`?6��2�V:���|���Bg�)!�#����?�;?ٞ��P���i�]����K�z�ӧ�%x}s���sESw�_o�v�Ƈ<϶/�އ��Z�����zq}��o@�M�>����0}Q��������~/�U�=�<~�>�i���΃U���jϏ�Z�g6��[�GJ�[�k>>�\�����������?8?�����.oo�u�h}���_�����ճ�OD�Y��핝�^��ɶԐ%
�`r�e��-�uA��8pȇ~蟶���<�󰑸 ]�w�y��/;"��j�+K�c�<������K�B�#���#>��4
q��T3@��Ѱ(ǀ���ڐ�۴\8>ܔ��#qIl��r�u��"���,�r�4Y!x��S�(}�Iж�OQ%�$���ӟ�ԓ:ۋ�cW�n��R���ԣW�:I��`�[d:vX�!
i�r�Y~�v�e5�R�E�)YW�PLj6��
�,Q��7�h�W�N��BS �9iZ�P71�\|��!�:x����m�t9`���o��w��]L[��r-�&��p�~���p����|#�G	�9��U���"l�+H�5��F�T碐t���[#&'��fv�!R��������+Rr+��1�g��W�u-|�����7�?��,���F�B����5�8.�����6����ĔE04L�P]���
qT�k�m�|�|!��3j��cr�6*MS�(����y��GĖc7bJ4=sߴ5�,`����A<B�c���2z��A:���W �5`� G!��8zE3p
#O��crp�� B?^�R0��Ck��� �M�@ox8a�� H�k8v��N	�YS�[���j9m]~Y)�W35��qԀ����MwUE}oD���u�ӕ,�N#מ�r񕮊=�`��U�q�5鬨R�]tY@:�U�d�4�h�rzU�B��J���"�!6Mug���D�b� r�L�1��Rݪ���S�^�d!��a�D�ĝm�v��I!.d�F��Ek+(�Yt�%��H�*d��<&5k�?�)�4E-�k�ҕPb��F�|!�U]��-��o(L�I����-��~�[��Y�궫��C��:%��g���ys�lKmQ�Jϱ����t,!�Nc��v����쾌��v�A���zq�p�:�p=ӑ"Q��t�F+EFS�����94�g*]��0�d��a�.�����|L>����7( ˥�ӥ�X����z�W��!������w�\����:!t�U#�ȊZ��^��L�+�&@Z>ߩйZ�� DL��2u�}����}�hQ�G��E�^ho���{�G�5�O��]T��a}&��L��Ҙ}��k��	QQ��Wm)%*��ԉێW�De9����щ��E��o��	"�H��*&~d���]G���7�I8d�#�J���tG3d8�X��"�� q$&U���m��5�=�D��^_��h�Z�Ǵi�^%�)���S�m�A�O>���1ek�����h��,
@)�hʡ�"
r�	Uh�����c�Ȕ05�Y`������>����"�[/Sv��O������o��׼GW��V�-��"j$R�h�,Y��LH<d�L0�e�kBJ�S?)!:�M�^�ҟ���1��Ή�nT�C����0%&XV�Q�%����*�_"�&��,���������`Ee��&=f-%ˊʭ!h*�Z)gϤiѕ!*��@��f��E��)N�^j	-)Y��ѐ'=�YM�'�(��'��I�Pm�C[K�LR��+�*�s �q���b��7��J7�ِi���p�&^?�����)��
E�c+��t>AL����7�r*ͦY�T���j���8k_���Z
G0j�r�E+X��U��B9�6l�)��M6�1-�j���㗲���s�R�B-���:iB�6|.\.�h4�� hFA�    IDAT�Z-Poj�T��� l��F�a"���Չ����!��>]�Y��/7e�+4NM�M�SR��4�.���d�Ǚ�ɂ���L.�CF�0m-qX),e#Y�$D�muM��D��*���qL���{�%�'�6�4)�3D�0e�CbJ�	l����Y|c���#ʪk���K���I��Bs�&��Q�T�Z��Y���o/m)Pn��1��B����t����>g	���et�3A ;R��tB��d+��c�J?�Ȉ��8��F�U1ŇԳ1uDMKd+�k�5����w5�X#��A��ko�h�`�.��)�B8���@~
pȀ��Ka���\4
B�!���4�d�c��I���zjQQ�8U��2q)i����_�豘y(������K�L�BSH�f]�Z�x�$��d}[Y��YE[&���b��pL?�&X�BME�[�+���U!X!=[�u�7���}G)�|\����b�.��ub�W�����ѱ?�y~w�GK�����{|{v8Z����h��X�V��]G;tt��M����W�O[^�3��7'>}�>i�w��+�>��t=����c��g�wު�3�'~xvX�I�k!.��sys�֏��yqw{|���ۥ��?}����\]>~�������ë����<���^��tΞ?{���f�y;䪯6��9�˶�]G(�ó�j�^vҐ"4H�nu8@�t�wU�����e���v�L�ӄ�2u�=Qݏ�(��D�<�K���.���tX�~���G4ZH| &�3�N�S�uA�*��%�L�&�3��AjC�Q�%�9��!�6?2+�q?�����?��O~� �v��{8���7�yZK�3�r[����uH���Z���r[�V���0�;�
�<(�f���:Ua1]_���tE�t��`u�p�$�~��@�G�n��8Nҭ�ɓ'o���m�����9�/~�����Q��f��_5� -���5U���*�Bd�����0M:�O��(P9)�H��e"h�Dd�NK1��S`�6V���%��S�ތ��-9�(��\[�mc��>�U|�F���K��v�W�V�[��_{�5�B�L/y�]>%����ҏr�a�SC�^�P�,��紷DZ��ٙ,߀�C�r9l=Dcm��y3tk����J�(jv���଻���t:�rԐ6�fu$���]���@"��v���Ԓ4A�r{Tg��Le	QN0��i
�hD�5c�l���"��.��H��'�Y!�^o,���n��ǴEtD�����r#��6����z�,*��S��j��f1]0��}ʺe�J���~4�5�y�j�:��UQW!m�$R�	@�#:$.�E��5�bӹ��|uTWW�ݓѳU� :q�|M���B�-�{�re�������X�bC�m�AYԺ|��*.K:A
@d-I��ݳ'uKJc�t��D�N������#�ŔN�#��@_W����n�H��9i]	IGku�Q��F�4� hr}��g�����b-|S�ƈ��=ʺE3չ7�d��!��k����U�(Q.ǰ	Dt_��iHѶ��d�Ⳮ�M�����$��.�M��RS:k(!���X�}���m��h�^)�G����/9�rR���E�e%qP;'����决_���mXMn
^���^�m��R�i!��]�^�^;��*-ĚN?"��;��M5fu@�4�����>q(�})u���f��)a�:$�ATWhZ�=+To��!SQ崄���~8��`��1���2���=�j�V1�{?��#:B��1H�@�����#B���RLU�4է)!)-UnXf�RpXY��BtE�uU����Y���jt]��� _	�jNYv�a`���q*�1����������d���K���&�0�1��Lb	��pS�:I�o��QPH����`:h�t8�)��6���83����*'�D�� 4ۮ�f��"�����P��k�@��J��dq�|�&Y~9�t^��u$��L��J"l"����qHe��x)�h��ֺ8�Y���A÷9��P��L�s~��ʭPvDL+$=��7j�M
�� �W�h2������v%��ī^�j�őhᢘ%��M���WL�t���9��Pz�d[��^��Z"������Ӗ#��Z��|��B�\3�J�@�����/b�Bx	"��_:�Z��_.��}>NC.X��]8�h�mr��s%V��ZCڟ�r5�+1��mES)M��P�JK��)_��pF���Y�~Δ�(k��")�Ch��5R�^I46ɵ.`6P?����#$�S3h��U�ʭ+C�)�&�%�sJA58	�"
�#��!sA����4�4�gG$�Q Y��p������h����u(�����o���Υ,k�Bj�H���ɧiP�y��)�&���'f����@L��,G�Q�ҁR���B�ׅ��U��j%f�F
�ʟ�D�]E����Gٮ�����!��7E�k��P�9�)G��ɥ��tŁs��F�/m��ť��U��-�4�m���"��U��zM���дā���-��@.�5���D��*��n�B�h��,o��v:B[�e��z� GR9N����E���{�il��.J=��~�%>k���'��j/��P�������@vK�O'%����X&P�%�t�b�
>�DN�L�ٶ�i[��L��R��%���W��D�	4d�-���yT�)��|U��$�
�g���gӘlU�hlxS4w6�<��
�a��5�$btݭQ�$�I�^���
G�h�,5�0�S�#�w�����1��i��r ����N�b ��5���#��,rvyq�W��W�G�]�m�~h�/���.�:��8;y|y��������_WG�g��]\�����/�=������z�����	������_\���z[ru|��<?xc��/��=�N��1ׯ�]�����@/N/�n����w0�O��s=<8=��+���r�/]?:9�ǳ����]?_�>=z�t��}u�VѩS��X�gM5ӥi�W�ۆ�� �I~�U�o�zV��Rœ"�U��B�h��R��b끂r�:j	y>�9B��UuYY{����-��D��@�a
�_���(Pc�����\%J� �t(T�?-�8-�nIM-4= 9@�kͦAjO�<���~�٬P/^���ײY~3�GL6��C�J���I�3�*�p9X��Y����I�b�>p0ɲr%J�S�r�dKii��K��JJWKT�sb�ƶ�
�SYb�zҋ��M�D(����x��_��'������Y)��Y�iȗ>C4Bu�Vt�8��������&��A؏R�ÔH{T���A�2�5LK��[�v�Bu�%����'��6�>�9��������Ǖ��(�=Q:=qu�!L��O:u��,9�%R]ֹE�am�"� '���i���UI���(�\��# U������+��e`�*���鉷��{W"��[����s��v��� ��� �F���8��]��b�L)HY}mוϊ�ZHۧ]H��:�i�5`�i�H�X�!�N��(
�c�ε�X���"��kL�n���B6%+����oE�Dmx1;O�{�A�FJuNgZ�&E��>FEwL�ķ!���k�m�BR�J�~4�wB�ӗ��@֝�� �4uX�p@���J��[ߪ}qUN?�O!H\?��(���ڍ
�1Hm�\/<_*�H�)�L.�.�|���\%���9F����hU���֢�,!S`M�|v6VuR�];��v#�.�R�H^ۦp��E��MEk���|�Y8���9�!p�Tu)B�T�7�%S�EGdVh�V!E�R6bZi�U�j>�,���pխ��?�` �'�����_T�����jql�1m#㰤D�MCw��%N6�|)eaF0%E�5,����n���(�r��v�&�ey#�;�6�_wG�I�Z��G�DV�40�y��}����:�,�{���l��н6�r��T��,�BZ�nS&b[��Z�QVj��P)K󦲤# MY�x�t70�X�Vu%�%��<q1�z�d7� S��c���9-J�z�L����Q��	9�5,˝
��*����y��B� �bׅ,������1��PQnS��O�/W4K�~����Z(�i22CÉ�h,Kk3���)��`jՆfZ�B�|:p=���;<F͸�+G�mIJ�d���cچh�**�&[K|L>�,�8�m���sqD#�o�Jg�/K�6��B.�T7�J��	�7��6�T����B��j�ۖ�0%p"gq�h#�|�oQu��)�&�"��UK�cV��P�h��#� D��R��� �� k���l�ҐF�c�I�X
��(D��~6)K�L�i�J�EQ+�S�7�,k+rH�jZ)+Z�t5U 59R���O|i�Z��`��B"(D�(���j�U��hS1�xNYYe*W�Yͭ�u98p��Ӌ�d���\�c���k��ŧ<餚��V��1H�@k��^���Z,��lCT�h����]eN
rۄD�h�拆S#��5�U��VΆ��E��t�G��5�C6�:eH͘e�k*d$���H=���-���)WyVѢ�ULGJ=��	��uX�o�|�,�M��#h���c�끳���ؙ��B�'>ʦ]��S.=N��(�'�*�5m�m��8r��Xn�e�����M`)h�~4Έp�����!�m��D	�A�U>~{"$�hR�5_QY��Yc�ԭh=�f:"h�]��z��tU-�Q���sY�EU܂�_�p�,-f��R�BX�����8�ѷR�c���5���8�j�T�	�W�'����N�lj٘�Y�#w��J��b"�b�օf��B��4�'۔�\ɥcpdq��b-�@;��cp0�6fSH>�O)�@�:J	d#$�f �mQ�Y;������QE�޵5&���\N���O]�e-�� ���͟�!��svDT�cچ�d���c�bY�l~�����4P�2�h-���Mh�^Y���w��O���\�;�F+q_���K�1(�P؏6��J�p\&�v �i`S���`p����>g��1e�ipLS`kRS�Y�Gy|O{����f���t�6�1`R@�p燯мR����j�5��8��"�R ���5��c�^v��W���#�G�|�ٳ��z��_״8,�#��[��J���'g��g��=�8;}������*�ѳ��g����7�uw�wݮ">x��Í�w����;�W7G�g|x��_�t:�{�j}���L��T�zs�҇A��ZY�=#�&9�}������ˋ��Ĺ�����������_I�ޓ�������C�p��g7t�ܴEm��\��]S��ط���9Z.�PW�q�pW��K���r������R��Iw`z��U5�i�bRVB��������g!Ѫ���bʡ��g)o��$�������r#��bcBFg�m���P�On�� �Y8���OW�?�6���(я�c��m��y&���_������b�=����	{x�JT�#o������h5�Bz�Á��P3��!�q�=p�_z{h���Gb�ZpCu"��n98pHg�u�Q�&�1�;'Fi@�'�rm�ĞPA�N���o#����w��[��#{0�z='k����!��� 1��f|N��`BL�=QN4�#4d��R$��[Q���
�[��3�zK�~ �he1];�p[����"8���6�s�>"��� �м���K�\ǲ�[Y���C\�zc�ڃK!b�.S���!�s �8F-A&J^zQY�`:̩i������a�N���ەeE�?�ؓRjg_��Wz�I�.K�"�z�*V�'���R�������!2����J�C(���	���4�)�F�B��1���`�q~=����F
��Yj��Z�h'��^ϲ<��8�����qsT��\/o�f��D�H�{�,��$(�e��r=���r�zo�x=[�,G:�W���=B�3��������8j���m�'�~�6t�yۂ�{�JX�5),��f�� D1��E�:U�v�Bt�>ˍ��fo9Fj9z�M�\�l#A4
��2buK��J���8v�V.�f�4�B�����2��l��&��n�l��t75�8KmV���_�k�U%\
�����L��ڬT������[�� �A���{H�4�\.� ��h|�|�]r��'��dI7���t����ru+}�B�B� N�t��pRdYS--�ƚ)�����e
I�:UB!S�F�l�����b��;��1A�I��bѤӡ&ݞ#��D�t?����צfd��<')E�[����p����K8�)�V�b�"c�t�*��Z�h9~~��%��.א%Eot�����K�o����'\tu��1�X�adCB,YK %�Z��\|�x"Q�΋"�����H�ńoݿ Ӭ7]E��[)&$C|�p@�Bh��w��;��+��*��ڶ�l&�!Z�t ��l,_��4H�����<�wl�U�HAc=)�f��QԦ�B�7��[�lkXT�,��c������L�I�>:41�e�9S������I��4|r��%X��tDYc�ŗ��r��z���1��Ҥ�s �i�1M9�ru5����VH��T��e��8;�������ǩ�D��sY:!k�2�]kSx{�~���O'���p�� ��T�_hj��rX�V����I�[\W�i�����Y��c��:��� d?��d� 9����,�B|:*X��)B/R��e�9�Ͷ:Y]�8�����1�4B�8�SV>[�����B�"B ˟W��I�B=�|�V�4��N�/��o�3��j�T���>NE��v�Әc!pC'h��8[�V*s��f	�
qD�9���[)S��V�)δ�f���M!ULY��R�▋�1F�Ϧ_oӉ\�ā����q�b��g�D�j�i�1 -D���$V���O�@c�Y"��9�Ef\��a*���|��>a�������tr��rN`��B�����	�Z���r��M��09t��-�������S�K�O����S�l�ouJ#��2ptځ�MSc�!	���d��>����D&�,��a�ې��ߊ8q�SK��B�����o�9��B|��$���1��#R֤H�1��yY��$��oi!�tT����l�vM�������q0������!U�DJ��Ĭ��V�4����M�SmZuN#�rq�d[�t����	�)TW���"#�M'�42�����p�#C(��@ �|�Dp8�tBs�p�����R\�cV�tu��^����ruBY�k�g� �_�B�����A�G1p>D�P�Ő�UE{$glM�n����d[?A?�����}~"�fgl������A3T��q%֒���GU<�k],�EFc�l�R,>���F��V���Bg�a���Ж���ݍ�.I��2��ol}�#�j�ȷ��������̯�=����+�OL^���������Å�*��ztq��h}B�p��g�7ǧ��N����+S�؟��'3�z�Ù��L�w繄�ɩ�h{vn����b���.�������p�y~tq|������Gj=�x���>����e��S���Oo�<����pNן�T~��������m���"�l�ڋm��Dñ{%��R86y۫u�G��t�Ф8��=�*+�+���t�����
��¯���׎SDA�,?�ӊJ�A�:��B�[�D>p�U>�ЁE���5���#h��M9�j��'Y���4�������xOQT����75�x�����sO]�xx��6<Qg����g��5+BAo|���U+P-��I���Z[|]Ǧ�]��(J
-��!N�J�e�>�қ�P��-�Z��s�&)X�,kW�3"V
�k"��&;��Uzk��������1f�����32 �F�ђ���k:�S �S��t�32ߘEMc��δV���Y?���ղ��\L k�Ȳ-�Cp 6�Ǫ�9�]    IDAT�Dk�>9���*���&���NQ�^��[��0�(��F�M�� ^�U����>R?z�d��C�B6/.4S!U�[��:{�|����R�N#��^r�t G��Q"9���$ҭo��᳢���H���O�����`�~�����du�@�.92�JБ%�lk�)��z��iz(��<�-�X����9,q�o��f���A�[�,|�|�|��L�R���H$�Z���ѺV����w���I�mTB�m�|WZn�(��T�� �E��V��E���B��`�Oֻ6D��(�L]�h���Th�D)ޕ�C�:p��e�@HY�h��	Y �IbD(W������|R��*r� �[g��-�6��[��GAcZ
�� d���dsp�Z%�7�h-p?��V���f	��!B�y��[<)��h����|â"૮ϗDpj�����B���Z�f�"hJ�E�K8�r!#��rER����D�,d�+R{EMG}@|
��W�#.�B�Z�����E���A���*����7ߤ�쟝�&ew���w�I��}@/g��j����*��h�W'�[��olG �\L�f�4SY,5�G�9�QVBc�q�7��M?^���@�H�)�-��%���BX)ۮU���L[W]\�����$;�
��!D�4j�Tdm���oI�pd�ϩ�VW�U���V�ԗ�V�>�1��(4��#W�
ռU�]"�8��p0�K�B�����r[`jY�l�� �mU(t�R��N]`�&3�@ �7jW��h��>�6F
b�����k�T)����n���B-�m�/=K��r|�/9h�[]�q��Uh-�ӟ*�]ِr'J-��G���GfE�q䖞����)�/�(�5�}��(�K���������J���9�i�N��M��R��!F=���N��\A~|���4�8>N [�R���Z5,T�\W9�=�im$�BQS�|jYS�QW,���t�A3��sګyQ�l8��L�8��b!�|�]:!�e��G�#ZW�{&\bW���N��PݚnWEN��3�YC��5(�H����|�)?k��hX���-�_�I/�ռ?'1ٮcuM���B��8�߾A��F_�#����+������k��ڎ'�9)���/�>/�5H��)�i��U�Д�1� +mr#�IYM!x�'l���>�ɢP��hi�����9@��6B|ȤC��{r뭺ղ�p:�*!8DXS�aQ��~RB�J4��s�<��io�'��"S�C��u�v#M95֔�c6M��BÌ3U$V�>�}d�W��(�T4�݆�D��g߮���Bs�L�㓒[!U��B���Qwl�Q**d@�L��:�� �Պi*Qo-vNK�4񧟗� ��uq߆�V����cJ�� @�y��1��\b�ьɦLV���ȓNM��C�:V�C��$k�����#`b��u��R��R�畎�T��R�ܲ����"D͔�~ʁ��s��9s�j[
��,Q���y��OR���|	)��a�j�VW�ZQ�Zq�
A��PJ>�r9M���@���49e��C"��P�i�uQ�V���|W֊���@���'�XM�-�0�n}n�Y��L�%dO�D{@G�� ������kϴ��pM�)�����C� ҏÉ� @ /@пp��s�t�'DO���#ۍ:�ogDuѫ���A�������&�c.�?�i?�/x��E2�k�e�S���m���0OO��֛�G7O���O�;�Ӕ>1�:9Y;����H]���/��^���g3�����漹�9�8�V��|���?8���� �7�t�Osnμ���νcys�W�z���GW����խ*w�Ξ^]{���\�;�}~zt��G�)<?9���z~��*}����w������+������}$����گ��%i���%���Bl������Tt����=]ґ������pWʫ	g�dK�,����D�g N�,) ����� @<����/�b�	0Oz��G����gg&q֠����4����į�I�0Z�@#��`��̞H��)=)�^�]��BC�ogpr9�!���������Ro���?�����UIV��{1�C
ٲt�R�����.ڞ�B��tS@��[Q���=A'n�#ġ�1L"���,�*�'�ͩ:��
d{ԩV�+�V��$P36��s��x�O��,�ӎ�ɒ�P:�����Ti�z6LB�V�@��ǡ$�HL�a����i�dYC�,5>�I�gE��;��Z���ҩ"�.��;�Ď���SC�@�j �6zn�O�,�DK�tQ�m��S����e�b�[.Z�hl��TEY�VQ
_ԉ��z�Ҁd��gKB�#���iBz���8��d�� ��#�^���9�2����`��ڠ�w�A8�R뭰��S]bґ�ï{Y���E��!8Pzʥ�A��@�,:��9FK��5Ҭ��1M�H�q�W�/H�=ut���mEh=�M�78E��	ڽMxuBD���z*ݻ���4�A�� �%���-��HW@���'r0!r�$�2U���셣!��Գ������d[&�D袈��(��כOn����v,q�@N��N$e��}��Z�D���8BJ'S��iVm �tJ�
#`Q)�p),� +Wu�K�-���YӪH�O]�v�>������'^��J'�e"K�aC�Z�P"�>|>>�n�5L��D� gS� )Ē��������M�������n�R��k� �s�h��KJǩ��Y���ت�r��1*�B�9���V[�V!SU��T���������y�QK������TK�-^�O��pC���JkCQ�����m�n�愣�(���5 �(Z][��!A8��a���޴�d��U�k_��������U)e,�)8S�^#�^)-�m�����L������m	��f� �洜��E��������A�f��S6��g�� Z"u]H)J���)���l ��J�������#����R|U�v:i	�N�㲢%"*��F�ժD���l
�Ӳ�Ut������
��0[T�vr�_�L%��l��|��:|���+d Cd�'2d�tp�����ю5�CD�II1�F�M��=$LS�֋P'���9AN�6�M�8U�\�
M
��wA����BՕk:
�բO��M1�U�?�D�SJ�
�U	�|��uX	SNc:��l�J,1�&�[�R��E��%6U����j�#C�ÑszF��,��rR���k��`��"�D�S����,�kM��î�]�Y>ex:��ᕈ �$[
И�1[H�J�uӈ�OǴ�,И����F����K�l4������U,d
g'�O$����(Ŕ��O����4��Z{"��BΟ��L!ӽO�4�Q�oi�b�`������H���p�A���P��DdLU�%������h�� R ���lJ�G4�0+aj7��Ł$R�)+j:�����C��Jq��kҴWYK��V"K'A:�4��DcB|�A?p6ߔ�(�`% }�`"Z�B�h��dCp�z)�F�z�+M*0�%@�a�D Z��F�9BQ!NmEb�oh����5bS�l�F��!�S����1�Щ���#�e~�	�őN�c�$?AVu�j��VL�)y���q�%r��+�(�/�� �����B�S�B�
�PJH��V��
-����KǷ�[/��anZo�!�Y�"R(�~*�`�pS ���E�E٢XY�Ĩg��CR�~ �Ʋ�Z)�094!3��m�ЬM��aQ���L��Yh�g�Á!d�45Q]'8R� ����e��\�^�O~�ڎ�6J!U.���+WE Z[1����1N>�!�_�r��Z�*�D�8������e���7�!~��'�t�˕��� 7M`N�!�`� l9�a�@A�Ѥ��lk��~?���o������Q?lÊT�uJ]�V�6��˽~�sðm/Bk�ma"Ѵ�^s���cE�V��]�\Z�z����3�7�ۡ~�wO���*��j����t�n'O�;x��G7}����ح����IMd�v�ՇǗw�T��ǳ��GϤ,��������k�8�������@��GiZu����hu�ޛ�9̓w%M��|��������c���sJ���p���>�v�Io��^_��k�٭�E/n�����N�w������d�vl��҃��k�V7NS4��������g�H͑�KD3�*ݴ��k��90J�j&A~�hҠ�ّG7h���\��B)���j
��FS֐��[͇�<���8!�t8�j�����K�N�8zFrH��Q�s��> ��_��'5mfkW��xU�������;v�C<�Pѣ'O�=i�4�3�GQ��qڥ.Y8��K��H)
w�Ėo��!��~!��pw���OS9��h��dV��ҥ�pd���P�z��.��C0=[k������կ~U��������~�ͽ��[��чk��LmDbK�5�T��JG(
��O�aQ4�ؽ�F��|)!�����B:���F�*M5@G�-�U��<|[�Z��,�'�VKbj9��S�ZRr FͣU]�n�p����_*�z���B�Œ2]��g����F�ԧN�N��)��G�p�Y.����u��,g�@�/��]�}r������\b�\��<I��F�p��6_�Y@=E�Ka#(o�-YI�R(2��p�V.đU�^��va��lUJ�O��hTN-�d��9��oxA*�	8O�ղ���6��%�o[�}����6P�:�P">�Qu���𡝧3R���w��߶�i��x@��9|SmK'%�#K�2j ���p`w>��rU1�����\8����tg�ᾩnM���x�05�!�+��Y����R �ϱ�D���\�@�]"m qn�+d�����b��iid9t��������D��<�ê�C�PPwR��:߲�_�#�4�����iji��B-�t�A�jF�FM4f:0Y!#�=�p��ZZ�J�~4 W.?h�㣉f᪔X��]d�ڀ��rR��4��@��a�f
R8R���c�OD�t�[��p�X�G���'"��t[]�ƀh^��Meyu|��_V(��8)4eq���F���Cwr���۸�J�(�-�����Ek[�v�����%�K�!�@��}����Y�i����r^�v��{��ZGHiV?^������1�(��*�^�����o�������#Sko)pX��@Q�pL����GF�s�:�7�&_�rӧ �����rz�Ѽ�	5
@�C�_��۩U��0�߾�4j��d}qqA�L�9���0Z���	Q�n�+
�?[ѭ�e9���Im2��Wζ^:����W��E�4������됅狶��h
AP%&���@qL�R�@[�q�"���]�o2�����K��~���S
5�8�J���@d:|N��R�G
�n��F= "��pR�$�2Ĵ�K��%����Bk����^jG4�N.��*!�_.g���n���{�T3��4k�BYI�FG���ȥ�5͟�
���Bl���^�R»�#��+Wd^���~iK�mK�e��!Vg*r��T�_�(���^j:�ǁ�bG���EA�/���n���0����� ��^�������FLxjҫ"��!��ZdE�hr�H�?ue�qD�:���R?�) p�tҤPb�!�������C���LRK��B�iFÙ�R6�-�����@F�T+�-�Z��V�����{���<���!�g� &�o-�U�ZkD�ȶ
N
l"�O05���KӔ�Q4q
��D͔R?|C�(ۀh�H'd�(E�T�\Y�N�8z�7Ф��J!X��p�4<B�����C�)'��OG�P-�_(-�c�_'%�}�XkO*�B�!��D��b�
������r���ޖĬ;���&.���l�;
B���bʙ��^�MS�5�#���I�^'�vCeM�h�!�Jj]�Z�	m:E�Bl������ k�m����!�+�Z�dCh�5ʩ�4!�n�u�
�'���Չܢ��K"@Rpc���B�R�Y��l�H[�'T�}�VE�Yu�A��|k�
����`۵��x�a��!��6eKϑ��GI����4$��%�@G"���[P��ˏ�v��\��A��$5��"qL�M)Β�px=ho�n_:���[�(N��j�Ͳt؏�4�Y!��t߶\���ϸ�u��_�Yԭ������c���Dમ�6�ɗ���b��6����p�S�kf[��w.o�o/L�K�=I?i����׷�O|��B��{���C�>v{z�����������zu��}z��z{��������'g�z����f�|�s�x��p�?���jx{+�ٍ�G�����=O֟����q7G��̧_����Q��Z���l^]���r~z�����n�ϲ�N�'�'�8�>��:i�#�Wٶnە�Ԧ�J�z��U�ܮ��Gh?��bW�o��2���8�p��ԣ!�WM���t*�DJN�"��	�^Y5)�Q��K����4>0��|����j�����rg�6q��*�j�W�B�����T�W�����o��Z�͛�~��iz��)!�mN��=u��,�ه��2�����Q�2�Q@SB�tt�f|�#��GЧ,��?u"װRLS��pT'BV]�����!��Q
�-�(���Ch*dE|d��E"]W6�[*��T���޳c���?��[o���RZ��FEsȚ� s�Y!�!�r���d9�
�,Z"���yq�{_4���&���!zh��v���`��q� r���\ ��(p*�vu�J��0kHhp�c��ȓ�1JaWK3R�V���5��t9亾p醓PQ�t �8;�`x���D�2Y�ΰ��X��'w�`��`=�U�'7��^{ͻ� �z9�����XC(�.�Q+ECD#�i��*��V� �2C�Roր�TʊR��bI����&)���2;EĽ���7�>�d�ݼ;(Y��ѻt.	)�Y^�.��5��Q�r쳗�m�5ٞ�*���&�������O\��ԕ"d
o��ҥ�RD���h}������E[�&u�3XtܤH�w������i|:��MB�":�hV�h��FJ��̶�I��������m�Wd��@��+=�
�X���x�騢���%X:���l[QŊ��1
qڱ�|&ZBJA�>��h#�%��#����jZ��X>Y���"ȭ\)�L:E�9Bm������%" �]M!S�Z�V�4k)��#����ɶ�J��nH���:'R�|�a�K��>&;�Y��͔�Bd�Iq�6�ٍ�/
�^���rY�^ns��3�l>g�5��W��Ѐ+�/Mz5�� �;��Z���* �D�C�ju���{i.:��ۑ*��z� ����p�A���CJ��8v/B|]�h@úuwj���q��ņ���:�o8@��0�9�D�r�tlTN��p�!����Q��-�)����_��tS)��&�_"�i䕶�R p뭴�����m\"A),�lQH����o���` [,<}:�r;TBh�G-��V�u�j.�tmS3�B4)p���߸ks�r"$.
�G��Df�B�4�e�Xx�)_Wv�������I/Q�P�BQ"6�n�
�B�
���2廾��cJa�q�}�t�LG�n�[�4����w��cw�#�u�w���e�/rb#� ��CІd�Nҝ���|#�m(�8)�H�@�Lr�������_��d� Y6�~ֳ���>/�]g��ϒ�6�QK�R���'^3�����OI)s�E)C�7&�t�m/��ьr)��4V�@��2�����N
1`jK}KI�,&�)4��/׸����S~��i8
U¢I�;h�X�ʪ+s�zpL���c*��ьf���@ԭ�)s��q��&��I��"Z��N�ݸ���)e��nF`�N���
q�Sz�zm�P�7%�V��4H0�i�R�$�*�̏/�a@��GK0)�,�p�hH�    IDAT�5Y�1Y�q8�EMۺ�����k�(qBu��:A(��$���D�p�Є���D3j�ǊZ;����o�N#d��C��)c֩�(��YR�B|�����V#�$���S@�}�m��H���I��8�q>&0��v�/�՞�����ڏ1��|��8���l���tcl-��W�t�˩%RL�ľő�2��h|YUƌ܊�t_��\"B��"7��g|�8�3r����1M��v	ζ���T�m��	�f�BmQ
��R���B)���66r!��`
7m���0pT�d�z(dڍw�J�P
�Z�zh�Z N��8�8pp�h��r:�,E(D�>�)�OxWq�h4��������f�V��Ԕ�K7J����ؔ��	�ٱ�hN|Q��� X�č#>��5RpH������!p����O�*�@a���p̖V�X�޴*�!�{�V�k�~kL��1����#�u[�ʵ^���k���28����%+7�t~�H�ק_���:�f9rG�xj�Om�/G���vC4���X�Q�BY{|;����O_?4'�T>�6*h7D��B)E��[?��ZW��]n���`
���!��g�s���~������'W��ׯ�޴րǥ��~{��p�g����}{��K/�ţ��y�=�Ǉo��}��{٫�{gWVޝ}����痫;o'.�Շ�N��ݸ�n��)�΁[��������/�=<>?��O~�7*�8�߻�|<�w�ׯ���]����mߜW���/=}�p�C���n祏��p���Q�Ǿut������f��_e�Q.2��Fx�1%�� 9�8��3�#&G�(j���W{o��N�7p����$}̺�s&Ħ�i�S���Vnd�F� ���^��q�P�12�1��FyS=m2���e�,�/�Ԏ9RIy�����wo�t�*�i�K���]��oW5��=(77�C�:
j�H{�Z������B���!��uA�y+��%�%>GԝP�y�L���1Ug��UQ	Ȩ��Ȥ�U������,о���Z"|m`:�TD.jD��!�������������˗���6]d4q*���Y)�q�1Ӗ/+�GЌh��T�*�I����������&����'��@�����E�2E�![��$.�t>�= y�k�%�"©�U;f�S�N���[�Z��$�lJPtV́���Q���:Aj@7"�"z�˴]8Bp>����h��r2;�<]r���7��g\/?ݬ'�-u�#*b����ȟ�#K����_USKJ_V]B�ȟ�͋�DEiF����-���rC��5�sb4��=�C80e��V�)�ur��b���R4�����	:6�U��ގ���.G!��j8���O �Kݢ�%��=��!�)S�zei��ҔY�Dp��0��BL�4�J�$�a���_cn�����x�믿�	���=�9@確V�N�ҕ�-�uU�V�Jג&� �Գ(D�ě
)��H	��=��`6�F��t;/j��)P"Cc�dZ-"� ķ?F��ߘoDh����q��$ߛ���7�0Y��);	3�ו�&\�*F��Z ���Ь��l��u+�V��N�S+A ߈	�0"F!�ӛt8�m��]�`�֭im4m���3}S8GX3�j�b�5�Q=���%Ą��|�3J��>�L諯��
�wfV���퉦S1�S����oC��FáO��?k��3�B�_W�]�I��r,M�����bt�M��ݍ��DMR��Vz��XH��v&��*���Y�,!B���6Ǚ�~ך; �?As?Q��-��(���TrEݬ(�;�+�o���?�Z&��F4:|c��IS��u�F�tc6|ç
�"PzwrQS�k�0:4��,�%%�̽"ķKv������JKp�II�H��3!�A�X���G-S4>G���C�C/W���S�2_b�Q�"�T^�S`m����b�����!Dt��8��66=W�X���Cm��I�����M �(�$�rS>C0B��M�\�B��;�V�:.�v��Yf�+N���q8�"axS�D�u^zjBY�|����rȦi*��i5?SLS��D�k�ފR��扄��V��d��C8�CM�i@�N"'�_)L�T�|"G���%<�}{Ջ"N��5&[(�	M���k58��[��M�W-3m�FR�}!
���`4SN�R��C8+�+N=��gB�4��C}�;"98M�t�E�D���f��s�6��]-���[�,'�@���SQ�(��s�rf�>C�srk���4cD�?�!q�ZqV�@���|ʍ�1�Ӵr@:%Rk���&�Vp:qV�鄦n�!�kLJ:iN!S)BR
���NS��|�SBJp҉YKRF6�*�*0��)�]�������CR��6�*����M�5˧��U�>��.���H�ҍ���t�I��@S�`{�Z��K�Sۣ&��f�|:����'�m���0>�zh9�־:ێx��L��<Y��t��g�P �C��J�(�O���n�pLS�\`1
�pL�%;�@
,<ߘB���$�S�a��:�f�["�i[�������,>��)��B���B**SW���H'[	#3�a��B�-�ɏ��1�+BY
\�ٓV�>'?&B~��V���ȟ�r����@Әu��~��CX��7:�L�J�>+g���I��Ԟ �D��S��eD*W��TH��U�@Q-d�t�r�L4A�~��WT����X�4�n���@Q�����eCTqoT�*�!	VK����ȶ�
��%h$e��hL�#Q�\c�PQH�SES�������d5��B�Ζ�6��N��roNz��_��F̉�G3�l���*�]^��j����R�h���n��k�p��Lg�ù3���:������yr�l}�����XϮ�+�@�����/��yK�0��t�?���u�Ӯ���u|}|s�/Zj��)��G�8�r��z���t��\�5�"���� �����u:�t�󠾊�n=}�v���gw7�W���������}�������g3=�����⛳����Oa��~�����?��Wv�������UOV�"��l���^�عY�Vhm�6��!�6c����aj��Ԃ;XF4:�R�w�`��8����_-�d~��_}���W�V���)pp�5�~:�BKz��g	�
Q�ws��\�d�0ǔ`)F~S�Pˏ^�p����)�N4!�F�f���/���CMo����3�nv��˗�!PFn�P�@"R�	!�I��v@���.^�@�h4M�7��VH��b��)��j "���s��Q6B��WB{�G�`�A��|jLiQ>��p�q�ސ�����'�e{:���+oZ�BZ|!R	FS�2���hQ-�B�eM'���!��ؐ��D�g�L�V�TW(N�Aé����dҤP���WG�5�RQ�vIB��X4�4�(�)��S�i`|��E�E��:�k�	ԏ��Υ�:�h,�)Y�L���V��g�RR�YU���)Aә���p�z��������2RF�9���q���Ժ���~桦|*D�2�mkﰍ�v8�E#b�X����D+���
���u,�IDC�0H��
��#Qtʅ�B�-����$+ݙgJ��h�A�}F[d��AV¡�;3��t}z_^�s��>�d�fK�����+_��[�T�A�(ALo�z�^9��W��(��G4mw��n��8�Y����F�̞��r�0���?�X��h��[]!��)�ܙC|LTcN2�_�dI�B}r�df���f�2��ŗ�r4�%`��1�~*T->�h��wD�Z�DpR��2|�Bd@N4L�:7��X/_���b��~��ҍڞtQ���)��40-+f�П)��A�f��q*r&��D�2!�(��O!��������5�T��S�ЙS�FRE'Դf�n�M4�hFS4U�?<�
A�͙r�(dL�[ q�?A���r-����H�6dg5��D"�QQ4#��B��L�%��xIGE}�*5wL��ݦZ����媎!峞��y��;�7"8q�)�J�S�����BQ`OR[)|ZݷͯQ�fJ��~+�>�yM"�]��K9�
|=eU�,=K�7�Mm�5B��?�_��_���K`"��B�e�ג��Ѧ�`��̷�6_�����W� \�h��irl��i�0��`��a�N�쿭�"��%@lN�F��6%��P�Cb4m��K_iL��<����[{8&�4�c
Ĥ��A2�C�|
.)�B���D�&�,S�_�8�|�:�Z;?�@���͸6+$Q
��Kwkf��a#ܸW(]���&($=�:��;���D�3j�5�,�f�7VK��@"9����{29�R��fB��f日[xʜd�4e���V����g:��,+d�9��%.}�%�$�RNNJ�(��0�r�Z;@?B��k[����GJ#)�(�iJ�ͩ�c�IS?�xj��چ��l94�m��	�/��V���_4�j�2�����
B�Y&5f
��0Sh94!F �qX���	"�YEYā�@V�|�����YE�sU��":
Ɋ2J�սce��9��Zk���H�4�"���UԈ�_����ъ�"8�1�rRj^o�,��Q��7��&]���J+Tƪc*7ܘ�HY���Px#|L��s�B-P���Q�_J��SJ�4�N��6�V�O������zS:@���Y��V��z}��D����Xq��U��
��J�֧�N�QP�����)��p���5r�!"X���<�M��� ~�,�U���
�0�q�F������	L*��/�1ZZ:!���PQ׳i]�&��E��'��|N��~�tL��0x�F��B!���+�F�C�2eh��J�i�S���>k��ƙ*@��;F|�v��.���s,4�ǨU/a9�! E;^�mLS�����`���l��!j�ǑŁ��hBx�&���Ak�$�)ʧ� ��&9q�c+1���lvRKe	�o�5��12�κ������5J���d��l������%"$ר#5�G�i�֓��}���ı	B91)W�-EpR9�*-�&���!���OS"����j��B��^Ti�@u9u��at�2�{BH�ᦺ�^�j��P���QK9���	�-5�+�� t�����c�k�Y�ۘOo,:��!:>>�A���6�ڧ��K�:���v;O������W���������w�GO(�^�Ϯξ�{�3ή|u����������v}w�����o�a��>�J&�#�����R'�,=�?^�?�9�n4N%�V���ί/��7f��~���9���;}�0�����OW="]'�w .��x�k����p����pyuy�m}+.g=sݎ��ky6mB�d{��ӭ�~
�;�8�:�f��t8��v@��ؽ����A�Q�7tLo��ՃFo x�ٙ?�jC�֤��e�و�n��0��_�3G�&�oL���0+4U8�9���)�a�,į�qR8k�L0�:+��o�w�w��ޝA	��r{���n���(Ѧu3�(�{Y|�Lg��Y���:#�:��+d��,F�ˍ2�P��������t]Y���Vu>3U+���r�:�wϑ2U8@�4�8�+�^:��m��W�)E�Q(�6��@�vO�[?���L'�p�n�������H��i4����1��4�/n��)e+5ZZ�����|4�ݭ["�����W�<��Y�Kq�8�;�@�8DƧ)}�o�	�OJG�fZ�!�wb��BcQ�t�a8��B�1�.�fΥ8������M��`Y]&��Q`p�l�=d��9�.=��Yvܨb*VH�+l]�����ej� :i�B|�̴� �~{Z	 �c)��SU�����N�0m�
���F)�$r��u�T��FO�����j �MD �
ۧ�)���a��M�p�"m���:p�3����.f���]�k*�����@�ZUD�h��!G`�p|��0!�kF.D���z[��\��r��͛����$������[��>D����|MJ�@�w�H�ꫯ�N`��(���tR:�D��q �i��4��ƌ'�9uR4��������r�FNU
A�&��; �څ��O�Z��yS��aJg��Y������Y(�?�,��±9���3�B,�}Q8�I���.����p�o�+�r8pS8�)��7�S���X�� Ae�8#�ACH�3�l�W��&�pȞ�{�����f3��Y�嘺�\).���NZ|���w�Kį1���� ���UD
5�T�� 5�[�F%|���#7-I����$��Զ�F��X�K���^
^� �TM��Rr�1��$����[g|:�����dn~FT�]��=!����8��~2@�kRK�Z,���H���zp�q�α.)����BZ]#��Шn��X�JK4�O�TEdf�	�(�)��C-�#AU:XB�*�J��K!?�|��V�'bRCVB?@�>�H�ǔ��p��iN�I� ��eiH�Z�׶#e!�D�Ap(!,M#YS
�oZK�ş\=0S�8,�p`�U��p�h9���ӟ�\f[4�4&'�#�ȒfU�Q�������4����%)�L����c4Gʖ��,�Ītp�hR��új���H��V����{��"p��5���G|��,�~�p�"���q�5���hU����7&���7mT�u��B��"�T�h:=����α���	���˯7cV:��t>S�HJz��Ulk�!e~;0��!5"˘Ig���X#�MS��I���l)ш��qR��9C��,���_���ӭI��e���N
��R!c8ߘSW�@�A�+�9I �Y|N�@HөX�Բ�O!5�@#D��2�p
�uEV��ɚ���R'�O
�HQ��ˉ\��BָouR�.Y�|�3e�Y�U��X@�����ۃL���=dۊV�A�� Ь�F8B̚Q%ZN����#��@��u X�t�_H.D��ܑMA(��
�[>�B�n�Fd:��ǜ�V��ӎ8#MN���,c&*=�nVp ������J)ڢ�J� �3�^#ܨg�B"p��?{bZ����>f��49p�t��~�0��g;	�d9���H���ٙV!��D@3e���$�щ�����cJSKz3�T`��݁;�(.�hʄL�[�r@Sx}�|���Ye�R�#�%H�	�D����ڠ� DHucj|~)U�s���s��n�+����TOA��4~mU�]B����T�q��T��Bf�ï:�M��!�I_��d%��|�����cDvL�+ĉl�i��Tk1F3�G��ïB�t�oy���1���F6�*j�uնh{k�t�7J�O��th"U�n��9�d�%V���8.cuG$��LSQLLjFRF����P�HM
�RK�,�ۓ~�������{���EI��1/=0T����峳O���}{�9u�LVn�]�V���⹵;f�I�T��g:�N��_�7��-i�����G�4������̃�C^�����+a}i���;���å���0|Tҷ����̋�[���?�?��__�1�9�|��X��.
��������z^z��݃�ڃԇ���?���?=\��?A��=�����{vx|x����[_���4�o٥cϝ�߁{<����Þ��ۣ�y�y�;��"�)�!��d���9�m�ڙ�,���9�F�S��Qz'�È�� t#Ļ
�c�m�B�_��x��{��#�y%DA�%8�����aN1����`X
D'|��o���ń�!pdc
]��f���,w���k�Ȅ��z/�o��o�dM�F��]���sGvI�+����s��C�;3ރ�Ɣf |�"��"u�G�r���j�\{޶K�8�ٶ0E�p���CĢK�T"�N�� �?<�U��<&�4~[A�'X-!��A=� �Ҟ$BfԆ�#���,��c; ��s�=9���ݞ���u�XK���ۚN�@d��9B�+&dRpDC�h��Kw�!��b��QԞ�L6ܸ��A���y!�3E�8�샷O%�(���!�Ҵ�2EN������N�̆    IDAT�ӑ�V�4r=1>C*����_S�c��"3S�oqh� 
��Nr�� �I~d���&�)d�`�����'�}j��"��'�\zP�$�!����:��8�.S�b��U<��!*���q��f�U�(�r4G>U�ȖJ�a*1�Q5
�pJ��e�@L7%k��q��
S8A��pw}J�G(��,�\��
�x���|�����8.r�d�`�$��~�uE:��uQ���5 _c�R���E���\�**�Z�r�`��(d=PA��۝�q�r�A�裏�"�\�k�,�49^#-���Q`�rm]Y������~����k�k��)WWJ=��!�GQF->?�>��R­�N����T�
�(�Ԥ��T�)2���pӘ�54������
��EÍ��m��F����h�
Sc:�m_�(���E�I�'1g��1ud�7�dҍt�����%�ȢnjK��n 
G��8F:B��ɬ��TH���)7_.�`䏓Ό���tJ)B�M�� ��@���BW�u�Tw]��0e@�L&Ő�N��|SE]8�p��ݻ<$��N���:~�	Rs/�\J��`hnqR�*�r�Mqtkʑ�c�'cw-7Iw	u��[Ѿ%����3r)4��SW��_�c*�c3]�/�zce�%˸ֹ}��ZR�.��)����[�#N�5nz���r������)�j����)�1Ҥ A����*D�j�2L4�G�إ�,��]�q�)���1Z/GcF:� v�SWm��(�t����+�p�,���I�D[�h��,W��[�I�B� ��F��83Ն)ˁSH
�����F�Rn�����v��"��J��DƇ���.���X�8�*��,�D[~˩����DY3���R�P-M-Rd�ꮞ��m��Q��)~LȨ�ω�\�>q�
%�QKBY�=��2NK8SK������"FW���a�D�����E�"wđ�ؙ�,D{hEe�ib�c����.x�|&�h
Oܘ��š�g#Cn9�D���S�7�Ñ������-�~8B[�����c����8�S�*hI��*VK���+��V�h�����m��\o�Т����岖�o�OJ�7��B�d[�~�F!٪�3����D|�IAK�S���^��ß(0�(��b�A�爖�B��|Y�OG_N30Y����M��eb:Y�� Gb#��c�Ԅ8c��FL`|�h-��S�4Ίd�r�ƒ2M��
Xoei�>���J�4�"��]і\�i�T
f#���.?A�D�P.\��e����&�-
�?#T��ǡ�g[Q��A�N��� Y��c1#�jO�g�"�A6���W�)MG*�ic�Mu�|"8U�7��S>�)�S�1�F:,�B��)�-�����{Eq�!Yp�7�36���۬�U�3S���'.���h#��a:mE�ZK���s"�Iʔ��d�i��D	іY
p���%5�u"��,�hcY�� �Q��q�!��K�M�����Y��?C��*���r�ۊ�pի��T�#U��i����L�Eqʆ_n+m��,#f�D�f�M=���Ԕn����rR�LE��B�d�Y6��
�ѯ4D��'*���ep��5� Џ��2
y��ȷ:"z0�2]��&Hӯi~��k�]�~��I���^��?�`�:O~]�6ӓG�<��� 3@̿�C��K���^�������k�'C['�E��t�z}%,�����9^��W_��kc���W+��g��<�shݟV���˃�O����kn����n}�������o����w69��G#������=���xv�ͱ�M��,�g���;�������K�����gZ��g�ח@�������G���㾹{�އ|���o��H����\�w��������P�}��5�Oض��ַ6�ήh��p�̣��l��Vܺ�h÷�\�+ˑ2Ev(�;�k��̥w�K�s�CT:3�� K-Hךh���1��:��;0�^���\-#�C+��7���)��Í�'k�D�
�t.�Ԉ����h���B)H)˨V7lMC�	rjÔZ��{_�����k��-�nx���?�������W@�>���t}j�m���V�|����p-KA��>�,�S!��!38�����$d*Y����2�R"��4Iq,�i��M�0��)�8�;4���9��q��95��硔iF��$Z�,F�HV��Ĕ������)Cۏ�c�@���b���rK�[u!H�"'���Q*�[N牬z��\��	K}�x[_:��85�Hꈌ��Ud|�F�7
�"3�Q�STcD�P��>��������"K�[#C���O��K��)w�M����Yv� G����>_/��x4U�Z�O/����>��3/�P���������ը]��"�JM�1���#t�R[F�)p�|��t:�����Z�M)pd�5��a�Ub|�ҫ5S!���0S�:.`�pU ��>��m��n���������E�)}S�J8ޯwr{&��C��M�U�N%͈�?�0�R��	�+*d��@�m{�����ws'B-��Y��8���(��MJ-V�[�g���4�E�[o��ՕC ��_YHn=��!q�ҳȲ�/�Z%J�@�|N���3�i4�60����@��[40�i�5C�Q(�ijd��98ՍP�m�)�)�H_:g��.ISR����,TQ
Ä`jRV�zHt	�J��X��P�&��V	�3��d�@��}::+�-gV�Pz�Պ�h�F
3%�~Yu^]c����4�m�=��u	{��8��D��QM�M����h.F�-�u7�� �
��_4m�B�
�z�cR|��(���QTVk4��u"�6L�ء(�����A샢�4!:i$e�D�8�ԝ%Ь������r���ʕ�z�1%*�f�F�?���O��-�t���3��-�'ejdc�V]9��L��ɢ���QWm5������\��r�1�B�m��,������{����V$�r��jY�,F�2��`��r� >Mc/d4���_�>���6
@֒��Od8�68��ɇ�)�����01[~)e�UW4�ꥋf��pc 9e��1Y��̏�1�D�n�4P����B853jÙe�)Q��K1���ҍ�aD�>���Ѵ&�:��N���(�%e�?��ᢦZ�O�b]�r�Icd�\8������BLc�*����v>Ǆ3�.��r'dʧC�Q�@#58�E��g՛���Sho��*0��E9�Ig���)�5%���l�ۊBY8�#�K�8�zf������iR����3U�S3D���Y:��V�K�i) ԛqIo��N��:�E(�ۃ�%E�pD����B���B�J� dʯ�,5!)�U�R�3x��z{W�U�Im���:i�q(S��1��:!B*
�^n�;�h����Y�nx��)d��9�1��9eqll��j��
�Q�L3���hG�Ծ�z�:�hk�*F8fc��>!�j�S����mE5�߈ً�t��H���id�������8rY�қ�r�wJ�5Ƒª�)���)�\9�h��0��δ'%B
��\
�u���zU��HфgE�:��a����Yd>���X��v��Uy^S��\�HL�(�4���s|�LG�t�r�[��+}��!�f�PLj|jFV���4�:4֛�(*%f�@�19�"BE�)��qZ���-2N��Vn�JDJuW�m��!m���%�ҪMY"�)H��l]�8�7�!�dr��T4�,4��t��+g[鞆��|�1!��}� ��dU�����*Ȇ�&�Ӡ>�e��84Y�r�Ԍ�K,�)����rj�B)��$�G0m�&4M����+W��������O�w������N����"���Q�B�RaM�2�᭱1Z��pzY�p~�iT��n8��wI:p�3�o�d�͗�7��z���af�R�N�>���G��M��+蓎���Z�q�`�?�Ϙ����}du��y�u����#���*��sO.}*�#?�&�<Y�I��KƤyx��������8����;�G������ʣ���W���*:7�^�����󋃿��6|����I����g�q�'&=����(������z=h\O^��켴X׻v7w�]9aϟ]_y�����c���{����<{~�C�v�C�;����7���on��By~{ュ��C��� 
=9��w��K�n�i��A�]ߡ�;��U,�F��s;M;.��`���Ҧ�iF�8��)kl�i�IЈߨ2Y'���D5糩S�իW?��O;�|; A防8�����ɟ1f=���
A'5�:�d����*�<��)�r|�;R�8΄ԌU:
�H�=����/������������?vM�O��w1�p�*d�M;Rm��2���Q�r���H�|{�����]�8��(�O��F�#�9�d��!�)������a��IG`�z_�N���P�����1��_}0L���[L>��'�<�tz���O����6��~�2�3NQEY�էi�8e%(](�)C��r���>�ȍ@46R�V�4t��Ȣ�&5Y���?m�3:�8���DM��)5V?�g��BD�F
S�	���d��h��D�O��a��j�pƏ��L�r��X	W�WC�Vʄ�=��7uڼ|�ҵl�c���_�x��5���&����Ŷrx��g��VahFS�Qa隳}�Ԗ�@Gnc���~�8<P��Я��� G���B�8�ʪCS�>�Ș��%wu���-�`�86��F��nB<��p�{��i5MMg����vH�=��ޱ���F\�ޣ7uhu.�yd�S�B�Ɨ��Ck��h����u	Y��Qo���=�v2P�nW����D��[�>�ˬ�5����Ok�Wnm���4�O����0�E9��!%�C(�4�)a�eM��MyШfJ�B"�#)#k�K�Ʃ.bZoȦ�B��	�ܦ<�jchBL:�#�U��x�Kn��r�Զ~R�Ą�s�ȫ�V�HG4�z36E�B!5>�VK3)>'>�)�IA6v'��G�����[�p`����s!>�pF�S!Q��C�(B�jE	�3�9�P_���%2|S���J��(##bբB�k�g�)�����j`^�}!�,���O�(�i�b���]}��u���pנ����<���	1�rvC���md	�j]F
�j�ӊ�P&0喀&����v'���P��v4�L�\��@��럨r���7�Gm�;-�j!&�x!S4�H2� lO"�M���S�� [�ж��Z6��Ey����C�:o��D?5[�<�c�'Uz[gJ_ifs�Y}��)�Ȓ�H���bBf�ȭS-��k���g#������S�����t�e6V(�Iߊ�,ʵ�\t��c@
8�Yь8�pV�pQL&j
��B��p�������q�*�Ak���٧�:.t��z �:��7�kD�oJ3��:��;��-��Ky�,)FV�Y�D-q�[�i��)�U�*��-�Mp9t�R���'bL���Vׅ�i�~}65VŘ�N{b�V�	O?�äc��T!E���ɟ!�p�i�)Z��'5@��'�N �{�4Fj�ʏϯ���@c�io��D�2S#��XM�Z
���TŴ����j,XWƜ���3�8{�r	�b��1��D!�(Y�M~|&�Yz�_��ni�҅ʒ�x�[B��SK���p>}����N�ش;*�5
%RB��2�\#�d]GS�D�$(3��R3�&�(������Y��p�B�SuY	�L'7���6J��h�/q�J��A�J�R8� Μ�^m'>mW�4DȞ�1�@�T�ϙJ�)E���ӹZ�� ���Ɉ@���V=��IL��@Y�!1�� �)SPH��E:�'�Qz��p6�U�7�ql�( �D9�9{�ߊҬD�YY>�נr!�� !��M�I���8B,ǘ�(A8'�cKK�Xt*�a�XR#��bL�èK12Sj{pڃ3���,�X(�i>\���h���18�(���Ϗ�ش�G3��X"�L��ܕ���G+eӞ(��@�L3��J��Ư��B!h�3-�Z�3�L����n{��,��8�:��j�����OaDҟPSY�v�� B�M;
B_�D�r�]浵_��j�/h����LѪP���#���B$�h�,���HĔ3 d:�[��D���Ƿ�
�j�Fw������4�`Z,�~
��8팩^� �*�M����RΠ�B�ͷ��������6��[�1Moy:��â��Z��1�s���uB�]y�����[7Y�3�\����̇�g�����l�1O��mo��;s�T�{�Ʊ��6ϯ�/�=��;�����:��.�O!�����ª<Y��D�.�����-���O�s�n:J�f�~�&ᷯ��o|������ӟ������+h�oo�|���}�powgW�!�.^�E^<z��z�ݫ�=	��ѳOߓ��/��|8�����uw�QL|�ϱ��yE�t�������O���Z��}L�i��h�l���t?DP�q���~��۽�O~��Z�����ʉ�j��U>fVW�p����Z|�ҁ���֋��vZ�P��|����F4��l㞆�r��0s��z�������J��o�jѻ%�$��ݠ������p�|�}S�K�q�K�̔S�!�~��>����ar��t8L�"�Î��z��B��2)� �/K3�<�'� �a�N�D���V
I�Q��8��4���)�Z]�1|� }W�;�'��e�~=�PVNn��9Bc�uB
�A�c���F��ƌ�  �|G�VqD�C�)��Y��4K1�m�B��UN��tѪ�������Yf#G��4�ld������:\�-�$��E-�V�c����A�)��Ĉ�4"p\�&:����E�!���А��/^�p
�NDd�y�����,9x.�v��@<Ʉ�����5M=_���AQ���4�������S�n��W&��b.�ʹW9!@�J�N'�٠�b�
��fL��fs�Jf�\-�zD��'�t�ٺXK�8r~��f��ʖr|�����A�����)D٣G?���4�N8xV���q=E���N�h���l��%�D!�~��h���>�����?��Ok�����욤�����U4���0!̎fP�!@#}����0��<�DY��Q:�Z�=4�hF"�b�1њ�G�>���@��F�,���W�-M8C�3%�
@�Z���	1e��Zܸt��}c�,�i]�/�i7L�^┈�;
ȶB?�4�F�`���c���)�qY�~-q��#^�Z��9-'��M�%���P��Ȧ&e�:��DngD9�Y�M0
i�~g2�BB��@�R�r8h̏D!��\�RH{kD�,ъ�Y�rۚ��^�1��\�����t�PH	"F�Z�-�*$�6LC����_��,�ïCS�*�����E�)-�ٿ��*��$�)Dp��3���#�h��&[�J�Lu��B!�b�M�Ѵ�C��8Lȡ�(GJu���I���)�9�F+U���X�%A6"����FH��19 �Ǌth*��/`�:"]3�:��ҵ�tU�ܘ|d銚S3�z�D����!I�["����/ݔ%˙�Z�H�BdȢ@S�I!��kʁ��#4�r��DD��1�y�F���m�";'g'b&.���FLcUptX���VJ���r uX�X���L�:	42�D?�ڮ�v�?:��q8�(LN���`2N]��@L�UȔ��ʁ�3�)�t-ďS�w�J�d�r�U]`��)?��%Q	)RM��G���B���Ut��}3��խ\�e����hB��i�f�%��F�t��0!|8UȊJdpSQӭ��rj�1�O�O���K��!t�r�DgZ��Pu�(��Q�9J^K��Yѩ.RtX�z�[��{,�M{#.k��c�Aފ�N `)��h��D��Q�8B암�!M��G�#ʺ�Y�;?2�9,��5¯�()FX�M1�
ͱ�.����s�[NL)�S	H%���D�\�ӵ�    IDAT!'�O\��42S� �r$ꍯ���K�\.�I��ͯ�(�o�#%���'� YH����ߩ�)�Ao@W�KhJ��$Y��6�6B0��ސEьl�Ŭ�ʉ�tj&�|���	��^�/�f�:�4��s��r�1��Ʒ����:["�1��o�CR+Zx��9�̚��ƺ���1F�
�E�B?�	������"j���Sb�[����0���8�6m���D��>N��IY;����:�����O�Ȋr�9)�@H#�N�G�H-0f"᥏rSR9F&��B�=�����k���i�ڌN��8�7FH������q��SJc�Q"Ę��O�"�Yې��*L�F4�%[�@S+����@Rn�V'B��z��~�{���t_�Z����1MJT�Dh�
.�)�:�v�_9�jR�U1e��ތ~�22��� h@��"E�hJM:2A#��n���z����P��v����b�ضW��%��NSQR�1����_n�uk������O���J�S?�����W�.L���#۰E�m���u���{�6Ҧ�� ��Q��0��	��a=w�d�}P��sW��gw��z�^:P��R�Z�Yd׌�7>!��eZ����;��ֽ�]���4�e�^����~��������y���o�'�������ǜ�|�훣��g���[?����}Թ5��[?�]\�=������G�~�Xo����t�1���l��;Rֵ%��������#4�[Ǧc��0d?���������Y��o �˶y��su�!H���t�qL�2�;�n8C�V�,$�����9S=Pz���>ʩt���蛶K������͢����
��N]V��m�����U~�*M;..@��
�j�|�{E�_�Rh|V�Z�S|S4�m4�|)��'���8r�D9o��%�*mG6�d�9�z��g��#��eJ�z�Q� Wz+�~�2��[�=����7�ޣ%|Q��W��M�=:U���-���P�l���ɟ��er��DW�mK[�S!Nfʡo���P���i
7�v^z���,]{�CsK:��fݢ9彔(k�rE��F�Dd�8u%��
)�5�R�(�Np��Z��>$\--�%�d|j9@:��"v��|pn�G9�M#;s�d7��9ne��7-e���Z	�3a%�!��F��T�)2`M�8���JT	�֍� ��jCkє ��DKG�T!�6n�^R��r��b�M��Cj�f�>2����(��*�yl��?r��J|����:|��ji� ˗�1B(x§\��;)M�v��6꣏>�nLn��/�%�'R�s#PZ�V�1��t�e­:S]���|��_c�ݝ�3`����#}Ul�TZ'�@���W0NV�UD֡%�DD��i-&��'�LI���z���!puk,�S�1��P
?)c��MqX�KS�/�Ab6�s"ė;|C�b)#>
8Rp�j�옕�1 �P�|N��&$�4_(H�Ƣ|
B8I�_E�L�=�.G}>�,�*�3�V'J�N��F�z6|Qd-ߘq~��Q8UdՆQW��-J�er�U~�4M���3����b�&=P��_	>>���9�
ĨNd��hQ���	�a*˔qj�J9�
�X!)hݥ9D��4�)��\�ȔK�݃�2�@���.WźݗF"�����(0�,>�,�h�,d���y�6����己Rl��l�cD���EVQ�O��� ��h�ESK{!@���49�
�Ռ�%��8�i���m�pQ��҄��ߋ��ƷWt��!mi�(dJ�A���u��>�h��t/
9�Z�wR���}��o]:�7�ޢ8�LQcd��&UTϭ��ȦJ���R6��)Y�1�4S����f:ȜLT]K�8"e���������5\"��RL�	ր)Y�j�ަ�e8%�lsb!B2LƩ���zÄ�!�c��/7�B!��e��B8������09l+a��'"�>��!Ȫ
�S��p`��0�|�g�Md>'�)5�pN8��`��8C@�%r�^(5c�LN���( Hge����!�lKz��!�7R��8���1
��ɗhԆ�U�>�뼵$�7��Pz��
��Y&�8���zP1+�ɄL���6�X?��!S�)��e��D�&#� !�Ʃb�sϗNs�8�~�r��O|��Ɠ��Q}R�D�ًO�N*R�:I�,�%�!��!���C�~R�{e��&L�Fe�ِ���X�*"�'iʁ�s�&�	��i9�Ҫe�8�ĕ�c�i�4�<?�&���o�D�!����*�"��q�|���_����KE�4őX�1�-����jt8D��@c��W2Յ�E�]ʥ�T�(����

�n)�d#�J�&%+E	4)S�C$��N|S�F)�+�B��LgQ*�T�Jl*]�t��V�2�n�ۄn�@)u��'��J���!�No��ڧ�dj/)#+�/���" �2Ȑ���[r[�iDh�t���9B�R�K�RW}~���b�jM��G
�ꎦ��!�1�	�7��\�*���J�B`���L����Q7�JA ��N&QT���ÁԘh�YQxʍ�׈��<7UW�~!%Br�3���)@��hHY��X�K��Z�V�t��KG���G�#B{|�e�F)�R:�h����@�S�3{���{g�믿v��V���չ��P��@�
☊��p�^ɮ���)8�41�)�r�7�|��_-|Y�6�U� ��F?���N�ۆ~�M\-
�EӔ��D��}��ѧ��<���DȾ8u���j&�V(
_�mܘ���j�MC���ˮ�M��ڑqX�^�y�Ǚ>y�]W���i�cM;�<+<;?<�������s�{�8�[of�o�Y��Zwi�բ�icU<U��_��>��K��g��g��=W������?����(��}�o��&�����o|���a�����g4�g��7g�ǋ�3~/?[�o��aы��w���ח>.}�ՖZi7s]�m���wt�u��#�/��_{����+�a�w:�~��ر�LDȏy��Ӗ͸O�it6D+=���AL#��L��y�I�P.�.rm���Ý��������*!�1峉"�Y�J��~���_|�"���~�m�6�/$�_��N�B��V'���D��@o�� ��T!LY��S��a��m�Y�hʽ�b�����f�]BZ��`�eǚ߹�q�i��J!�MJ'��s$&�tE�A�E��$v@!�D��!��� �M��f$:=��/���O8�1A�%�� �Z����9�T�r#s��Y�����L�s|�V־J)��b�Y�XF'��%6S�(�o�)d*�~"��~R@��W�Ԉ�w\�F��TqR0K���bJ�0]�1Jtd�+�Ӂ����,`�s4`Z����3��1�^�y��y3�����=�� ��Z��Z�-�7����ގ:�Ŵ���"��UEn�8�eiEߑ�-_h�F>>k�-OH�02� �!7ny�ZR`u.�C�����U��V���QE{��Z��r"TZ.~�#�[�Y����8ӿB�g���8�D5S?�9�u"�?p�#���0;	�Ч��)$~]�7Ꜧ��t�m�Q��@��!��//������;���w1*�P�B�j�g�MS ���2���[&DԴm4MӘ���h��75��&� �����B�����B0B*��1��Uc����ۜ	R�+7=�8��|Y�L�MN"�/�O�tQ�)����[���ګ� ~6�`�y�,���b�15eR�������p��n׳P�s��c}�T1~ʥ�M��l�V,c��yb$�,#2�L!H�I���ܴ����dJYnU\;��VWSԅ��[)�T����� Wz?H)ǈ�R��6��Ȋ��CHE&�5�S��������G����xUeV������@���_�/�B<!��_��a�m����ߜ���R����9bĈ�s�̪�쬢�
�������c��M���-U	��D��ґ�������C���y&Y%��8������Ψ�P�T��p)x)�%��JM�洗�3���R95|&�-	�rK�Q��Ğ䙭a�q��K�H)����^p&Fֈ��gKq�������Z"�IG��[6Ij�0)#��7���p���/��D7�%��D�-)�9�-����i��B�C�l��"R��"�-�ޙ+a��/�8�ҴԔ����[,U����!�(�&�/NmW�=�KA,C��RI�XА��1rx���)��SL�%H� A�'��b
"ol����"p
���j�puڳ�����ё���n�e
��3��8e�(�D������FJI�h�t��X���D��Ij���`��b�pˉ�������2�t|i`����=����JP�)� 1�'^`MW��זek�7����#+E�C�/n����J�-f-�B�SG�������u���L#`
�ȫ�]9���N&�� Y���u�l�b_;��0�3�l�xK6K%���r��l%���YKAj�8�Jo/˪����_�dw��v�ҙ�,1�A*AA"<$�Q����DHD��	X9D�մ���9�d�� :&��p�o᧧��DS��Ӣ�����3Lʉ`�N
Jpd!,) KG UL$Nd���#�.��qʑS�ES'ͮB�
��	NV��zՈ�E�*畳t�R�W���̀&+U�Q�S�Q�=�p�7<�%O���7� H:�x8WՎ�Z��"�3��
����nZ�I����/���SG�Qkȶ��U��e"|�<�.@&&S\G�)�������ډqx8Y�}A����H3`*iq�/�38�c�C�D3!�lj�/�B���gʆ��W(�q,��`)Ț'}�Z(70���h��W"�6wQ"8��M�r|���&�g�S�Ip�	��+�ZƏ35�&��56r���Ï^m��0}ey�t�bA���y�h�z1RL��['��9;m�����a\
M�o��-�
����:?�z�`%e�WG��	��ԧ�6����X%>}�ε[�D�
/���֤��L]�;C��p�˰�ߛ����{x��)���{�¦Џ��P�EL[�Z��S}$�|�=���6o�K�=Lt�Aߩ������~����o�O^�z8]������������n����ƚ����K�p�=�]837��G�]<�ո�X�w���|�����7�_{y�Y���w�ϗ��O~u�~�x�G����k��o�����R2�����o��N��U�����n�����x���7�k�}K��-�6��s�����Wh,>�Y��ݵ['V���Ep2t��r/A��p:zYR�#>CF�!��{[���@�ĥpC�3KA���[x�@KC����Aq��S̋3�vt�e~���G����e^��裏�xp�����X���>�#�!ɢy��,����U�((l^ʭ�{1G�!]���@!O��h8���:�8d�6b�bd?�Av
�Ęq�u�)iˑe������'�3�������+��xı{�ًx&�e:;"��oR�����4� A,`�8
��*�iپ��]��
J�m?�<���Dl �ZV�BK�\�>����w�8F�N�;7Y7��q�jŘ�m?�JT	��h� 3L�}�~���H'�*GJ��ɺ���&�QyK�&A6���I�F��N��e�`�� ����m�t����^Ǩ�?׺���=�ӻDz{��ֆ9�f�|��E�a�S�m@� �m'�RCc-#(���}���+Wh��Fc`v���1��g55�=v�5�w����s�R���I����΀�zXM��鷃��1�9���B������\�@w�Q����N-���)��%�8��Ĩ��2�^� ��TH����R<}�>��|��x"�1�(��pflU)t� �J�$D^�%���9�e�M�2)�L��rg����A�q>�ctiĽwU���c7�Q$Y��[2�<D�f�X�	PG&KY˺�3�R�j�BVb)+�o3�j��:�&��0�#�`	�� fh����^q�d��=�UE��{��6I%�qJFn�6�ܲSEp��Ʈ�	;��ԖB��wW�j�mKRt�+ƛä�i� "�º����f�6	� �
A!�!f)���cS#�A#ɪQ����1�&���{��\d�8���[�D�� qc����t
lH�.p@�0R���p�r�vz�֗-��V��'@U���B�.������l6%��T;��� c1-e��A&�lH
:Rx{�2pΏAʤrx�f�B#.���S�ة�)D�Ĥ	��/����/�,���|KWٗ�L�0
��P��!���!�#�k�EU|j�,3|8o���RGN�N��p� ۋB3�B�X���&(,�o��������p�*q�XU�o�g64�Jp��\}���Q۲+d���x&�ɧ�b�u�i�4�-M��4XY���pK�l�s����M8k�)>�j��� +����(Ĵ,��u�79?jn�d��Q-)�X����;�n����b�aL��� (��1F�\Vj�
 La�	2��1,��3d���c�l���݁������j��ΤɔG�ř��� !��qt=�(��Y��D�#��������,�'���M_�/����%�@����l�N ͪ��j�kŘ<�%���N �Pܨ�x�r4Y ���_a�8���7�8D9N�}���'(f#"���
��fU�k4 >B-�]��&OM�9�r1\/-pt�W5��%�^�SX�,�N]�4u	iG��-}m��pRb�̄��a�s>�lÈ��N[C(��ǔJmjU�1���I$\P\;�,�R�,���є��Kb�R`�X��C�F��J�#^�ґ�I��x)�v�ӷ�E�y�.��Hӥ��*�eօ+vo#H��FM��DxC蚆�Ԝ� ��5C���T5���L ���[�ww�ˑ�Y�j�T��. bU�M���^��}��xt�(i"mVA
g�I��Bh ����т�u��p�|-Bp���в�-c�H�&k�30�,M8� �B���-�j=�)�J�Gx��5��ZƩi7�|q��1��-y;���$KMb�����U+����s��ٝ �2k�@�h|��+�b �UkT��oN�((6�.
}��C�K�157�,C�4	�M�9��e`�շ*?����'Z����Rb���?�Ô�Y�;~���F�$}4���h} ҍ�nc7�O.�$�f4�k�}T�}�Rզ���F���*�v�}I��~�/�ʃ�EZ������t���g,��X�\��[�'?##�����Mg�c��§K������Y$m�Kn��}H�����{x��e �-A��C��b��tuw�Wؒ�7��/�"���?�1���	%���D�������Ϋ��]�l{��ͽ��V����yׇ2�Ū�7݅_l냣>uz��u>�����=��*.�av��Ǆ]�b�u6븖�A)U<�*[p���ϓ��k�ּ����M�!f�IA!�,�Ɔ�a���v��_ ��pJC��M.^��FЀ��0���\�3/�)�������|�&����ǿ�+�����J���i�y}=���=�R��z�{���n�vAG����6AUZI��<����D)���(ʺ)�R�S���e��G_c Mh$D��f����X�����Jm�@	Mf61�RUi
�裏������.1)����żlK��ƛ��E(�"(6�@V��%f�t�g8HU" ɦ���tVp&�6K��p��n9dq�C��5��9IH&��2)l �4!�D,K)1I�p����M�5����iI�QSS�)���X��k�Ah��QȲ@�WS����$�2c�A챀�l��u]L�!�֗#- '�Ԟ:	��/pw!����;��Y4"5%Y4%z���mc	��H}y�b�g<�v�"������e���H���M�6�al֋���>4Y|OanG>}4Rb�H[�.�&	1 N��쓄g�    IDAT����Y�q�D��xM�G?�����M�5Cs�ͩ<��F=) �ʲ{�6{��b�t��R�����Bl�뛤����u�����wVn^l*���nA���) ��F��0]�<��%��f>H����,���6�T1<�.j�L6�eH���A�Is�L�wD��d6@�����8�0�k�A��Z
l!�Z��(�X�5�q�)~�$|-���MUm'�)����Rq�S��^˙$B}��l��S���Z�0�+1��&5ݧ|�-�/5�l��ۦ��E�~8M�BoZʲtRP�Ж����N{�����t
�
Y�^{��J��Jj�����)���>A�8��jH
��D�3�-�lS�3D
�D�'"~O��G�
��03"���e�<2��L�oq�A��ҳ�'7�O9��c�R@�j!ju�嵶w����y�*��|4�Qk<�LL�[�r��<�i���Ō,+V(�ZQ.`8.�'[Y��%pʖh�h��!���TeHH�x�����W7b0K�P���&��Y��;�.y) A�6{�Է���3L+9*(�j�[&[�;�A1�/�Cx�{��tJՋ'��O3!��b�LeI����C���� ��ڔHË���3��#����@�Ҭ
2����F��f��ge��#��k�f�j����ŶO'Y~�\;��,�ɦSUj
�X�Z&�Ԛ�#H��!)���)��H���
 i
0�3ڌ�X
���@^a%|`�158�!w�R��U �_;^#%�����0��²s>��W8K��5R
��22�4I:��D�pd�5m���%�*46٤���jo��e��<K�*\pA�?=�,)���Ĭ8�Z��S
RU����"O�Z�<CH罩,Sn��-��t�Ĭ0�!7�e޴<ڈ7	��e�Z�`bx����رe
��5� 4�\�:�@��WV9���x����tnm!��R�jkQ-��j��D���|NƲ�Ԉ@����85%�dZ kb	7F%�B|?�Z��S�����B�.� P��R��<Yk��rfc"ն���z5	��X�!8J쁹��ށ�tJ)��phm�$�.P���y�R��h�Ğ��.y�L�T�.
)LȳU�.f�.e�{4�j�O�CSU	�ë�-�i�jS�T_�6A+ې��	JL�x$�E0�@��"�C.F�c��i (�ź/�>�@��T��[V;����������b`�tR&�đ�e�	*)8RO����l����j��!-u����Ŕ����JO�kR�$�W�+��JF'}~
ōZ#�G��Ff�e/<��&�� �ڎ.�d�t��IsUY�xlH��PVP\L��(Qk�'��,Ag#zeJ���:��kA��+;�~R�/E\�)>�=L胆��A?����-����O\v��e��F��7
=�l4)�3DhH]���J�y=���o��z���-��\��v�}�!O>�y哐�r��|��G���g��\��xv}�h~�����4{�{�J��ɮ?��x�����&�z���kq^���e
��<=x_Ҭb�O^z��|�
���/��ݻ�~����۫�\���i{su����^��w�=Ͻ��Ʃ{�����ӻ�W�7����K���,���\A/��4p:Ů��{�NF�r�݂�nACpAy
�L�;�vn ��,�|wZ-��'�{c�� ?@��R�}	�0̆!e)���o�G+@`�ҷ^$2YK 5%�귂ZA8o�H`�](�d�Ox����/h��O���O�Lg/3������x)	.V�����}�kM�^�N��DV��790/����J���@K�7[]�X�2K:���؎H�Iu����>}1��P�D�ˀmp�6L�P_Mi��X�Y%<Ck ��CJ0���R�4�7���E-�Jo���C�lP�@� ��IRԢeG�:
�7�,�#7��!�-�Jl������l��)i�4y�vQZM�!;XH��1)�H
� N�%��eI�Ψ)7C1���\��noj�{�)��F���U5C�8�Ь����HI�����p?o��O�H9��(໅<~}�_�٫�?��%0�R��^�\or�� �(�\: �X�84�*)�-n�J�X����p�*|S�����2q�����Ӓr"h�rjHܖ�N���#��F�v��M��ZqV^ef���q>fk�k��7��75=�H�吖�B
�i)�5-�&#�_jӗ�V�� )�����)���nr'@P�jyxAS6)�0R�. g�)�B,y�<}�I�He-���/N�g�
]q
�����@	�j�h�V�#�
x�x����A`J���e_�Ȫ�=ej�eM�OAV\�2Axc�b:��K�R0K���V+V>�����p"6̙�GVk(�[5ަ�<���<���C�T�ƉD�'������R���fI�m9P9�r�D��8����y����v�&O|�������;���+�;
y
6E�-�V��ŇXz�!x�!��2�̜}{�r��$E���F���F�'[�)��\��틍��+��⾕���w- j�H�&6[^a;�i��۷�ǝ��j�H�gK���S(Z�4���e^-0��ڦ�j|Y��Bmu}�-�y��/�jw�cI� ^H��rl���JY5��T�C��t��w~��7⎨�b��(,�xM��z�Y����*�w⩥9���
"೘�H鎏�,�@���qD1eY�,~�+�K6�� W��C�"��U�@��MsDX�	d�����i)�KL34��CG�BVw��
-��v#N�x8���QjR%�Ì/�iȕ�[���*��h�-S%���H D
��G�,ϴ��	��U9��l�5�l4)�r`��8<K�e���=T��Z�}"�y /+g=�G�@�.&��H�.z:|1���p��W+[;>r�q�8�B�J�>}�.(Gh�eł��AX
��%�N�l�����4$N|ڑ0��5��Hu!�'0��<�)cZΐ��
ߛM
G����]�2-q �`˘s	v��S����_���m-����6�N!B�?,�qv�g�Y�jZ�r8�~:�#Á�0aU��S�4B3��vlZ6������B����d�/��z>�*�#e1�	��ꮰ�i�&�l[(�ՑI�F������!z��xK�[�Y_4�E"�ڼ�WI��FL �+�
(��_=���7�2OAP�_J�`ǥ0��5Ō���X-��"�%kI3$5ٚ6��;yHF
�n���cI�Fywpd^1+k	C����KUK��h���+g�L�M ��{�ĕ���w�!<rjRIgF�r�6A"KG<����^S�����Dn���'�t���H�,&ZKj�ֱ��FvR�T�fC�qtϣ�&�D��,qx����B|1)��?��[N	Pm�ڥ��8�Ld|����
pLp�3�h&�.�Ǐ�Q�@�^��f�:r��S����(�)c���O|�c�d��Q1� �51�i�ii�Z�1�,Zc�Й����i�H?bC��@A/KL"��.����L���1y?zv&�Y����M�w#�d~�}�\�tFC^��z���phkؾ��:�Yږͥٝ`�u\~c�:���1��N6y�h^��f��f�7�����ʧMyK���a���V:Û�kpu�x�w�^>����7�����^\|�ܿ�}���4>����W�]x����཭�{�~n�j�:���#Ǩ����ޜn�/���Wֻ��,5�������~�ſ������ܜ�?{����9O>�����7�_�y<?������i��͇���������ս_�{{wy�#�w�%v��<]���Ӥ��6d}�6G���=�{@`�fW8=����f?|d���g�8S.Ջ�V�2��#��x�o� �)F������W��g�W�[��g�����������3���'Y:
8yAR�D+�PIw�^�杏����^�@ ���J�k��� %��g^i��R�!8C2Ut�a��i��{�˥1[#9����W%n/�7���Z�]54K��x�uA���hAq�dMN�$h�*�F/f۷d�y�Zq5�@P�A�<��xU!Kq���צh2�L�p��痊��^���F^��*3����5���ȯ
GIL�)ID��KE�Z��T�K1��e"��cDt�������g!�Ӌ k�ɪj��<��kl�р
gG*˔�q���;sH�2Ad���#�&f�$5A���#Ŧ,���(4��C`n~@����^�������-t������z`�R�m?bmzIT1�4�bp��DY�X�G3�����f>�̍��]� eVKR�oC@tD�Û$�%]'KL>>��QS�?R��Z">����C��)yU]�p&���Ѵ��1�&B"p��'V���i&)�ƫi��ɛVa��-���]~�DY�$
���5���^�xf�_�0Rb�@�{�l��#����1 ̲-H�3��5��y3�#(a=ک��8��L6�A#|q3 �S��Rc| 1�F��<j-ќ�V�����L�Ў��q��5U�R��������iJ�%�>Է���@D���8�z	��k�К�^�4�Zd^^j������m��WD�����o�R!M�o��";U�dъĉ`t���Ш�]������7�\GHSa&X߆�� 5!�V�˲�
�Y��A,��)@Z�E6'Z)��şC�2����۸i�-��x������4=�)AcuLG�<M�w�{�����ŏ�ތt�+�fqB�haM�|,=��}���`_~#?��<w��Ls�^Q�+��rj� ����7��N
8��J��*F���"��[��i
!Zj���B�b�h�8�*�oK^�����5w����hRd�/���9H!�b��1]Y�����o9�п�q��
K�q'��ڑ��'bY-Вի%ϒ���k���G+��`䂤d���u�
� ��	�e%1y)�!�5mS���tZ&�������X� �{��/���(!"+ �z�i৉���59��������E���Ҭ\��Ym��B!���
�Z]TY�)D �8����Ǚ��T%N�0)k���$���T�p����{,�[��h�̉�J��%�2~�Ծ}��ŝ6'�������M,���X;ݥ&Lbf"�X��ܪ%+0y��=�KtW�x�&�A%L���-���d;��_W�Nj8p�:�)�dh�SHR�8��Ő�נ�pT	�L��x����)Gw��J�,n�숾%\y>Y)A�8'�,/�Z�Z��;����R�0��ε��-w�5��ʎ2D�_a�y,�w�%�Y*�� hzձGY�T)QX	M���8u��!Z*�њH��d���N���p��	U�e��,��$^/�.FȚ(�L��3�F!e��CN�q�
�N���Q[��t��`W��3���w�hB�J�X���G׾�7�6&N:��-yj��&��hr'	LJ�r�	(0LU�F`b%�b��-SB��/�T��Z���VG�atI�v�&��d5Hm`�)�,�c�㫥#5ٙ��MS��@!�y�A��[i��R/�D�9M��F9�j���z��$�`~��p1�v�Cx:�(Ǥ"@k��{�p�<��� X�w�S��GHPU�X�ĒՅ�*����O*2|�)�,�Q�jy��8��=��N�{#���Q��G>5��M�33��(T۲�曤P;}�M��IA�m��
�2�L���٣���c�#XIR
�T��؏6t������~�i6{����S ��.m�os,hp�8,�V#�o;�t��Gе���Ǡ4yjhu�MM#���U�>�3�>��p�mĎn��W�(�AIW����y��������$��W��M�W{�~��s�F
=��s�������W7^J��`���if�>.ؼ��*�i�����{K]�>g#��[��v�������w^��߬/�o֟��^}�����Y�q��2���u^�n}���ۙ>�y�]V�#������[��P$�x���W]�n�;�o�qO���������ܯ���ś/�\�o�._���ܟ^8���7oo�}������_{Ly_�;�n����Q>uz��]������O�ޜ��j�P�u��I�#A ���n}�]���C9Rޒ�S@��{���p�f�e�Q�@7�e1e�8��
h"H!�v�	"Ǳ�DˆlY�1��p1�bʵ��.qTI��!���t<���������׈����G1���xOp�{��K�Aj�`�bj�e-=f�t�p���<N�T88���j8��(����*���t!f �"��8t��z%<C��4�
BP���Lk�F�G�jM� �N�!+Ƈ'�%�X���l{���?���'a�qyY�+�s��XR��)3� k� b��V� ���*��d�o(���O��Z���QI����VK�H�ɝ��AI�,��Gk�"�c 1���*4��Q���P-�����++�OP\/� ��9Yd4x[ ��XT	b���(wwaz��,p�yz��WM^v�|��'?��O�D�vZ��`��������-�!
i/��Jp&+F���<�٤T�c
���gc�쿧]�@����.�+��,A9S+n;�?g��̓Z]<:�P�
LY�{B����!4���	����y7M7.��R-��f08}L 14���A,&��n�Z;CK8M)}U��w�.b�:a(�>��I���G�(xLoR<#�D�04 Yc	�Fb���⥘�^dݢ�jі����  WU 0���%>�	X
�I���������uOϡۑl���CIx/Ū�B�ά���5�B���9�QgS���0�ዻ�S�QR��	�O�W��&�`-���6�jU%hi݇S^#^�,+N"Vk�l��x8+(;K��jk�Ϥ:R4w�%�^���ؙ׷���f����R��&%�#��p�S[*��j��r�ڂS�-�G�g	�6�3��Tv�=�M�#��f={�{�`�ăodޜNG_��<���a1y�8bSY�G�i�p����숤څ�d
{r�oP������~����S���u!��W�W�&�Es"7���\՚~>|�e�o~��A(�QUkK�p
�Y�6ժ���Yx}1m��}��:����ԎH�)暒�/�x��,2Ym��..����7��C���(��N�}·h����H�(��.�p �d'�C�������<�9�%~W�xǦh�*`HU2��j�5[@חB[N��!�_	r���@d3HX�E&^�^p>��b�{j��b"ę�IՅ�CFÑe�/q��Ù�U#W���m��Q8N�`������] �3x������$`Z��,�.n*��ë��O_Mo�p*�j�Y�0�	ĝN�ǡ��V!�S�ZDV�qH��h�_A 0�rK��2�@���Y�*�qM�I)�/���Ç�)�lڪ�:L4�vZ/YV�Ȗ��-��Ɉ�PH
S�C�e;\쾢��i�汬|
-�@��j���rħ_mjȐ�K��e���.��ٴS�r"�� �^2��`�5^���[�f��0�dR�30A��!�&h$��G�N/~�&0�h�%4 /��עچIG@��F�#C���ulI��3�Y*�'Ksl���@��Y�iT��eM�0��"LJ��l�ŏI_�j!��gJJ��(I'2���,mT8Sޕ���ưd�bvbM�3djbLV|��u�7m���tZ���S2LH{��jw�恓,Z6Y�6gUu�>�x�Ȗ��.�+�-CR���J��2N8��Q.LV�*f9US_6)�N�$�$J�0�ڈ�9�A:�^SR5��(��#����gڡM���{�k���a�֝	���S���1�lR#.���ep�RZg�p�o��ydV� ����r)��R/U���`�7g1?j鄻mүJ\U��,mY�5LKw]{I�8��Z
���׬J��JX��&��%G��]���a<ُ?8���+�\���&�0�    IDAT.�[�)7@}��O��F��55Ij�@1оڸ��|�C��3DSY�J@�����Í��=���K���&9�>���	J��&(n�	�ILo���[��d��.O�g��8n�t���Vs�K��
���f����s�-w`�\zc��!����~�7*_�=�z��G-�;�������7��X��!.�����:�ۙ�����~��h�Vk��\o���{���zG���W��7_=��a���Q��{���ë�_�����W>G���������o�}������}�յ8]��d>���~�.���u�����ɳkW������_��;�uD�2�!]�uP��)��ڡ�Q��ڑ��(T��v�a�
w�%q��M"�\#�w��U?��I�y����$��]�]R)k1P�	"�C}�SD�Z�(��U�A��<(����Du��{��MW�|�IvCR�S�yA�������ѥ'R�I�/���>���؄� 4Ō�Td��䮔���@�t��Z���0;Z��󿪞�\�DT����(�]_����T)�@{��n��I��tp�jGb3��@%��q)�ʦ��Y�Ĵ
�,=O�
�r��_��|���^�#Um���l��D��	:"����M����e�q �^	p�K�h|S,�p\e:H�D�]{�j�i�=A"Z�g��.`�YKLU@'L��#��0]���ApD�$��Wv���T��@1D���C�����]7��T�=`�	b�p�� k��aN���78�w�k$��U�H.���=��Қ=K�A�/(6��Z��ze-)@č���i���@��TdHK��a�@�m$P�^h��l�sA#�`��	:�SkY!���Z��%ҥu8��,0Y-���G۩��4M��K���AU�,��j��!)��+��ꈦ�A%uW(��T'g�oP!�C\���)�`҉�F�R� �h-������lJ	�������B��e����n�b^�D��4�ÇD�6�WEH�edHj�D��Ԣ���O'�SI�d�0fckǳ�DX�)��]R��a�D@klW',���l��>-V���غ*ם�<�zim%��d�d��b)���2$5���;G_`wf1_	͒��M_`4%�Z�#>:@����1S���l�p�X`�!dˬZ����d�=�x>��}DSSKS��c�� �,1U5OO����
"����y.��,�O9\�l_
�U^�8� o�p%pc��������<ٲ��{�x��gSa�ێ��!�$�|%q�a<��׺r��LBВ8r�b�Y*l;��k'���e���7|���?|)����.�/��&��B��t&N���bL�]q]|s�Kg�<#�A�h:j6vRL�T�8<�Sc�e!�Q(��o�!x&ێJ%Raʐ�g��Hv4@J D`4�i�g�n�Z�Ya"�ČԱ�TW���8fHË�d�Z7����B-,�P y�i��*��y�I6�Q
���Sp|N_J�{qLH�RIU�w��4����T����o�j�3U�#�q���C�FydUn q���
d�ܒY֥�j-]в�-�Z��Ǆt�U�kS��X�x���wG�"R�љ��h��T϶	��+�xJj�|e�_����|svt�K��0Y8K^�h��u}M_��ٔ%S�ٌ���j���`�Ų�,i<1�M!fgA��S�/��31ձ;܃�o���L��f#�.ŤRN�3☄/hΆ	T�(4�Y4`G-�/����̒�#AaRHѱY�I!0WN��Vpl���s��#�zf��R0%}�f<��{Mxc�����d�L��)�m�m"t@q
�,������ ��5�z����]!MV���W�Z��7��)���b���� π1��ٝ w�R�5�W+��ut���\m��jqx��3oeUũ�@�1+a��QLA9��W�����Jv��h��pH��j�m��MR�W5�lȦ5U@��i�C��������=�T�,e�J�����Չ_ǙM9_��h�pqK1��SHV<˪��(C�XV�{�����鬪���Ԧ����bj��闲}���Xp7��=�� 7���j>�ٔ$�)(Pi��S2����`6N�R�$|:���;�`J,���|�_|Y
�i�� �O:]�N��;���J���PPk�5m�Ɛ-�C���h�]UJf��J!k�\��*+���R�e%��#�ûR=����'�75���E�Ƥ���������<����>a%���������s�ד��>ݸ�R\Mӟ���R��㫯�~��o/��&/<��<�>]��>\x_�����h�	�ӡ(7�Vk1],�۟�뼸�?�y!b��Ч���Û�>��������H�^��ҫ���|�����wo}f����ި���Λ�_�}L�?>�z��=x����z��]^]�ýx�~��S��������ɔ�'��鉨{���u2�e.�4�K���eLy�`t,�ۘNǞH��8}>���B�y����U2O�)+����H7����3�ױ`���*�!�|��,�kn�J�ʪՋG ��� <��F�~���t�YG/�����nG.M���@�+�U�8p�&��-I�Q����1��mG9M82��I����#�L����iHx/Q`A�֚����8�b�Z��g���8�15A#Y�"�����j��(����A�"(��"pg�.��R�4���@�pRd�de-�4K�!�Yx�)5K1����/�#-4�	>)�`�p�мېp���#��ή+�]���KS��Д�j�ۗK i�␙�N�2��E��"� E��*�J��ƃ�lw�v-��Z
p�u�*�ۂIt��Cl���u�#|���s��l|S!���^��v��$���?��{H}��ؖ�f��C�4h�s�ڛBjM_<{Ӿc +����\r��&. (@c�.�x�:�Y3%��)��\��/�T)�� {Y�!�L�����m���x��������;C�J�KRw"�r�N[Э����>�.(nx]H���2S�]�N����,�9��p�!h��Ř688�e�h��-%6���5P��@��hR6!���8�x�X��p��2�\��6�}r:�"�1ۗ �,Aj<}�f�]�h��c2�e�p� ��v�u���3O>A{��dJj�$�c�&��RIR�(�$K��}���џa�� �0�Ӵ���NA��>���ɦ��@�dR�`G�eW(�VV9�l�x�䍑TM�O!)�@
�s��*^��&N�R܄��hL\�G��ęv
����=�G��,��� ����3R`����SS4��8]T!xֳ�e��=����������¡o�c��%0��P�/�]#g���{�t�=���_���H;ٞ��hT4"͓�k�Mx�##�Y�R3�Z`:q��NL3����;�eK�mJH�G(��H�`˦�/�F��y-���RJ,i�� ���~u�A��BC�*�����Mȣ�p��W.�5�c�[�#q�R�KA�]$�
�`�c�cU�7m|j~Ud�<�TYd�0"�*�莜��y[���}V�c# >×�{�vpU����v�ӽGA!��XU-\�.S
e�fk%��PV��&���R�r��������8�h��,����D�%/���Z��ݴ��Й{UGKd��h���$�b"��Y��1��� �W��2�,�L�M�2&��vw���I:��\
�h�L��=P�W�,��)`���m�i�$�
J�.�ɧ�,AV�iG�ZI1NT0ʂ�D"�9NO_��Q%v��5a"�Z(w&����Rމ	F�����7�T��i�0�4�#�T���7�V�#��D��"7���̒9�֘]��<�zO�Ȑ�@e���y
lˉq�:� �uG�*N-"H5��f0;��;�`K4�b̔��Ka�-�e�X�p"��<<q8)��-��(�9��mgJ��'�o)41����բ�<��C�D��49M%�Fj�eq��c�!�������	�M���Z ��v�q��)4C�������*��� �l��C��[��zR�ВNd"5�U1Y�8�8n�pb��&pk�;Y1���j��<~"-1���_6<��En�tC�3@qU�';Kp��L͒�Q�I�rj�.V�x�S<�Iu��Ӑ���b������;�LȐ=��R-)(n �uKe��n��)�m��b82�,C�ڋ�����@�"[S�6KA +��R 5����/�('��dt�xUs�
GpJ"K)<��] LK�~���j�1$q��)$ˋ]A�&PՁ XF���!�mVG
<ӂN�!�˲�ϲ��~t*�uD�y�rބ�@��/��#����[sK��/^]��Ӌ�n�.s����������$�>�K�B;��F�߻�w��}��q�~���X]��F�ׇ:��8}����y������?Ly����f�'��	���W�7>�5���]�>��v���^�xv�~�	η~3����N�5�����c�-�xz<��l����>k)~\G���߮���K��Z�ϱ>�L����5����W7>y���u���~r^o��7�}��C�׻�g�>���}՗�[����wAvd�nB��
:@��bb����,p�c]})
]����v*���Vy��[��F� C�K�ݽx�O��Qش���<�C�x[��T�� 9��1%�}�]R�#��(�i�un������_|���R
�p䟉ۻ]����33 C&���%Z�6��ȼ��5�XF#1CZ��~8Ϗ���?j��ٚ��]h#u�ፇfw`^8R�Ī�(i�J�y
�h�Ɣ�Vd�x1AA�^��n!G���~7y���K���Çx�ݎ���C�Z������R[_������h0޴�f�.���-ߓ�3[P�,1PP�,�CV�WB�	[6R
���%���C�[&�cJ�CP��`:�j���2A�%�O��`�Q�S���k�������av��5)�\k�.���W%P��\w8̎�F4j*%�|������п�P�������6�ϝ�+M��H¡�;}��h�q����Y��( 6z�-��bb�x��2%��~�w��3|d
@�Q;����w	f��,)���G�/�Kos��R��@6AM�S�]D0~�5�)g��98���:

�:*��=����'�&��J�.HP@��(FF�������u���Jw �U�E���Y�h��eY�\&q����zO��%�[S@��؜62`8�)/B��@bɧ�7��ȣ1)^�	M3D
�g��w��L��S�~4�{�:������|�#R���}�@a���-�3g����M,h�-�dʇ�����*��Է� ���4;I"�EM���GV0�]�J�Ԕx��*��# ��G�pԊy���Ҝ-��~g� R���BTY2;�D�)�9������T֭b����V��d%ek�
=3��kWk &ĲB|>_wߚЇ˚��)@c���35݉7	e�<D����2�-���_�����o��׿z���o�d��wEb���[L�7X�k�}��U��T�M��,P\���qH�W��&�S#CH'egb<W��fvh_�t���	�q���L���� ��+���v<�o�ӷ�噑�p��=��S7��L��䫪�s@��-��?BR��lH��p|��!�J�)�Ȳ
�:�+��o_:"`6���� ����y�%�C���u&����������rsεƇ{UQ��n�Ktui9�V��1̬��I�
�ӟ@
"�C�.%(�@`�,�u|~L�͌�Y9o0:deyKx
b�l|1\̀b4 A��)I�d��}�1�j�qZ�-��*����r�B^���8�m�!���w���@�ID0��@4�쐉��Y�4�'U����j�o�Wǁ8���Z���z�k׽d���:.�����R� BAR��&!�l<��,�P�H�J�FC�&��� �̤�f�t���I�tx��W�ҲS�B�2���G\����X�cߤ�Jg��w���X2�3	��eA%bRb��;5�q�t�Ѐ��Pa"q�~�p��D"4�X��$+N9�2kY9�����]h�0�^�Z�Z1k��a�B�u�RS�OPU.E*��=6ؔ�Wax�dSN3B��dJՎLA<�f�I�� ��0M�����@֫fd��<���%)^�sv���yL���m��&T.�B|�ulJAV��/��2��� _�A��d��Z�Ywl�DXUK1�!��� �zH*A���j��-�*KقD�Zj�L��F�i�-�t	�Nd�IavE"��Ϗ`c7[�]lKP(+%�TXm1�D�IMI�D�g	�T�D̖�>�@�p^w��$L �͖>��S� 2|@�,��uN|�=��m��-y�H}�DS�!��DkT����؍8���H8b%���(�L���M�G��~��_ٚ��o�*���g)[IA
�ڠ ^��󑟳<���T,P2������(8XM���gRE�W��!��L��w2gkA�2�r�m��	x#�߲�{X�6���6U��pφ�:
��<���S5'Ado��痯"3�t/`���K�j];����0�~�l^aޟ�_�<�	������ށ�My�x����t���R;����+�;n��Won^�,�3���u�2\}�
܋u�l U�2ݟ[uh�ru�`�DLh��n���Og~�ի/����s�_�2�գ_1�p~y��>�W?�럯��ߏ_������}�p�Yo������o�ݟ�[G�W��տ'����� �@����� ���q��u�{<��A�)K��mC�B�;'��Q4�vbO��
(���}#��[���᧓�
�H�7'�ZDC`�M�f	BY�=ĲZ����+&��l�N#߳�8f
v��z��o�R��}�ư�����t�֏�b"�W�2O����C	O���#�(�*Q�@<����\�Qch፧_a/sI��*�LS{T"ҷ��F�e-�F�;)�M�l٪�L9AA�Bx��d��fVB!Ax� +�4�z;���'��� y��K^Z��i�G4O��r��ew�r�y�*ɧ�V���p��u%�����y���C��δk�dɚ�rg)�Ǡ���g��֝�Bj�L�����c����>����(��~��>D�����]�ѡ�(`j'�JPܖ�ߖy)�9D�[�	"w$K�u�ysM�/�~�����f�=�9��­��b�������U�dz3�����"E��l3�;��H�e����IYӡ ��R޴�hA0�8~;��<��@9B������z�V��xīBvVu�/:�h/�����^֒�@��N-�l��y)%��]B��������(d�b��^hK��:�
��!g�8��D��Z@���S+�U��<��ҬQo���,��0�#`�
*Oj�	��SS���H ob���~�tAf-S8"�@�:.Aq+l6�b�!�`OD�R3�%����eC�Ť_/^�x�=���B��������K;�AШxF�6HM�8&�CȈ7��^
k���4fk�5�>C1��hSXm|���_��ūU��
�8J�Fh�e9�D��b�\�6�����e���@�c�Mb6|�8�fOD�Q�;�p����o*Y���'A>1�X�RnU�� �Ş�@<e�%�\G����'@L���1���y�TN�BS	��g{�f��j6A]����s�~[��f��w��<�|#l�WKV���K���k;4�8j��������A�j��4�(���r-�3��)@��	�]H��!UA�Y�˿����=��C��x-��Aܙ�֗�4y��?�X.Ћu�#`��H����t���|jS�-�8AA�Vz�(��$L6A�T���X���'D�{C� �F#g)8Ip�U    IDATU��������;m��:�<
�&)�����$��������^"��
1�-F#�K7�ka~����uk���<O>�d�s��v��1K�	1�k�FͦU.~��
>Ŝ%������8)G0%h���6�,Z�!�D�_	QV�|6��hk� 0�d�i�h#�D�,%��rZ�N��iV�hf�����l5?��q�=c�p�t��@h6� ���>Q�kZ��u��������ь8�5"�*V�i��k&D��Cn�H��z@�(5~���Vz
с��2��N�S���!�� 81�Z$��lj��*��/�	�Y�i�.�|"LcƩ�A6���-8����#�'K�� ����Nʊ&W-�ҦBF�ڈ`J�Os1�P|cR�#����OЎ��)e���mg�=�B�$@��L���|;R.��QV�B�(��G0��[+�[!E��o��rh�q�1Ӑ�����-=��ժ:P�l�%(7���$���m~��N{Y:i.�mi��M���=�Ѥa�|�N�V�QNY@�
1��M��Ͳ���*jLR�����fҜ&+'�~j	ȑR��R��99�cZ�@Y�D�oZ6���aR"���8\z�G0vB�b��ӻ� ��r�ig��2�M@k�8)UА!�YS�BU�sB�΁�0
ħ\"� ��MK���c
%�q�C�F�3!-m���p�S.\nE�+��b�+44��SԔ���.���1��@ӱJW��aUc?-�����J��tS��	�	|x�CPi�iV�1'P�i��������s+������M��]�#�W�i���Ӗ��Q�͐��ܲpJi���U`3�DH�įm>��>5a{������s�)Sz�y�@�1e�2�M�K_��:a�v�Q�f����K@-�љ]�_��_G<'Nќ�H~����<�C�����>G��w�>`}���×�����t�ɛ�\�}�s=�u�l��7W�=���� =�=�\a_K����=�M����⺃X�.��k��\_X�x��o������ʗ���������+�9yy}�>:�����>~�����������_~x���WWo>xq�����W<����Puu��W���U���p}v�E�8�8�����Fl��]G���e>�x9�82g�Qt5�N�U�;�8���N�ҥ�c:=z#�Ө"�Q����� ��l���c8&�aR3���+��Ԁ(Y�eZV�Mi�4)�H
�R�t��%J������Zq��y��3�_�����EٻF?��=���(�Z��L8d��rp���m�m���(�h@׸'��+�m�P)��Hm�$"����d���1�F`]��~���XVK����c�e
S�}�r�.�ݦ}��>�.q8j��I�3!4;Q)��!���0�<{�ɖ(&��JO�C�������[�$���+�V���#O"��k�����t��UxDk������J�7�Y��SC�q�z�o{�x��dR)�FS4#Y�&�����j��R��L;�4|�m��~�����?�q;&˙�z�������A:ǈlԆ3�O�e)0�Q3��P"���Y�~�t�Zb�3-�\��<���/~��O�S�#�L�Ə������o��.pgm�jt�Pi�t�o�p���A�o�FY�R���}2)`�-ٴ5�Z�����9�v'}��,!dY�o.����PE���z'�\%XmL����cY
�C�lsL��\s �_4��?���3ʥ��R�r�}��/e]�ޮ���y�*]2�약��6e${�ȼF�M�J�!�}~����:����z<NZ�I2�1щw�l��p1W�mw핑��[:QT��h��}��N��<qE �4L���j4�$9%f]�P�ꦶ�|�T��D�mj�\��홫��03�=��;ٶҺ�膩U?(l����k��*�G�����/�w1h�f��6�L֨gI���yS;=R��aE���^�,�_!�66 ���3��@�)�m�Ma�9�x�MS���XG�=4N.�(�+��nMa�@2�0M��n��0ap��|+�=��[��DI/�!�Kb�����E�FV�z�,�d�B�*��|2�a�k���+o�!6�1��NZ`{���.Uj�v�XG�o�P��t~2Z���$vMh�I��YY�)�����q�-ny����W�|���d��t?�ս��%'{cF�X�M�|��M]��+�7�k�_XV��oڵ 	�aIw󝭪-�m��R2����e4!�$� $5֓���s��I�ݒ�l��%�W#�����"�A������3�v����*��#cGM���J��1�Ο�7!f9ˠ7��1��'Y��r?���d����{=���%�^�(�0-�F"o��$f�d�([Q��<[l��!>�B(�lbT��ݶ������7â�Z��0>�&d�����˸f���a~Zh��C��Dpw�pC�P��ByhŁ�?����Y�%3�d���Ȕ�C{�gb⎤�-���]/��ʩ���Fu8��KW���OoT����ꄝ ��u7ySf"��h/�������9v�U��E��V�O�^��~kS���yun�.zh��[�ьQ4Zҳ�~�n+F�xY�p�0�:ɔ���_�X���[l��ܰ����8[�����/�M(���s����~�XY(�-�kA��٦�pL��۲w�Q��+í�W�ׯh\�U|��{E�H�@�UY`�T����WKO�g�7R��U��*���+���ל��cO-33Ot��ͧ�2�(V�d�jzp\�]�d/x�s� ݾD��R��&�����x�Í��_8>�'��'|�����!�7�c;����`��Ƽ����[��~�nXc�v�s(�k��OAgϺ��ɥ�ۯ�S��������&���A�]���x�U}�a�W����!�����C7������R�C9F�KQ&`2�v��\��_���.��ʬ��P�"w����:P*�i� �͎?z��a�Xӡ��ۃ�9�zai��O,�C�H�4bc�+'j�;�T���J��1Ne��Idx��J���0,�N!�יs�{���˝��?�*k�W-#��]�wSbY9>�n�ώ!�x�3Y�0����]�4t)�H�2��WiĻĢ��6��_߱�BS}}
}PIv��Q�rAۼ�]'w����WS����J�	��G}>��X���ĐR�������ݥ��uT]��)���e����R߱�a���˟_��Ǎ��<:h�%�u+��}}�u&��w�&��#���r׳��nQ�&V���C�`P@�������ѝѳ�ϖ3w��{�]�5펇U>-����RvV�_�|r4���������H�a�|-6��L�I�r�/��G!�'cϒx^��gf&Y��zu�>x�7j���/*����8����`/���x\��t�u4��жbǁ�.���A�����y��aE`BA.����8���ｏ�W"w3�����G�ϫ�$�֧���C��-3�����W����U�5?�<W܄�4��y�Q!Cȷ��A����7�ӓCze�۞=�uCB�)9~�%c¢t��������>ˆkq!?㫻�sZ*�8��U�O�E��*I��j���&�A|  �ϱ���yS��G�,�,�"���<��M�V�TE�X�!v㚚mr8�'��p�&�O�$�i�^� `�T:1"}�i���\�KZ������%�T��i��%R@^b�C���/nω�wy$�{�nHƊ�[�����>z"�W&�}��q�w����#�c�5lu�Ѷ8�X��ygͲl�4iA"�r��:�������v��v�Gv��O<�6�j�p�����3d(�t`G�����i�,S}���BYu@�؜X��A`�{ٟ��f�Lƕ����/���M&a���>�Ϯ�m��xy̧x9�������>����e7�맛��-S�rAc0��Qb�?\BE�cSI柝�fx�������+���E���o�����x�1$L~��ٿ)��WǷ"�Bآ��s� ����(�=�N�B���ǩx@UieȜ���m!p��%M�K�[��t��������;�Ϻ!O�x�=�OBY�wX�$`�hP+��9R8׮�����~���U������+:��a��#!ޏK�n��)sh<�:Ǫ���.Cv���`OAGA:v����h�X�s'�*���6��*Um��q�����%�!��@�a�� E��<�)���!��.TO�UA']��@̔-�����~@J��]q83<��{��~�6�T>��'dR�r�m��{]Hp0�ץ�Ƚ�`�4�M`���4K5/����X}�85R�$_�W�z���ǖtW��:м�]|˛��o�}v%��P�y�<#���GK��܍8GIG���a���?�3!t��tu���j/��V�	�ʻ��YXs B&�n>Z�GA��� ��_)nu�P5��j�8x��g���yGYs�!�I�ɍ��WV�[ܲ�-D�\�W��� X6_���Ф��d�`���	�w�P 
f:����9
���!���j��W���o�2ߐ��<5$ŭ���h��I��^��7�ƫd<~L�~Ή=acA �"ĔY�#�,(����x�~��'�jfؕM���
���H�gb�.���q����Z��!��Q>+mp���жs��������_��b�Lq���hWH�5U���xB��\#����U{���r�z+Mg�@ca��Q�AT�Y�
QB ��8�x>����U��9:�=5PA�O։f{2�8S�����- �Z�������K�X ���)�.������O<BV�`ơ�\)��O�������4�l�,��ݟ-��d�+�3IR���	� ЌO����1"�lBf�@"M}�Y�2�wWYS�u�3�����M���1u�o;jS�#gd��K
�t�9Qi%�#wb�M��u��"o��VT�.+�Q�V��	_���@h�?�2w�s�++t����mU�:�C]����ڒ��+-;Γ� 9�)��'�]��֩����K�F��>�~t[@�)����{�j+5 ��w�'b����#'t�<|�cfw����枸܌���C,���'��,�C�Krn�_���'���Ծ'7Pk,��]����PB�f�ʩG��)���d�l��X	�Sc���//*~\r�ޞ���$68�"��i>�}a�R6��E�_?ؤ68�*ٓ&O�[�����{voX�йT6�32��zS�v�6��яy�O�Tq��B>IG����@�m�O��5�d����>wqEZ#���H�EM_]r	=ц��Mύ��h����H>��^&�u|*\V�k��<K�0�K�>��D�m�̠)�����R��>JW�Λ�3$.w��~	˓e1r�j�җ~��l���;�����8*b"+k��]ѩ���3�Y*���I��._��y�*��$3��m�>5P�C�6޺��v��5b�y�78'Z8������g</_��Y\];��.�>�E������Tqi�]��q��Y�ڻ+Ȧ��l�D��3�ŵ<煝���-�˳��Ͽ?�M����`� �
��[+ik0�Q����	y��߯v}Z:�;�ר�hi�����M)H��ӽ���K_�vKU�^<kML�;�x�@W�LI��[3K�pқ��ܦhS�R��6�?o�`8m�B+�z�޸S�n}$e�c��� �ʧ���צ�"Y����m��6ȱ$��ek}���h�t����ةn����oX*=ܹ�v?�4�wx�~��xs��9%����%�q�v��̌t�̇��Fd+�^���ws������y"2S���5N�KO�����~�5�'�O��ra����4S'����VF�@h����0@�w �AF�)o��8Qn��H�P�j�i��q����3� �}YS�C�5������w]�1_��u��>�`�Z��)�{m���F|���8��L D�+m�YS@�=C�j�l�D�r�C�R�s5�ۂL���}����s�~��J]a�UҭtsLZ���M4r���X�T�lNlΚ�G!ً��?]�Vh�k!�C���Vߋ_+�u�g��Ϋ�W�L�=����\'N��3�y��[O6��3aغ�z������&�W7���#���'��Ns)����i�1�1,�45G��f�R����g�:̷l�[ћ�ׇ𿂓�9T����"@nDs~�.�A�	����3X�&>�^q�Z�����k�_�{�a�Z�:�����pT�	*w�uU"�[jTf����U�β�2��~�����Yj�rl��DȄ��r�b茐����2m��U$�
ӌb��O�t�h��~�Eon8싫�$�J��&WW�c9�W�Q��I����3���"O�+֯<VH5�5M�X��,���%rB�i��u�}fiD�i������~f�ת�|9��]򳚢DN�eyfp��.N������i�d13L��#G]Q��@UWÍ��#����0�:l�De]��)ϒd��?��~��=��{���aLMcp��3�M�MQF�R�K�V��j��]����4&�J��^����j`��r���8b�ϩM7�F��lp.�3AK�	/&/���k;Ws�(L>q����D���!�뻊x{;p��yX!��X�R��U�oE�X}uB�&����dCW�[M�T|r���j�)G�����?��h��Tx+��F��7
�O&.�N�N3:������Y_3���WJ�Bi����P��v�I��,x�;�V��0q��a�"�,�(~�]����$�d��O��+4��;[�٣Ql%���,R<ޛ&	(N�!,N��k�M�#%��)$���F_�Wpn{)-XG52X�p�O1���dVO���,?�>��b���q�9��F�"-�([m��+G]o���󑫆ҍj���N��>���� �,�I$��Um�#z���.Jr��	�f����%����9�:?��ۜ�X8��X4�);.Q��Q�R���+F�q^�9j��1�A��5��4���ԑ�ۭ�a�E����U�oz��Pj�o�v2�fW���c��98�Av�ʕa�Z<��"� dv���M@���A���0D�XX=�v�˂���t�r�.���b�V���d��TO�
�s�$���n<�au�yԑ�:qk�� �e��*�c0iZC%����E
 �Q�}l,I://c���F� .䗊a�9z����=Z�W���U(�S����΁�z`g��.�pq|�����wy�}}M^nsds�k��ѐ-��:�B%89�/����Å�D���C�uQ�(�o\�_|�8��z|L#ԓ���4��)��Q���H*gR�+���BH&��ML�=�w���Ѓ#��'N(iy]֢i�T��NO��ɥU,F��gô~yD�#5+�?�Ͽ�kǉ���6�r��x���le����8��}Y�a!B02=�n��]ϖr������~	�fv^�0 6`T��%�U�c:{�i�Qv��tV�Zg�ћ�A��H"߉��?�{�S�Y�}A9��I�NC������*W~'��И����M�HA*�4��'�+r�~L�	 |�{\_Qa;�f�嘕����T3HƖ��B�/�G��O��'�G,�:#�g[����?DiIT�ڞtZ�����x����@����v����&O1�e^�o���?k�d=8��a}��'�;�eI�[~��"����-����|��s�9�A]����/�G��B�)+q#� Iw��cW��ꝃ����vq�=*?h�Ɣ�����as�w׾mTz�,m����.��dY�Ѯ��ʷMQ�f)qy�A[Gsǋg/C�vr�;�;k��洖����]�8;[͝�3�,�������3�1����^(*�<�.+��}\����7��_���䪞%��m��֎giX}��[9�v�M��m/�L�@����C
$�^S*Z����_�=��Y�Wu<� w��7g���o�f$S,�s"E�*ɠPIV��	8&�Ą�!��sWq_�����l><|Fծ�ْ�D<vY*,g�Ru���#Tj_�v�%}Ih���,���'3Xؖ��l�����}����j(�$�v���坵S��aIA�r����ҹ�}�Ҁ�)^OE@��]ڏp"�����r|�k�]�m���?E�G�DD������������q�.e�l3�~��<��1���
:�j��'��'�NBq#�f�y�)��ɔ��^DM��U9sT����A��*�P\/p�j������w��8�8�WX[��>�T�1a�7�����߱�ŭ(��Hg���um_$ּ�;p��Mפ�SP�1"b7�
����K�!�Fe��r�8�2���R�sl�o�����+ѳ���v۵���x�nM�u����P�%���~��߈&��U�Vj��9����\F�0ᙆNL˂��P�t<#�@�!gLC�߁ߗS~.:�RGh-�v��K��#�s���N�����'�Ơ�R�L����P���`�ye܇����V��p�'�2ho?k1d���󰷥�D�"\�W�C�,I��O����QnC�Xh�ʙ�X�iP�D"=�l��"� ��	�+e(��������[��i�������<�ʪN`|>���U ך��4VX���u��:���d�z(��o>@��=��{�ᱰvj_E�0i�}  �Gu�yN�JsV���T��%'�"J�Se����WO�JQߧ`��yrY�a�N#���K4F��ޖ�Ӎ�����������:�ER���AÄ�/�v�.�U�5��8�;����ZǢ����9�w�P��Z����Ʃ�K��I�X�y�dW�K�D���"���A�ы(���k�]_��m
�@�y���,��u�"�g���k���1@^|��Y�*��I�ñ�=�#���qq��5mgz�
xZ��Z���lG�Ev��UH5���-��
�ĿD��-�?�|zf �j�5YP8^�\�Ŧ��WcC�Λ�]���4��f��a��]��0��jJ�E�J2`�R��@��f��"�=�Cď#�i Y�ꨄK��=�U����j��
3(���s�X��q-�3>g"�Q�j|!�����n��F1�VӊZ7�@���Az��w��/�����y�,�c�|����?��.`�O�W0���m_�.���,&vVr�5P�+`uޝ	?Z�u��neVp�3��
�QZTȨE��e��dfx��6Kl쐣�z�>xH�s���h�o�xV�X�8�o:܈�¥o+�v�2���ơ�.���GN�;�(�⏛�K�q3�)3r���nh�����f@y�n�NL�7�8�v@7/z`����0�Eа'��q#�愿��4���z�\��2��w��I�	��L)u�5u��{z;�'$��_h �sN®a)��
>a��p��Z�m3c�W_޿�VN�}ˋֱ�32��9��SI���8�����)���0���Ճ���'1Y��z8N>m~Ù�*�p=Ɍ�q��$�~���7����W'	(����/���u��{SQ�L����v��C�}9�/�Y;��/��b�J˕�nXD�7Nt��o��p��	���D�Nc�~P�.���1��q+�fA����P�ށ��J� ����<��\0�i4}��.���6	؏m���rfa�ԣ�E���L��%����>�yЍަed6�Ρt�Gu>b����I86V�#s�c��9ן����|}&���٩�|}�o�U��>�I���l�%%{��'��E�Ǩ��e0
D�10:��+�Qw��~E��S�����D��(!���W��y��v:I@_ӧ��l2��;��D,�2�~��N;����Y�&�`ҲH�Ο\1)�K]�G'nf������˵6���d���a���;V�;�]�T{�����	�9��h;�V^Cջ�D�oS.#��6�v�^����L��{�{�%�Ck��l��_�y�,���G������XpZ@���7����/�0/��
qmʭ�s��I.y�&u[��U�ܭm��-�y���gs��' ��E��������$Cᵤ9�6�M�x���_�_ss[�J�ɗ��bw�W(��n7'���*�->�s���k� �.)�#��hKMiɟn��S�u�7���季�H��d��w�r{�hI�&3wS�T�)��7;/�e���
���$��]�4{�i�,e�sÈ�� �z1��IM5IL#;�q_C+�.Ҹ���Э~��e��P�Z?٤��L��o�{1ׅd������>�<��kեKKp��4���AMf�%��o�8���������b�͟	|1X�*n6���m4s�FCq�$�+`Q5A�4i��/ F�"�e�<��@�OX�ʻ��1rFA꾒ܟ�c�i�-�1�P��tk�W�3��j4}�.��[�six���r���=��ph� rc�tI-��i��ai��;��>_��l�W�����	x�pڻ3j�O6j�%��N��֎}�F����v��;#Z9��╽m1m�}1��|��|C� ���(.@Ǻ�í���}+o\�M<EC�n�h�@}�4TV ����i��	�d�,oZ"�;�r���5r�i;|i!���+��+��{�%&��9�� ����9Br|�ցM(���d���G|Z+���"�9pH0x@>C �ٺk��C��O9�W��kc�V�k��ܗ^���ܬ5��M V\ņ�y�d������Ϛ����2��b8	4�'�۱Q�(r3�G{���$��]$'��C�	��̍"@�����������w�V�`*�ʟ$����	M�˛��/�ǒမF`qƺ�4m\��5C	D܃s�:�7}\��N���� �*0t\�yG�-@�(]q?�JX����� ����{0� (��@��`����0!w�L�?�&�K��,%��2O� ���>��nͩ����OEJ5'��cxBŔےM@cb��)�w�?�9ڵ��U?Χ6�N��������>��7�������9��d��L�&�E��hS�s�^����ot�S(���Ъ02�;�Z��0��[���;��'�f�� ��;��J����F������&
�>��).g^|�]QY�u�D��ժƼt��W��*�:"W{?�S��M�x���^����U��$`�r^���x^m��d4u�Lt¦5s2� �A\g辚�(h��߻�Xt������p��;�B�-h�ۤ���7ϼ�vT`��A�$M@�͇��!����zYA^7N�j����CYw�^�A�!Ӊ�ӎ�I�Bd�GJ����H��Zo�Ua�-	��)T�I�6<���a/�,�����kck��=v�t�TFY8�x�i��1t�ߴ׬�P��Us�R@��.�LQ�夡=������U�ʳ�L^d����0�}w�T�7��x�2,��Ć��K�إ%h�A��k#�X�5\�le�۹g����%f^���6�$~ԑ��w�gĕ�+�C�5�����	��A��L?���&(kb�Ԥ�����*�����l�܃�7�=�U�N�>|cѹ�*�Z����"ϰ�ӹƂ���A�ca�V���03�c�d�S�X����!?��LFBWaܭ�176nL5����{S�iI�����!���Nݝ4�q��F]��j�c^K�L�
?��|uk���z��݀>[�Z�|�?�'���@8�A��#�M9_gIy�V�8N}O�1sL<Q<�(X	Z�r(� \�/���dс�������;2�o}^��O\��*�`�\h�\���Ut8a����h�t���>	�W�`���V��4����t0�pܝr�Zc��$�15�r����f6XDNu���nȄ���P
(�a�I�(���dE�p�X"����V���9�]>���.W��|��$}v�e��z&���V&3���*��0*GnW��@Q���Mzb<��cb������PDh.�A�/.9���M1�����2�OK�������B��ɺ:Ą3��-���|^���w,/�A�� �Pع����E�]�*O7��H���^�<�r��?nN�C��KU$�[4	�p��y���|�<�)u�d���� �>CQ��$�@�C>x"f�%o7���t�� �c�Fu�lǞ�{���T<..<(�%�QSM<ڇ����F�g�.��Ѹ��5�&��+�t��y>6v�լ�̓?�O3��`��g
N��\�ԥQq�/�����-������,�峃����X�����CKO:vm�7��meޝ=�[�x���<(��	W3�{��P�Q�F)��KYūLQ�	���@�>����aKm�ǻ��B��cqqL�m���A�#����Kr3�.]P��B.v�j��ώ����^䧏]�W��?|xux럗ĝ�Gy��U�EG�[��_:)�S�4&������w~p�_���<ݺ�l��>��;�Ӵ�9X�SȪ������o�.Q���F�o�h	 �E��%������ū���8&u�͸3��}\a�C2�Q��/���eV��(��_�c�{��ҌP��a`2�����j�ܳ?� ��W[���m�,�(q�6f�6�� H���ɆpL�-R��]�`��]���^�y ��`
�qҰؐK��"�%:��rr��*:���,��$"2g�͔g�̿��S�e6;C���� �_,��ˠv�l3ڴU����T����(�	m�8s�ٲK�iq�JϚ�'%o�/��}���� S3g!o~6O�����<ƣ��s;��P5}��*j���Љ̥ư�]�H���*����ub��b���ָ��OEK���A_��p����V�T|l./��-J#o���e�X3G�^˘Z���T#��^����/���ލm�v���Q��A��q�w^}���n_6�i�8�e1�zuʪ�r
�cz��uܶ��Y��fFt�e+}[�H��T{j�Q�<��r���E�'w]=��@����n
���_C�*>'���Zέn|�h~$N��}�oI4/M:�K!r�w�Y˂n��յ��.��Oi:�π֜��nE�|y����o�
�pF�����z2戆w�yu~ik���ism���sU�D�@�9��3��������j��"��V�Qo~�f��=��u�oΛ��N�j��YF3�jW�����*ûN~0�@%*�(�Փ��~�p`�mDB�|C��M�Uf�L�|z^��	����8N�1���&��F��w��"����SM�Ս��D��mˊ�p����~_�dL���;C�%�,\7M�	��Rx����ㅙ7)�S4��m�����O��@">d�6xZ}��t;r$@4��g4��6��Dg�2$��"��[��#Z�+ò"����@�����J��;J�)�%@��3Ӈ\S"�oj����Γ�8�vy����ux4�m)�����M��bhd@=P���
ȣ����:?��䏄�2�z@)[s1���2�~������^G�,j�~�W�e�a�}�V"��l�@�p�l���@���m`�է��mS9/��9�$����X-3���Y��1�F��s�[����\��I�+rN4}s�� ���,�B|Nn�Z���B�.���0@U�z.Ó��Fس�d�9��bUDYJ��m����~w���X���1�����R(���*^5ɑ~}w��]K��q����+6WZ��/�7M�T��p�gv��BNG{��$�nM.�Ky�
�"���h�t[齦�%�m�:�|��
�^�K۠�.30'D�rk�P����@R��PWNQ��1�T�8���Y%!5��w�+�E~3uƧxY��"��e9����dZ���t�X�������m,B1�ux2�'���U,��!x����D��9!�ĕ�]�����(a���/��X��C�=Z�d� 铤��T�®k�T_/%�������c��p�ߝ>�CW��M������׬��|�!9Y)�H��[�LI]:j0�1�^�ҮV�z��� ��^��	'yR3+�_�����ͯR�f�H8H.a5�;7�����j~��[�[0��:����$�*�v������M���e:��(�x���d1}�2{7�!y�"#x��p�k�QN6��M��V:C2ȏn�^-�|J�a��G:���+ <�B��<x}��#�J%b66��Q�I�ue���/����Ba,m�z-�+�������s?�>��,�f5��v�;(7v𔙭7�HI�2�Va��H	�t̶hb���1<��0�U�@���d-�lȦ�2���;��P�ܽ����CVZރ����6oYc�����V�&�!Y�nO�a�6�#�,�:-�c�1�
`���ѵ'��=	
R�]Y�rJ�B<iV��ڗS�����L���d 6��M�u�p�?�.cw����>���϶�;2��LI��Aq�����Q�J�Oa�#'��50).q+s�O��Lr��d3i�x�}]kK�#�;���u+����9���?x�M޺�����vH�i�:ɰ��,e�/�|���O/W�SXΕ����@yi�6�%uK��fҺYٳ|o���}R��r�	����Z�{^���=�ιk�
>n��3�97Ȭ<�9�����ϒ��{��%�V�388��?�EK˃���|������ro��^��tk��~d=w0����Ƹ?��<Ic[m�ĥ?]O�T��X�(n]�i�/^�Ϥ7j�]"�I���7�3>ꂎ����b����X�p�1�:[8ǵB��7����bVˁ>q(42�ނ�.ۼ��:�'V���7��P{��iu��w�z�n�������+��[���
�|m8Žϗ'�x�is+Df�E����-&�DTt-�y�up/K�k���A������Y�>�4�r�*/�8B�I�&K���M V�<��/09T�W���?�h���U+V$uU�2r�<���y�X��C��~��v,��^��[ƈ������V�Oq�K.a�ʄ��T>��mT�{����� ��\���C��~N�W�n�L��B:͓����E�����j ��XG��6Cf��i��������_�]���nk��j��� �^�Y���C��<����^[=���%�{���h���/��W�Q�N���g�����4Gl{d�f9n;\+����8�*�E�5��?*;��iu�A��CP<cS���K�V�=A���zQ�-<�Ϳk�\�T������{�Q���H�T[�vK|a`8�)�a{� �b���),By�.���
-���yQ�M|;m�T:��:�B���-��fM.�ۖQ&���к;�܈5ʫ�4���9z+�B���kO�YM���FL&�ѱ��j��k�h�*y�{%�ua��n|0Z�aeP�N���U��� ĩ��U7U��s\Z�t� �K���eǁc��B��������S}����䠯b7���f�j����"�ߒp�~tZJ��2ݡ�MҀ�?E=,kԅ���<o���sׁ���N����j1���w@�{3�	��9R�\�����s��Y�ɟJ@�.��ͽa�׌�W<���J=���d(�F��Uo����_�3+�aq�ØWKa��0�Q~��i�<�-���LX��Y���M��X��V	��qZ�����ht�d��r?>��rY'H��U�s	{��t��vSm��^ۅiuZhD���I&?+�6�h{�d��ڵ�o�C7�p����d4�,��n�>3&|�~��H��3G�.c�`��|iG�ZW�1/x�~>	�R��*`�[�.`E��6mTR�BP9��m�.��� k^9��]��0��|���9�Ь��U��8A�i�r��fk�Ztc�5sS>=:�ЕT�9��?w�7A�Y����*���ܣP@Nn��,�:���3��h�`p�p���7$��Y���ئԐv7ѽ܂��|~�P�Fp��V��(@&N$���^�� �s���>���^?6'?�Ȯ%��2�b�>�Z1�N��EӍ����=!�%���Y�V��5�|C�|)S)������sV��4S�
?'��޴hI;g��1����Y ��)f)6{JZ��FE��l^� �S�����s`�O��N�^M��"��5�$�$�te��6s�Ϭ�)V,(?���"3��xt�N�� �ra�x�+_�H�,,���\����$�c����U���I�����w���ď��Suh- Q��A_������D>��,�����\8:�ߛx�{U���3�y��F;?�u�6���O��'���>��c�R�Q��C/�����b�6�P>�Z�n^�Ѥ�'�?�R[8̈(��C�>'�>d�|�
6]��L�����e�sG����O��b�1wVo�֣M!C�<��9�?��]�ʤ��U6��n*N�m�%3�)ӀP�V�����s6��/2��E��J���]��)��mq��l	������cfil��	�Xq �����KC��oZ{�u��dz��dy��9^@�ᢹs�;�Xl�� ��F�XD�7TR��̝5t��E�	�Zk�z�=��EU�¶Ӟ�~�K����%�
z"�s|�/�'�}ܰ��*3)Tu�e-
��]��|��\q}S>�UGy1pE���h��m��Ƈ����V2Vѡ:���c�, ��7�Ԏr"�j��l�ҏ+��W̹-G�쌯n���w����$�{�W[p{�d�z\[R*JJ�P>y�B��V����z����"J��:{�U�+�<b��I�{�L��l:+����w8��qp�^���<��n٦ϯ��K�f{g��w��[52F��^Ŕ�����Sǭ��-9o��ё8�EDg/E�q1B�G;��[�o�ר���8&˭ِ_E���
�._�&)_n\n��V.dF��ZV�z�U�#�H9�`=�<���S��rYx��w�w�����JG�����ﶖ���_Fj'��|���݊d{H�x�����`�j�'ί'�49G�2��Y��W�$��6'�"I��0`h��Iҿ]m���IE�7����ܒ���ᘢ��!Q!䌮�zG��i����֝�O�=6r����a�!/T���7S�I���b���O8��nvRҕƆ�af�X`�� �YK5����ؓp#A�N�'�0jC����
�2�6���'�?f�=����-gUTns�Y>,&���	0��c�<?�]԰�c6�j���EY���"?���;�B�Q������z�x�>)6w$�� ���7�w��� D@L�Z��{�9}L��ߔqZΙ=�n�7Kt}�ɑ��,�u�w����V?��=��܆�܌�#�+�I<�-b1uT�ۯ�_����LSU�i��w6�0.e���!�8�2Η/~=�0���f�9�����x/��C��`t<�3}�[v�,����(������=�b�.OJ����u���e�H����6ZĮv�����s�-�ud���?%��[��W;*�)�A?�r��X5�O�r�Pf�񴮦����;��y[��<�A|�a���2�UxQ1���cuG�_�.{AFdBc�w�,��e~�bT�̸�s���G� 1�}#��97�7&���k����'��Jz�;.s��BX-ĘX����=u������3z��9Ӹ�.p�����qx��G��P�Xe��zܘUK���Q,g�5��J'���i�}�ro�|��O��@���جU����s�!R��'�M�m���j`�еr���{��;�`�Ȥo�����}���w(���X���Ɓ���3)oE��5�1�8�2��	��֧}~sW�P}�lUہa(��Ժ��ެ��V�+�"o�ZHզ�R��a�
Ù���L���1�}�� =@¿�!ȥ�;��u�[!��1uB����0K�B���8���E��:��ߵߔ�S9��'eĬ+�:�R��b�q�>G���
��~����l/l^�u[�G3�Y��`����/OL)x-0��p$qLY�±
cmPcm&.ʷdM��U���G��x�j�F���T�&�O��d�*
q,ٱ��~!��
�	�@8�t��<)��4I���������8m�hmo��N	��E�mmt���Ru� �֐��8L
���#5c�K��8�D����X�h�"��
o�چ� PJ��9���-h�����DJ��|�a:4�	�X)�F�����1�rj���a4��ߢ ��"�ϡӊL������|G?�@��������)�J=@3�+�1��t>d�A΀��R?��!j�����R�'E	�SW��I�Z>�ˇ��p+HG��x�S�s�Jw�+7SN��A"�N��MI�S�8�F"����� �����&~�%N��-6:1D`t���3-n��߸n	́6�l�k�|=W´�!��R
>)1��M6dQ
r#[#fSQ~�?��mʵuB�q$�F�j�l��iM���$Z�ݍЪ��kAc�8�68uH6��4%"��IAJ`
�ç����˭�8�hN�8�F�u	�K�ç��श'D���������}C"CV�6B�M��@���F�)�PS%ҩa�t��eŔޮk���.����*�CY�ᦜ@4)�*'0qQ+
���Պ��7��6N�F�Fs�@����V��L�#r�BB����~�U�_�r��b/��F��.�YH���X��	U=A��R!��i"���Z���>ۥJ�*��)䓍�9�8M!����cZ/M��Q֌�E�|��	��Ɋ�9�uR�����"�\j�i*e6*D�UB6E�p,��2��o��|����d�k�*�q��X�Nf���
�pSY����݌S^�%K*�R��a	�L��h�!�#$�)�h��JO��oJ�XJN�����U:��Qtq攃G�����D�)�����YR�MƧP&?)��|Q���J$�(t����O�%.Wnj4"e��8>Q���v8����$M:�(�[�BL�y���z�B\F��5�Ԓ�B�Y�J���75�!~����[6󠌖0}-�:�.�R�;�ݳ���������~tquy�k]���(�>�u��;��l�e�Щ��g����³���	���>���G�~s]��T������c���D��������~��/?�9�;q���O>�����������́�s�z�Юܿ{�����.�>�����yT�O?ޝ��?����ӷ�߼������˛��oo}����=��Ú���Z>\ܭ��^�#�����W{��U 7����/����{!�3��iNǨ*Ʀ�I�r�l�MU�.րlo85�aj�U���G;�����0��ڃ+mۍ@�Uѕ�п���vG"�*�h�y���O�>����l'��+�)�Ȗ/do�-�S��w��� ��PT�,L
h��~�V�+m-B���0oѠ�BA
�{JRԂ{�L���w��O���)�ڠ,])N�&�&Ј ���������|��G]���6J���G	4&
�'�A�B��#j6���?o�R( � �)�Vp��Qb�!��YbQ>>B���q��!��,��D36�M )�Avp;m�C�g 3%n7��{B̒M5�ZBՑ��pQx���{��F�m)D�4K1�d|����"}n�9�ME�u�(��h�JG��(DT��;��5k)]
��ֶ���UdpH�*|lT3��Z:v�c��HP�	�!rŴ� �jj�� �2"���45���S!)9pSS��X�"qE�wt�:thG�&%��?����׿�5~���H_��)?e{d�(P���̚��1sN@�;�r�.�*nJ�U4��^4���L�jm������v�)8�B|8>&� ���V8���7H�Z"�DZL>�;u��a!{�7ֆ(����T�o�`:F���X%���W��D�MG��1)�iD�LH!Hѿ�Ѵj�jވ� �� ���9D8h�PsgD�D)uXM+�Tv7e�Is0mi���Ɵ�QÓ�_��:�M����j��N�B�����i�WqVQ�)�\~�T?p
c���l
.df��)�\>��-B���R�^kc�[o	��U�2|�x>-�'A��6SQV��Y=��ob��THEf�@]���G��)��^T)W���#��bZ?��9*TE4U�$�R����غ�&ɮ��}��� �)$C@�R�����~��׫�FP���2( �[_�����ߝ,����Ƚr�����:�Ug�*2���\�B��|R��I�|���E���ng��0'��bOdLu�@�q�̥o#qP9O�����4�R��e!�jL��h�F=# K7��NҊTqsq=��v������$J��gd;p:���<B�(
Ԫ��ܑJM�P
43�o�����[����R���Z#qC�i�Y����-��ٞ?�H�B�����28>�(�c[ү�1�8�R/ڴS��9�+�VS�@V��|�B�Yh/r�mD9~�Q���	I7�EΐY�9��G- �Nug�>A��[T�D������j�Z�Ǐl�hR��U����I���"��s>�!~u�DHmh%LY�h��i�����m!%�3$�,f�����Q�b�h�Y3s�T?���&��GH	�D�;[�	d��	�zG
B�>M�݀��OJ��J�(
O|^?�BFR�եPj��J�H���K��.�2�N���8���P�S&��o���4��VQ�|����%�I'�l�c����^?���H"�8 ���N88l�8qtߨ��Y��!%"��d��;?�9RRXe��0�8�I�w�L��@�˕R�Z�!8�ɗ�c�9pVQT��S��xj��D�����9�6R�&%�l��
ωY�t
ё)�����\�#b�U=2�(�T��'��)��%����/Q��8����l4cSLS��	���69X	H��P[*�_z�D,��9�Q�-�d�X)hE�����R��mdM�iE���,�u t�'�B� eљ�E�#��o-�DF��k`����@(!5#}��-���C���U��R�s�-S���Q�O�S�S��
M'Z�$;`%��PHm�ت��䰢�p�zˇsB"75`����0 �+r>)�*m�)��'B�B��Eƥ�)q���Y-����j�T���x�L�d�qR�m:ǈ#jde!z��aH�r�P(�N�)'�|��rp~�8�p�B
y��п�8n*WbW<����ED��^rD�8^z�V!S��!����OV���.A�ڐ5�+y;.��K�С�o4�R��w�y5�O/ {WWC��.}�e�3�us���L_z�>�t�4���9�sڙc�(a\�^p���T��ߝ|�㻯�uS��L�+����!K��{�~�ҧ*�w>[�8�y���E̻���l]1/���}ODҼ�����g>��n���ޟ,w>���za{��Ov�٫�U�����l�a��xg��]��������b�;�����?��\7Q|%���{��oϮ�qr���nŞ�.�����g���c�~������	���n�^^��_��{��8��8۽��}}�zs�ܟ����úJ��7��7��vFϐ�r8_3��֑�N |2�Bk��_�F������@-�RL9��0�BKqqv	1��8?�B� �#���	�NDMSHĘ�X~N�Q&H�B��C�����+$� ��Iy� �!�ù��ǎޘ(�QiU�h���(tQT_n�z$��C�,�Ø_�F���K�.=@�q�}��0�W=�r8�[E�B�C��M��U������C�~�([�a2���1��0!�0��Sf�D*���s��_���-��ddzv��z��\<==�X
�$�6ʅ4V�/(�)r���a� �Yj)q"�;��Ǌ$V����Ȣڞ'���i:�؍j�P:YS����Ch"HL�Q�b�D��@�|��'>����  �[rMA��G
�Ǒ��#2�ؑ�L�Z�ǈ,dj�@�t]]�-��F���N"��=����1!��J�tl}�tg�c�h��KT<$Ӷ#if�(VG���Wr6H\됤�)��2&�h*�fT:P	!����j�����_����Jd&���[�)d@�����L���#�D�'�KL�c���A���Z��@ʪ�2:z��'�B��2M-�T-o�R�n�=���>Y�R��B�� |�R��(�8������
�	�DHK��W+g{��'n��r��� �V���Ԁ���z�%��*F�r
�q,ު�1>�������G�Iq05�15��F ~�� ��!�ݖY"�q�/=`
@4
F~�4͠U��)C05ζ�2Oێ���~�W⤒U�J9���H����H�[!>b��	�r�M"��ȁ6���ah�ւ���h<�K�ض����4�PKre�PQ!��	$�tB�6)d��M�%�1�ČS��ѭg�����*M��\"LeI���ad;Q�KЕ�i
�8�sd����5��OHk��R]�D�	1�(eVE�W�+ea�iju8)l���=�;FF��ݮs�GnC��nmz��lQ�rYug3�Ĉ�%��A��*�3\u�F��u�a�B�ҭ�hC0�,�z��׆1\Ì �I����Y!td�0�L��W��"$�o��֏�9(�TH��-�yh�bi������j�Hs:�
D�a
Ն��M�8t8BL��i�4*AV�tƜ��=�ɧ����
K��S���W�q�|;�D2�$V������/�9�s��7��^S#��B�~R�D��2%R���RF�?��-ZEg)�A"�I����t^�8p{��T:35Abۨ�[�b�r�8�䛾���\��x��A�L{|�h�Yh��YHb"|�%V��l�>b9��:�o'z��Y���h���T��R� ��K(�c	ӡh��Y"٨4�(K�6��H��������c�F4��i�#[��$��IA�i�D�(t���
�
>Z�j����0��ڍ�h����# �F�Z
U��:RU�D��!�8�N"�pc:9Dp 4����id"���Mu�T"äf���k�X��@�2֪�Y�)G!)�G�s^�!7��Hlcq��9���[ )dm'艌`�hD��>#�+lD�ԕ\N�8
�r�U"��H�F4���BUB�
ČSz4 S���):�B�<M�Ĥ�����0����=�[�����f��J��8��*j���STV�F&�%WW���!GT]L�e�R�4"�d�
D���vS!�#"��e��/Q
G8�����[�>�TV�`�5	)2|)#;~Q{R�t~�|vX(��E��Ro�	�����˂7���ut�\���h�	
�-�}(2:9Ʋ��N�̺�j���������r���}-�r@��h�p8FH`�|!S�h�I��,�Z2��b}����(ĸe�c�o�������N���H�I� �Ռ�4&�TkIS�>5
��&M�Y��D����CC&2���d��7��̞�F�JV
�#K���i���%������=H/DqV��S3eLfQ|W�����m��yJ'B1�ʈF�(�5�������"�n�m���@+}����n�1%ee��:ů1�d�����"=��;z8v��IJh�O;w~q~t�~����٤nO�N��}2�g8}:s=^4~r�{8���<�x<����ˇ���ㇷ�;�)�ַ����w�K������r��A����oJ�mO|D��&��Cz����<��u��>�<����N��!���ӝ�]���[�'�pw����s?�s�p����ۛ������ɝ�н?Q`�;9�>�B���ѝ���}���]��'W����8:�Zߙ�9�z���ޭ\�8�caہ�0��x���O�:jO�9��!���Ǐ�>�:���tB�	7"gdq��=����4��Vݸ�'��=�(�O�)���<��w� ô��^}o�;j+U�����B=@L�{D 9��e~��罽�F��%*�	OD��J�D�'pS�_>�3L�����M�PޛK�8�.K�\N|82��\0��6�Ti>��4����*MG�(�Ėǈ��	��e��&�O���#�HY�xӚ���P:�ե ˔>�n�2�C&EYKt�)b��&�U"��Ԓ�p��ko|�d�[��D���	���r���A�)�>+�	�ǋ-    IDAT$'�8��G6�	>�D����OV��N-Q�p�FY�)��X�HM�m�r-�����F��?�᧟~��'��#HG9!L��iء�=��h:D`��a�g��TZW�Z�!·:�����%�7�F��c-7���!�kLm��>"�Kg�~Y�__���Gz���z��tr��OB|`�dlU���E��K�:�oa���#q����Zo;���@S��W7~�����������o_���_�}ـ�ǥ�Nb����݀��zT�z�Z�o���~᯾���g�޹��D��I�����^��m���GO�A�xt�DF��:9D��B,��o�2q��3_t�|ъv*ش6P9��8�p4�p��S@�[���D�=��QRnb'�Ď�����]omN� �aZW�k�g)s ���o-%���)22
�F������:b�B)��˷
��VaL�Ð����� Ghr��"��T�@TIޔ����Rn|��F����C�	�YW@V�O�XkPe���ޜuF>������p�i+�m�1��t�~�!r1!,c��X9�z�Ж�,�he�$hTEu�@V��E�4� |c�Q
���,��e!�!�zj�T!�P%�)F��(�i:ądq<xR�
��� �t7��t҈`��>�hQ"��(�NB4��h�\]I��W)8p��\a�C�T���7�u�֪K�K��~�;
����t�5�E^�8F��у�=W?�����J�Ϥ��I��L�Z|r���gY���2*-�����D)9M��җ؞�֟R�_�r��֩� A�6�rV(8��`�1~K�c�t��Q��@3���,FPV]q�;'��şVq�R�Չ�=jL.||S>D�5�΅(0Ӝ�!�JpdM�Sz�9F�|����Tm�1k��*���Њ���Q�V-Y�II���9�MIE�8���9&��)'~S4����v$����u�NW��4f�{� �Ҭ�P��r�T�NR��	�ǝQ.�!����8u�'� �X
?�8��09ِ)�������p��m�)fk�Gn�s��`!h5�
��B8���hj���P�9~SL�Ӂ0њT�x���A�+c��b2H�F`>S����a�8R,�Ƀ����M[,&��%�u%3�>sNH���h�D�5�b*E����߶3|`�h���
1!>PT��ܜ#�ZB���'����9�˵'8|!�d�Hґ�������JH�"��	�7`��d�#0SQ&�	18���GKD���!����@����P���"Y�J�eǩ���IA�@�nF�,4��N"�9d��Mbxk�n-��G��!3e��I'��\�L�c�ǯhe�AbRί����� "@L�,EMC�n𤌇:heUN.�3}�"AT%عǡ#w�q�ф�ҍ���o
'�,��*������tUf�bMį\;Y��q� �ei���1!�t��br6�Ǔ�C)E4|�?d���lBj�)� 1MHW����d�)E�BE�0���-3��gKZ�bz �D��ǳ�rS�`�����H��4E�
)��B�O:)�DH���9)�C��8�D�� E���d�#C�3DJS8��c�yen��#��q�-�xE�|yt8�C�Z}�s��l�@:��u�"��K����t�r�s5��rR�.�M���V{���@V�ܖP�)�����ؤ��SVd �!��z�6'U}
1`u)�uY�#QT��������k���$�buR��^�Q��#��G`�0Q|�|f�Rf�hӁ�ӇH�a}�毫�������=>fZ�w�3�!I��'"�n����w^n��R7\��C�ue-R�e��S��v+%���:=�~v���v'�۰�/�Ο�%��ս���9KO.no���1�gݥt+��]��L70�o��y��=D7�_]�0�[]���]׎��G>��pw��u��Sqrzsoin��)K_C�탡�[]��y�q�?����>.���N� ����c/��ןdׯ_�_}�����������W��k���7��zr��f����r�����M�Pon.�~u�՛���ś�g����Z;�ku��|�K�}ӪM�<4���W�㰵�|A��s�mG�ȷ��\��}�N��&�l���D��!@�	LC�������t-ş�S%�N����&��A@kQ�s���R��9��� �h�8�ɒ����ٽ�b���������b�_���e�?�9�ۨ�*�����Bl�LY�	�V�L��./W!���-�C���hS�8�v|�jZ�8ܔ��;t���W+�qWE�ͪ��U���F���#ΏI$A\Ϧ|�MH�H��U�K։ѪU�k[9>�O�[Un\}�;�	4:���9r�tT1BLCf�R���L�t��jn��r#�Xu� ��X�D�ҥtbp��r0#;:iz_�3�fGGQL��1�sD�~j���~�ӟ~��G��jO�ĲL�'�@��d�k���
�׼����ڬI�'q��ђIu���[�#��d��?���)+JD�[Z|d�U�˿���~�����g?[ߒ�i]�<T:<����r�L �TO�s�������K�7�L�|�C�����q�U?���/+���'�~,��3���������z]87�g#O�:�僋d�n��..���8YW����3Ϛ�'������3'g�}q����M�ޥ��g���pl�u9���|�ű�Y�&M�8�M-�cㄈ G`����fut���혙��ޞj^t
u~�2= ���"�%F�BZ#�)x� pNR�H�3�@� �@>����4����۴�ˍodU1� �����ÆϩVk"�#:xlj��\>k�j���U�����)9Y���ߢфr�:/�W�(���lʑ��tm���B�f�'��?p>�'b��/j�zN�Mn >�%�)����g�4���&��U!�tD�������*��̹-Znd����k�:�C2����R�*�f|#�[#~H}����H�F���L�u+h"��j)��Ei� �I������1R��W<!����O��p�
MK��.��='�����h-�ޮ?r�8e�azF4"��lՍ��&"�YC��yS�)x��X8��#(��/z�B�iO��-���K?���|Bl{���U�) 脣"��m:��ւ9Gh�[�4-D�_}�>F�*�J٨O�>N����3=�a��m���%F&�޳hՅ�<.|�J���h|��`� �@Qfϛ�Z&��)k��fZ"U�*�<E��E.j
o�p��ү�8E�
���p�6�*1�@N���w��M�&I5�I�Ρ�i
�P�>�;L�hSN:ٶev� �щ'2�*��@�q�ѤKa!c�"�X�1KG:f4�@>B����{�p��&�S'FV.��Rc�:���)d�#��SΑ;�t� ���O!r�p�BCS�t�PӢ�҅�t�����"�\�K	�`Q@U�ʘ�
A#S�褛V���_|S�����UQ4�4#W�άQ��Ƅ�/���L���磆�� �Z5?��z#�Y?@<��d	
��)|�m��Xϣ��đ�f@��~6�Zl�FYE���
���d*Qf�!������T��)����38�BE�[`�1�����eh���%�V�E�l�9�`Q�'Z�SE`���8$P���D54��L9}����V���o��H��I��!�d���pBү�h
����jҴ�r�����8@Q���@c�8	B8@��iX��Sb�����1u�YS��\�飉��)ā���B�%�[m��H��(_9!S �dq���sƇ�4K!���5�t�d��Dn�,�����S���Q��)��������&G�D��p!�P�]{Õ��hS�%7b�m&���d����|!|����7MgJC�VQVk7���J�C`5��2�!�O�ooL��i"�RL󍬃X�6�Ek�a8����%j��
"
QG�t�/���)Y�O
>>�h`�� LӨD��j')�pv�Wژ���6Y"��ր36���|�S0B���ˢ�Ʈ7YB��/}|��Bk39ޠ3����V��qA#؆�Qc�(V"�S�H�`I��
)�,��H�g
I�#%&"Wo�уt�n�l+�v�Nζ��W�g0�_Կ�|��>ƩogU����n�[�CF��O6>�~�ᇣ���o�u��=�:Ո]�޿�^?t���\�~�җ��*�<�T��M�/��;�����AC��y�_���7�7c���;_{��c���������;�Gn������]W?.�>�*��8~
[���?�ܽ��u����-N_M��W�޿|�;;v#vw����;�~<��k��^}���/�n^߽ݹ��sS���˫W/�N�=�νo�ݻWz���G_\]�y8zsz���ұ��u�S�O�n�����|غýuuh����t��������q2��h>=�97:1�9k���H�X-����G:��D�fd���F`���X�V����3Ȩ��2S�>E9��� Y���֋)4|�������{�D�C�2K!±�޾��[�F��M�h� �J�����*z�3�jY2Du�2��釃l�S��ޜ�z�B�G�>˅����W�ڙ.kږ��$"˒����I�D�H�qH���V�F6}���h7�%J��)N�@�S�C(O���D��j�׏j7� �Z,MY�	!0Ȁ�r��'Y�J{�?�i��M�qD15 dE����z�MvN �5o��j%U��Iq:lY����E˭����o��w������$��N���-C��ק�>��|LGGVK�O�8�ŜG��e�O�(ı�h8��zl�=��=� �tNoi��O�~��_����1�$]9텎+I]����ï��kWHk**7���8�(�4_:�u��<ZT�O|<|��'�W�k��//����s��<?�]���ĔK������s�4/�{��g��c�'�������>pi�j��w���ˋ�`Ӹw��S	��i��GJ3�-6R`|#����X����
>�Q�`�0!����sB�'������r��k3E�=��l`*���iDV.Ad>���5 $+!f!x��C�sb�Xz�FS`��וB�zK�J_
C'#�gMq8:�!:č82���,�ǉ����1���R�|Ym��ę�e���B��3�L�Y�;��΃�����������ӌ(�>�h�6=ā#(�T4N�9�����h����#`���j��i�YT�L��i�#�)��o'�9dj��^�L�)�	����s�[��MD!���r[f��)>}�|�0mWg[���g8M�kL'��]F*qW�\d�8F�F
B#BYԕ*>Ĕ>�>�&�f馔����#�!x���5i�)��u�t�B�M͞Jѐ�	*�!��S>2��i]�ᖃ#��t(��!bu�MUa�|#sxE͌�� �]lY倥t�j���RN	S�a���f�Ę����)���6V��������(K��̑������׿��f&d[*�cO����g[$DJ9x �e׏�SG�B)�s�8��ą����W��Xh*TT:G"'M���tx�J~�~
!�7��|�)'�*����}�%�?��;4R8�q� $"�2���q*m4����qDs��<��.PԒ-�)��\oȥV��Yd��`����C��,7e8�!%��(�أL'р�D�֞p�t�B<X<
�!���**�8BS:N�P:P�?m�d��i��@c�⫨�;��X�IQ+��4et�&����b��b|#���7�B�N��� 2���S2�F-�>��n��'G>N�B�9�S"�P�?�a�A,mH�4����['IA�,|Sc�3��/[A�`��v�NYP
Z����F����$[�;�q �R@6-�X] �՛^��R0�EUD� LK�w8��tfZ���jg`>p���FEٜ�8�J��Y�m�ۚio9����g���R�v�eB:ĢI%R��i�8����
���wJ ���J�4�J)�h:��҃Px��dg��0QH:F������Y���îLC��8!�-�q2�Lx!=��A9Rh�B�	LĘ��,.��1���I�Dۥ��)�pfg(���\��C9�qJ�q�V�h�8�E���V��$��WQ��h��8G�|`�B��YU��D����|��b��[d��*9\�$���OsKzԟ*@�U����8E��FE�m��� �v�R3�Վ�/���d�`Hk�,*q	eU&7f�hEB�MkҔ�8�v�rY�1P��Jh �Ñ�ZBO�P)B=��||#"!�Y�Ԣ�	��5҇��r���v%�C'A2��2�t"㴄���3��F��Z rǀ|Q���P�ü�l:{S
�cD3"X�(��Zd�+Zo��M�S�~�=��=��%E��%��L�hUR�E�T����-M"$|�6p�"�@M�RVXd`|�]o`�˧�ߚ��������-��ܼ���v�Y���%�tM��M>f��vs�r��FUC�����J���R>�~�r}��ɱ~/s�`����a}z��ϵp����ѽ_����;�������8{qy��{R�G>��3����*ޟ��IýE7B]c֞��a�I�>ח������z/��h�~`�F����������W��^o���ԧ�<��?�_}zt���ڿ}�cj/���}�r����7�w�~���Z���stΝ�ݑ����߽ܟ]�x���A����/�u&{�r�E5��l���O�������ps�yO
k��cB�,Z盱w9�u� L�ME��l�n�&:����B$ͭ��cgħD��+��%��wԌ
a&8)�_CHvV:���p����+Rt�ljuV�#T���֧���N-~R%�~�L#_�~*�V����䢅R��X�ߛ3���`�=7ut�N��4��E� B�|jp
��U�/
���B��k���� ��8RD�����ҫ�é%�5R��2�)Ԍ\�,���6D�b�7���Z���LKA��_�OS�*�j�Ttʥo�	��Q���B~ʁ���1��'���r��|�=7�1|k75:��������7 Eg�e�14�����χ(�ˀ�?���W����wn��R(0��9�S��?��@��adN}ү[�3�O_��zS]
��Z�*=T{��U�Ҽ���\|Y�oe獪'Zљ|1	@Һ�W��!F�L���[L}���Q����D��2ᛰ�+���{�Ŀ+��N.����r��_�_��l=~�|w�[�O��\�/�ۍ�Zռ��Ϧ|����	������o�������?����K�_~����ׯ��3����u�����}Z�Pk���J!�QT�+r	hgZ{�F3�`��d}R2�E�ЦUE(��M9���:K����v�\=Kw���҆�0рS&'�����V4r��UEL�)�W(d{���kF��af�Y�h�qL��IP���Q���>Y|�����Q��4U�0��� Zb`�n��r!ԘЌ��۷h)/��g�I4�6-�c�����B�XzNd>g�D4l�������F|��n�X~�p����-*4N)���Lk�cV7�*��D?N|!S:)TŴ=1��l����M�)�� w�lQ����l�_�M�a2@
���T$�pD;M���B�*���c�C��z9��
�p�IpS�(!���0�m�SDz��qcLn�����L�9&}�N6��q����4�TW�-��3���뿺�餲(O����Kz��D�3�5F-)>�d��9%�n��t�뙃_h�Z��'`%�EMgMC�����sʕ�U�@#��,!� �Xi gړH�6�S!������ڐ��Y#��Z�do-���<ħ�0}?���*�;Lhl:ć��gC�]:ZQ�@R�1���(Qx��҉�SZ
�DE��Ke۟8h�p���DNE�ٖ����I�!��O����1�&�1+w�q
q��j�DMYk��,qF�R�aF����.4��Q���c�:S0�qv��#j��Q3
ѩ�ʡ�[�pS�(ٚ1e҅p��(<�d ���    IDAT�l�%X
F>+���l	���#T��Ô��X)�19j�&�yE�7�[�r�Y/�TBL3�!��D��& T�D�YQE#�E�n��������r��O�h��+�4�,����ÑY]�j-����!8Es��0$��tHU�L�\K�dìC�h��K���h�@����Moq�A�i"�r�vn�NhrM9M�"N��Ɋ���[bY���j�P�i�&��J9��h!Vʙ,��(¤כ�,�)�bF�mĄ�?#Α.QѺV���#��b�1ũn#��9U�iN]����t8F~")LR����i
q�%4�L���Y��h��ڟ�=!�(%�j�v�ڷN!)8%�=�J$�܀���UQV���_�1�����x�Mn����]Q�g��L�,�,C�O�V!�A4�)T.0�B�q��L�h��+������HRR�1�����#T>"��4� /Ti~��pﬨ�rU�!�ycS�њ"L'�Fj�w�d�a	>ӹ�3�R����Z�4�#)p�Nʥ ��!�(��[�8���W�jф�sҴL�����͘�9��>n#��\Lmh̸JnE#Pp���V(_($���6��F�u��ů�FQ�X���օ_�ȵ>Ρ_K��D)e%R�F=HO�Ј�C��L�n��NM9/U�U
��ņ�Tz[ѵH�DL�$V��j 'e�{h��[�N���ԀUA!A��22J�/����U��{e���n���ԧ$E�/���?{𧻓�����g;�yrq���ǧH��\euU�D}J_��)���9����O��WG��(M��<l�k5�vk���>���*��"�^�����X�o=�� �{�������_�8��[^����_��͗�n�|�iz�{m�Wq�f��^O�[l�f> �p��8��՛[����S�Y�����,�^_]?{�����y{s��例&7�n-�����o��[:7>�s���7��f���z��{ѷ~�S�������Û�5�{��}y����+g5�wA��s�:��1�帯�{:�{�u�u�i�q�y�,~�Mc�p�!���hE��%ӄ��	fJ�HA(��W�}(�[%��`�tRq�����?��)L8�"|;�kß.h��S�R"��D9B�����7҇(*Ĵ���L"���]�Qc����cu6�Q0B�"#�}����jc��/�4`ǀ針%*Z�Y֊L:�q�R���z���0}=��b��oL��})��[�֞�w�� ���T	u�:" �.K._�i�(����)&5����hF~���#�B�)�+S%�`K���*�%n�a�����S��8�R�1>+�)7Nx��Ѫ8|:BՊ#���5"Hg��cuh���v�ɯ1���G����禦[f��+D-�D�M�lc]~�����tYpn;
>���� ��41SPq�pֵ������*q����(�*���%��K�gS4��A{󆧐7����h�j"����?�ɻ��3M�{�kG���b2���C�bU���cF!>>C0]*�q}0���FYZ)+�3�킻N(��yt<x��M���g�>��������7�����pw�_�ܝ_x�7>�)�s��琗_����>��_|�������L��-�~��P]���|���o ��]_��>,��?�8:GӤ��6��Qak�ە.���e�N�o3�Q�H���ʱ�@YD�����mC�Utt!��'E�Xos88����������L�%������)��J'%���̔!S65�G�#D���;�ȉ�#W�)�&�f"�3M��!��"W7��)�Q�,����b�cR�#�~=M$Q>�6���s0��H4 =@¿uE�FVo��s:��R"s4��\>B"M�Ne)7�w�Ԍ�]�����CG>�c��dqZ�K����$�	th8�PA��C8q���T���I�#�o�!�������N`
��eVהC> �0Eq�&�PÜ��XҌ��sYVO!��ʡ!���ҵ���E0%ȧ�NȪt���Ğ��\�iT���TA�C���0�cB� �I�m�!��I�?�1ʅ�ʹ��g8?e
m��,�4U������f�p�"+j!���ާ�~�_!��K'���u/��t�ŷ�жr�O���ב���8GP!"h�J?Ȗ���'��nu֫Î5A4>�����T(����Ӟ{bEzC��-�@��R�#HA���D��\K��C)m�tQS��aruN�2EK�� H��2N���b:N!S��C�]B�A�p��C*g�XZ���C*j��Y"M��)��8찥�6��P%��	\i�Q6N	:���aE��pH_==�d�p�@���
Ajrt��ls��X����
���8uMG�si(���[���&������hʪ����ktLei����/7�q ���|Rn���S(��e�SB����K�f������/�g��1~�B)k�}>�_"���|Y|8�8p%J��@�9�< >G�s")�V���Β�s
�áfʐ��B|�,?�����}��"@�D���+)Υ��f��x��d#�i�t�9�SH�� ��~�&T�B���2j�0���k�uGj�2 ?Dbm�Pj�mD��7ʅU�N#���F��ڥ�(-Ģ�d�N-!]����[K��qD��z�2'[::��g��G�w�(�LM�q�$��O<Mx�2��w�M�����)K�So��L!-0�R���q����&�~���#T�N`��*�h���
�M��`,=�F���6*Z>�����ڊr��P��6��h�yc{.d��1��z����s��[Q#NN�^o���B��+��=!�� Bh!�,�MTVӪ�V4eS8�!�/��S���m���CY!:E��Z'U.|��)HLd�D�|`HδQ�i������f�@�CY�\c�_���IL�V��O��^8 ˚�� _��Ӊ�4/Z.�n�w��TN.P'�g����?�Ks�|�9c%���B�QVk�j���iu�^���cDKj�I��u�KhO�J�/��=��mu�QѢm�i�Y��t��k|�u"��p� p��eEh�"�P�HE��-��X/f�u���Ȼ����W���ɣ�g����_��y��/_߸?���nW��53��YKq}��2a���^4˳㋰>��c��8�;?��!�Y�����z,���[���S�X9�I������f=|��͟����]·{_p�K��m������zCx��������]�]���i�uTv����>��ߜ�����|����/��o'���ݼ;;ٝ�c���q�׍˵�o4_������{-p{��6���|�z����/�#_�{�W:o��=��󨍲k6��B��<|V�� �4ġqdM<�X����9���
P	Ɓxu��D|8��ߍ
7Ш�����v�a]g`|�NKS�-�T"�A�T1'|��)@��qZWj[��!<�*�|��F+��m���h�n��0�[<M� \�~J� �qRF���&�G��G �V8]�h�$,:�\%�j[�Ð{�%e}����~��z���<���0#����(&�MTS)M�z�pX��[�����SR�3��bl�8mE�P(G���JC�"Αk�9������j�5i��C�Ҕ�����)0N8�n��F�·l�[uK�P�!���HA��Jg	�J�{m#+�T6���L��3��!H5un��Y�=���;��U�@��.��o��!��-Y��ӟ��t}pjR	YԬ� �v ��\��*�]E��]��7�b�K
�g
VM�C����-&|u�t��xC�T['�ou����%�ijD"wVYg�F*p���8!��d�B#2�gR����r��4�պ'����Z�9�"�|��Ov܃���������߿�|���������{qq�io��ꏯ_~�g_�~����w{_�w�)�����5
Ԝ�W�7�.=<�X��/~�6�������?���Z��v� m�hξ;��5���+ۢl�#�rL��q2�t <�pH!!mH[�VH�������*R���\x��#A"�`R�����t(�Y4	9�![]䪛42�'��8Ch
�秬4D.Z-՞B�!�ǔ�H��(���O�DH�O9�՞��(W�`�I�9��j����g)�̴�V�/JvJ $aBE��|��(�񍻆8i:v��-�T����)��W�������+��>��B!��V��b�U�f,kR8UAc��HO�\���C3��ex�|
9�e��P��P&8-�d��ϔ��J�K��U��s���F�\H����袏)�r����P��\�j��+y���傏�B�r�(�@Q�E׫��]�D)�$���f����G���.��.�:�W�H�U�<�cʗHME�T1�lʑB���c�A�i4e|)�V�^����-}:
�y�z}��v�4��ܻT�Q���]_c~z|�f�EKS��'��-��9U3[�*��jjg ���/\����tY�z���h��<�($q����X�8����CL�Q�9� m5�����t���Ȩ�:O�r&�V]�8>f�|�F*q||�d�%N@�	1�J��������+�bR(�4�h���2��ˢ��#�N:�m�g:����!S�#J������&��B#�3)�e	mJk+$B������HGc�|!�HY�Q�y����婋Pn͘V�Ϊ�t��\.��I^W�i���kL�Qe�_8>)RD�7��!�eU��4~�)���A�@�E=x��[B����L���aR��i�C�q��4U���r�8�!�9'�|x�q�5���yz��̉c�x��4-���[K��J��� hG�H�
�Yo>����f|�� �A0�p6�1g+M�r�85�L�CP�F��E� �ST�a-�(�0˅V��M��@�����4|�Kk�$U!0d�{|DC:�R#�n�>H$���c�(�� Ӵ���F[�`%�"���A�l�4c;�SQ~j��IE�eQ��)4�ҋF0e墑�H�c�a��TV�!�8�I��p#D�1��h�� i�� �˪�Br�p�Haq� �3�i�,㠱A�ES��?#fS��1����9�Cd��Y�H8'Mx�� ��<R� ��rd1��F!7�l�5�p���k))��{����(�c*1�m��D�@
Fv��*�T:�Y��"�r��||����0&5��Y�J7e�O����)�h��%�e�~J���&đY��e�XMB0�[:3�8@N!)-���7r��H`��j�$r��� 56�)��p��
E�y(8{E�m2�zxL�2:�T"�8��G�DN��	/e�.�|`�3�!�6�R�Q9̙�P��M.$*�8=$"GNcc� ]"��Z����WqB-�hՉ�ҩ4�BR���9R�B�U1ʪ��g�p��L�g|�Q��t�i�� Ԥ��Ƽ�����R�t�g$� �����}��W�N_�}�WW�����ھ+�a]�<���%*J�����c��|�q��k���A��6-o����M�gw��#�^���@F��c���Ǻ��P���W����酕��ܻ���8��˫�7�7�=��*�}��d'���߮\�J2w�ۑwG��WH=�b�ks}P�i�<��z-�[�>���j��=����j�ȍ��g/..�=�v�Z^o���v��o��hV�/޽���'~�s���-���o�\�ʬ�7�w�����ٝϨj���קK���l���8|�Vg^�o;�V�Ǒ%Թaʇ�'�w��CMG-����BoA�{�����~ ���+��>�F�@4��t:��O��ٰ������H�(�!X�S�1�3�9�p
�C�[^ƶ��m⑂,]!�Vj��j��$2����,c;LX�1!o.Ie�K�fS�)���C �o�;(�R h���kr���:��7B� �:e�(dOT!�f�"�!k��M��C��2����� ��mR8@�E�.�T;Y?�p#�w��Q�NQG�Y�M0�q��1!�42�
M�b
qG��j,����<x|��U��4�3Yj-(b�8�	GAJ��-=5#�s؈���,Ĥ�E��v�O>�*_�s&Zʍ��pM�ol�g�}�d�o�1j�4;�#�-M��Nm���L����ޥ����oQ���;#�L�/����q,����m�7i[�>{ ���4��/�:�g�RЕ�~�s�R�W	���\�$�4j(��X�>fG8���H�����o�� 3,S��^x'���q���B��M�U��佟������?��?:�x������峓�_���~�����~�;�ݞh�޼���=�;���o�x�yF�/�>|�͋gn�����O���_�������u���_���?���n|�H����m��.;f���h�6|4���nK\��y��Ep���"�O"&}{��q�k�4�`;F3)�tY�`�8��4pS)w��"�|�Im�"�f�j����a5���BJ̈0�hI�"���J�`fqV���?·�s&485��[�G�Qs����&�xyJЈlD�ҒS�W�S�� -m�r9�����R�V�FYL���	�I*5H��(���b���F���,fQG�֥�HAsIl��!�M�?l#��|E'�%�-sBEu[(MS��u�?�EM��O9>`Rub�q����8h$[n[��L88���b��v	�8�u.�H� ��i)�&�h˩4!�sD�?]�q<�c��m�?\��4)��)�/DD�i�s�,~-��1[oG!�t�UgR\p(дFN�5�/��-�ĥ���U��Dk Q!�hس���۔h[\���DWiO��_��~�9ϕГ�'�|��7���?��?��?��N�R��Y�wqs����O��gt-����������!(3돿�D�G?��Ө�7�ݵ8=��O?����>ҏ�JwSSÚd-S-�2��2e��5����'V�l�f�^���i�.�>Y"ь����Bc|�L�F��'�?>��(����u��h��B� 0S)�&��?!`|u��!E����r1s���P�%O�äÙcd:U �FH��Mf�"j���YG9�d��𓂴4���m�qڤB-�r�)p"�Q9u+��7�2��%����R�����?)�|H
M�J�W������đ^�LE)T�	f��OUdq&�el�iJ���oY1�i����!N�C\�Q{��rN%JO���fd	vd����$�\�t�� �N"�Y�r��H�r|#NE;��CZq��4$���đ�O�� �g�Y⦽�ә�6�"%��E!��̴N DL�im���]6!Y:��W"�U�A��v��pb��9<5`:���h={g��[R--A�ZTט>�t�6�mğ�#rY� d�C���B8US3��(MN�E���o��fʔ���~��u�)�$�4�-�m][�Qb��.	a�EU1�)�|�L B�z�����Bx)���S�#���P�|��R�6�H����aEӪ�F+ޢ���L���Ԓ;���
�TH4>�\�ш'�3�pirM۫�t+a��8��SŦ���M�q�oqG�X�tZ>�}�G��)�H��q8;�0IU��ߖB2x4Q���G�Ӵ�gD�Rn��R�i�B`��A�p��sQ�w?}4>+%��逪�C��ƭ�Zo��UT����'�?�8M�#�5��y��1�%p}�1�|��P���lp� F��u��I�88f�q�M�h���������J1�Sp�ԪO
CN�КN�h B�P:A�dA��CX�q ��&D
0ZՅ���z+�X!�0)8^R{��d��Y"�>´7��P9mʍ�@SW�X]>PTE�NZ�)e��|�z��R��D�j!�g��4��M驙k�~r���oR��b['^SC܄[��������֭?aWKGn��+a���Vʽ{�Aֻ�����X�l%���o��Vﴮ�w�s75��t��}���*�	�����AR7/�	���[�༻���M������������t}��_�<>�~is�=kS��K[�+/@ug��Ԩq쓔Ǿx������~���as    IDATa�Cq������[������/�߮Ĺ|����l~����,�冫7���O�A�����<�ɵ7��v���S�g��H:�vCg�X3��·C���H�V��+�SN�3���3��B@LY�I'��Z�?�O�:aB�O�y�������&0��&�L3}�:7�h9Kz�M�����)�FBĔij4e����M�IEh�0)�|RNx�b��.�MbQ�P{N��QE���vX.Ajp��,[��sL���[�p|>�t4S#�.�p���"=M8�b�&^�.d]X����&����ǅ�m>�%J�Ȋr -Щ����nl-�[o"8�0!�P0�!~#�p
a�1�uŷ����apE��d�d���l�S��w�谖�ٺ�]ˮ����O4�2H&+�	Hr��$�m�� _�_��|��z�z���a�R��R*��d�d0��w���?1s#�!j����7Ɯk�&�:{oY|���.�gE ��� Pt5������4�-�Ԅ28�GC旂R"�fX�C��	Z�5"X�i�S���m�i�뇂�a'��Ⱥ�꣓.?z�;�A2ST�fqm�����/ݿ�;��(�ɏϗb���N���*��Rp�,���Z��N��-�,�F�!���Q|-q��^EkN�[�>':߆bs�)J`�@�s�-�W��UL���cvl0)�%&Un>�4Y�D(�����Ӽ�bD��������_~���rl٫3������뛳ý����_|���.O}�����yۻ�8מ?��ў�Zz�������������D����ƶ���m�����~w����_������_��ӗ�6�i#�2���;W�Z��

�h��99��r�٪�Z�=��e���������h8*1�g��CY�;�j9m&'S�Z~N�+ѺЪA�it����Y� �H�q�9�j����O���MY�� �
AF�'�T�i[f���u��	�(X�i�B�+Q
D�|�7�!�p%R�2m������A0�g��{XJ��u��Me�f��**j���(�%�12�Q(N�,��B�n�,a:��ׅ�@�iS$�Q��N�� �9��2�����)Á���ҍB�TI���_����G�X-~�F$2&���8��U������e�P�����I1繧��h|)Yҽ֕\!����z��jOqr�ޤf���W�g'O�Ԁ����H����,#\�8���TSj^�9s�ZŬ�DK�.�2�0�����"+��o���_��g�}&��U+!ݭͿ���!���O����zEw�ӟ�\]�s㯁�{��pi�C�Ȼ����Я9kxs{�#���������t�)5/��̻̿���#�����S@�b9VͧID�eM����˷WԼW����r�"�3�	�i7�hF��N��E��GK����*&YMLc!���#���F�(�r�����4���ʯP4���p�9JA.�Q�0�p&.�,��D����c�����5[��1���CjB��e���`Yr��pX��ʁ�͚VN�D'���!�p��x�4m���_�X)~ &����n )�ZsS4��hiIQX�Ɛ�CBJ��
�hZ��2GH
��(@J,��^�p�UH��Z�KV�1�o��)���1�|�"+݆����1�'��S��#xf(1��
Q�����
I��rp -���+�]5�����M������FEKr�jI�7�	����a=��a�L�2�ҧ~%8L8�D�B
s9��)�r@�l�pY���qL�8��*���);s�׶K�>���|8���WȔcZt-���6j���989��%�NkIaU�fD����M!5^a&��<�������-U��q�:F|�4YK#S�Z�Cd!'U��19�R6�b4E`|��L�I���V� ��8�J�y ���|�L��-��"`�Z�k����j%U��%�UK��|#F�?eq����i6�M��M��Rvn���:A�d1L8�3�-��Vj8t�j�Z��|��A`��Ȕ���qX�.ˈ����"��R��_�s-�L�AnZ�*%��Ҭ�JT'A�t��D�U�G}�eI��!� ��1��q�"�1�k�r!�pZ�h"�?��K�ג\�Q��>��(���c)FVQY�u[�Ԩ�D�kr*�J�Ĭ�S���Zm��;��ۢt«8C�lvhZg�wn�J� ~���$�4}~
r��2��G˟m�NB~j �t:�&�)$������2��W�,�*"�U��S��~%�B@u{�e*:�L�7��@s�[�V�F]IA��v�N�Eeq��c��A�A���n'$A�|������!�ÔB�������S��k�~���8�������8���f�����3~�riI�Ӹ c�[��^�9�z�CՍ��-��"�ԍ�SlU�#�c�FY72����n܂]�l�=%�f�O�1�c�Wk�{n=��o�m����������Gߦ�ε�q�ԧZ�@�q'���-���qJ����Ŷ����F\��޸ǹ���X��������\^���M��6��<~��k����7`��|rtm�n���gߜm�^�'���+�I�}ҽM�}׬����Ͻ\?'�m��@�^���;_��f�{����Uۢ���v�*;pF�Mv>�DH���Q�Ꙗ�<.]HdZw����2'��Y�lT�iCY��uR�r�L�&3�Db��p�Ζ��R0'ؔ'>��\=���#Q�xN��8�4��0է��!¨�!�˪!����
=�9pײʅ�,���W`�����m}Q�#h���`W�rdj��h��8����Zg_E�����[��!����g�čU�Q�mI_���b��N!"Rʢ��8��#�#*��4��QP��+!>fN�cҬ�E��w6�-7��<�u�)A�I�O#_(d�V9���9�12E�o�iJ�)$���ԙ�N�����
i �ƶ�đe��f3��L��(Y�Ǝ�,S4�R}^�=�U��咵�.�^�����}M�(���h�RL���W#� ���e?�@�\�E�')=� �"QQ�J�	Y!��Td|��c�1�#p�F�,P�Z��駟���/�ܗ �g79���f�d�
X9���2!���b|�q�&R�Bm|;�f}嬇�c�/~0w6w�]̥�_����Ǘ��>��w����?|~��矾z������/�?��o^������΃����ݣ�c���ٳǟ>p�����{���7?�l�myq���:y��`��΁���k���ŋoo�<���ή��O}��]z�+	��5�̙i9o޼���t����f��a�����؆ X����5v�8���W���IA�O%�s4��8�F&>&Q%���kL�1��
u�[��T��:�����C3L�>�xG�8e�B�Y}�Xn�8F�3��h�h�� guN�T�,��B
�B��*�c� 'Zd>'>$���B��� �>��9��!��4���-��Ci�V���9F��Ҧ�D6K45�"�kT���(Û�,��j��D«kD�%k4e�+�J�Tň��Q�GDϒ�v5�td�:i
�$R��8Bp~�q24��թ�M��jc�4z� TŔSz}����D�8�,:%
ES�˪D\JǇP�xKt������ h��t���DfZ"���^�z&�|
�S J��كc+8��Ɨ�}3M�\"�w->U����(��Q"e�\}j@:���W��?|��uvq�o����5���nm��ȯ^�|����w��m�[��v{}p8����*7�/���𷱛�>77.�6���g.o�}������Α?��O����������ۻ;o_����F����řf����/^�:��[k����.1�p;(j����|O�vOH�U�!t8��;���4�r|��P����a�ӕ/��N����6�%N�mO�DV"U7��*�g�Oc��,�h4mPCc���tf�xK��e�؇RpDM�q�8Fd8CX�"
i��u�bY��6
��ƺ"����Qc�����E�%˅������9��S&�!3B;0J���-���p��+RB���>pj#|��^㨴X�P`5��������Z��LWKǬ�rt*Ad�G[m2}�,c�R�UxS�9����,%}�j�ӺD�E!jK�u��s�r�^�Fd��`̑2���	d�pBz��*����NV�r���N�M����p SSz�d�fo�J�s�S�)�B���+�T9Y��q2Q)�C�k�\�[]��}�����\V{�+���L1E3E�b��҉�XP�� <M��:,�8ZY��/ğ"�,��/���),d�W{��?�s��DL����7�)�RЀF8>�̢m���Y�W��Z�U��<vUD �%�n��*�	���x���t�x��8u�Ñb����j#0|�K��3���jTiQ ���S ��R&���@�:��8UǄ��!j��Bq��#��<��ĩ'�N��9�T�HĘ�B�F����VK�h�5�,-����V��\'�K?�����)�g
�BH�hj4e��n�Al��ϩz=E�[�:q�g�NHo)��=dR�d�ڑK�U�4B�Z�@��X��3�2�$��Oc-��8� �A��B�Ͻt'���L�L����p ���%ݞ��RDgҮʥ ��UD��By�խ�P4S�x:�$�����xĵR�Bq���ڃ�V�D�8�U�HO0��E0�gS$)�L_=�ZrZgd�6�J �����M��E�s}[N��@��'��Z�(&�6�˵�U7:�[�q����҆h����*���������ǿ���T{R<0�N��P�nsb��0{朝�q#�����`q�t|�*������q���νÛ��)��us��ݥ�,FtWs�IՃ�A9�|�5�4�����n6�����������H��=�%��.뭗<��m���^o��9>�2��#�{[�~�r|��ʯ\��m�޻7j���;�`���A�0��N�5�4���5�@�G07nw��۶~G��]j{��wϺAzuy���б鶲�pu��ś��s����m�㲿�^����9z�-B;��[_ܷ�����^�n[�ͭ��g�n6�����έ��;`.׺۪�~��K����3��&��[v۩봁�{�72��8��(/�N$Q�BNfg��i��nbru�N�_�����/]��F�+Z�����(�~��G�Ө�j�,��k�������~亭+=�&�Ïɑ�;��M]u�����tec޵�h~�>gv^�r�T�ےӖ����1�{h縲ԍS��PhǺ�/DS���i!������E&�V'�;L|��u��N�pM�@Y���@f	�j����%ۥ��ei]>�T�E��Y�|�`Z3��|E	����XW��%4��32�����_!�����4�FHS�@c$���P�?���a6O�,�6�U�M� ��Mm;�At��L!�3��OJ��ie�?�m�>�/�A�V��JU�T�M'������o]�� �sLW�d�Z�LW�;t���A�Z+���X���)�"��Qi���[2<����Q|�zƁ{pe��P����g3=�����=N��Q����aCѴE8��W�H��$��p��# �Hy���2��kh�xL{\;:�����	z��h�opm�������������������?���G���^��ws�+ѯ7w��v��.��7��k�{�'�_۔�������>:>�zw����_��ع_��˯��vO��t�΋֎�"��';���^�w�OR�[���h1�ёc�AS�;c�v��3��Z��y�:ul��mO]4Q4���v-g�8m��Lc&љJ�g��Ҥ*�8|geY�%�4P-)�k�I���ӡ�7��!�RVG�\�iUi��n��BvV,:�������T�3�k�8�0�h�����~��h��$�6���S*Q��������a��9�arY�Qz�|�D��r:�A k,4����c�J�~b����S��&�%R��!��A�G(�4��4��8ǉ�־q -s��������H�o��Y�i�H�qX�Q��c�N	�@�Lb%�pL�g���1�ҙ�Y"�Z��
QkhU1�t��;��h���Y-�FO�E�X�W�qf//-p��R����WK=c�K'��X ��I�1"Ku����ܫQ�t�RW��h�x)"��n=r�^/Պ �hD�vF.��ƌ�h��2K�]1����������s���������p~u��W��=��N�.n�o������������փ����y����s�/�=y�_��?����_}��W�>zr�{v�v.�<�Z��9}�p_�^���}���_������޾;���oZ�U�Rٿ����?�3���������VU�Y�b�l��й?��mC����6�\ۂ ��j:�D��(SS�
q4�8:Eeq���՞+d��U�\-��K,k:�DV�NҬh#�qSm 0H�����8�d'�� ���Kl,dT�>����gbmHd�Y�B�Vݔ�� U"�J��ᐦ���9F�!��KIYH������)-�J�����O���:�)�`VTz��5��@�_�������c�TS>Zr�zh�K!�J�@c�	6�&J2e���?u�J��,���rJ��1�� _��l	�?T	��̝,
�
=sRUW'sp*A\�\S!�F`jE1B�)�(
�0᳦ш���[f-���+^z�5:=Є&S(k�tt�S��)K�L�2F�k*W!A#>GJ� p)�8�dE
��|ʕ�h/5%����vd�b�N���T])�����v�S�!:��\n�0K���^銏����3Y3�t6�ۅ5huh*]H����3EL��iD3f��@c|H:��(�lL������O����i|
hU	���f��/D�a�J���3��-��XuS!�)���(�W�4��Mbx�D�W(��Lbʦ9r��6q�@s����֔IięSmx�i���*"�Ia�6��\LN������:	ՕP˩4��9B���4�8YY%�!�C[T���+%�T��'K��_����p���`�0���I�˅[�fجXu8�t!��T�BU1$f�j�����LKMʬ%���1����4ʊ)K�)$ߔ������'&_h)��i���3B�Bkb�m��.TB�|��[�
����H�ƢtL�MkfV�Щ����/*�B�&(TV8�uqL�Dd��w�t ��CQ�SWD������h�єũ[
Lo�˙�.Dކ��mQ|Y4g�m��g2�U�<��ұ���փ�*5i�W:2�����
o=2zPi�V%2%K�&��,��u	A���P?m��;[��;pk����Gw��\_{������4�/�-� 7.����8���G'� 6�?�(�N�o-r�.��]�w^�*��x��e��Ψo���Nƽ|ߊ�k���|�/��?p	��\��;{w����!0!�vBߺc��3��vm����?�]v�}F����ڭM_��Õ�ne.��g!)&�
�5>���*�ܽ˃�w�'~<��o]�	��=�N�]�oo\]l���mo���ޜ^�lXέ������C�.L���u�ngo�ܝY�{��-7\ǆ�Ɏ5�������-�# C:���R:� ���0�e9m����T�I��rƝ��ϟK���2�名�����Gc���e��h�4�EM��?I��)[tҤ�B�HAJ�=.ZW�M�(��ב<��B������!jj8r]��˱���6M�?��\\��e�����c
G�Zq��B�����˪V��*Y
�8�Q6%��*�Yt.D�K4�&1-K����t�L'�n�$�S�`��N����<�9�X �tV�9��v�oI�0��Ln;�n��>��]�#���K�М�pj��%�����Mpu��ՌPY ȇpp�L��e�8�E]�k,j���_~�%B�)�m�!����B�|d&W��R^�M�Xc	�I��    IDAT���~��7N:�W�%v����9�.Br\=VT42>���p`�z�kUu|;༥#�~B(�D��t瘍2��D��K�$�������d7S-d��Z	�-pq{���5J���j�q ��S���"�g4���������W��WM;�Һ��Y^%�7\���2��a���󸺻�����O�ѯ=��<���ޣۍ�ۻ����{��k�Wۻk�;wW�o~�����'�}x�}��������W�_��{y:�&h}����7oO��W��z�vc���|��Q�|���E��i4�<�!N[Ԏ���-�Y���c&�
�0��ц0LS:B�B|�p�*�9�e�釉jO!~G��Nz��zN�m rR|j
�v����<P��oUȔZ�\>�L����S����cD6�[>�,̢@N�����0�t"M�@f
�)���R6b6�9B���,�F�Y�A*�S��;X�B**'*K.�*�I J4fpVL�lÔ�B���/��#�t`~:S�/ZJӹ�s:+&���	��4M���锝Q���'�~�O&���%�&<�&�r:��YnL>�/bC�T��m=�91</Wk�8�1)��J�3�MNU�+�	Q�	u.��3
,gQ�\Q)��R�Z!:�d%�@[*��%��j�#Q�|k(Yz)�ґѼ�x���HJ���	�"�Sf���l�E�{e���}Uz����$eN&��s����K=�5��%"�W��Ë�������ǯ�����'�����fw���w��kw���'W[�;�;۷�k�7{�O�~��O�|����������;/a��?~��xkϿp�6�8�E5�w��z�����޿<��+�~��bu�mw4��_��_���_�v�U���<
�l��ļ�j�6=	�[QO�R�Ԝ����1�"���4�F%dq�{Y!� A��	>}֭͛mđht�i
1H���ϔ�����R�>�^�Gv�)�0� pF�ZB%L3�j"g��'������t\E�ZMΊp�)5&w�j��i�̤D��d�r�|S% �d� �࢕2-ā$�YbR��䋚FéPM��!>S���g-N]���y����ު!|dc�pX�I�^��2���G悔X�5�a%qL��:%�� ���]I��UR��p(�� "j���(��B�(d�ZQ��4�R�&���)��<돏�p g�ā��D~x���)��i��15-q�,���2�����v� �� �u�F�B�f�j�6�he��8B��)#��@Jȴ��
>�f�g�g(��B̓�(� F�DZ��\Q��P��D	&���h���I������8+ʊ�8�NHS�%�~���@�
A���:�A��I(�h���\Jʢ^e� �x��r�5-�\Q#��&�2�@)�$�<��%4�9r[E����Z~|�PUf�pZK$�hZ-!G�)?}ӑ�,*�`]E�� ���8u�i��G��]�8�T���f#9�� (=Eʚ4Q4Ӭ����E5��>�\K�%�qZ�t�)0������15�G_-!3�rU�'"�} �D$"�9�C1��	��w�8�
�\��`�ĈO$��B�i��l�~dNjh8=l��YԒB�T_zU8B�V�h�Z� 7+
G��! +'+)���XV]YsDIY�V���E��'x��D#��hBj�әP@�~���r᭴P:S����e�����#@0+�� 8�F�Vg�)�Y-A�Rꡊ|�i#+���!2;�g�Á��-Tu~S��1ej�0�^�s�L�2��D.��E��O����%f�0�*Z����(�~�l�����J����I���/��a�0��H�� D	Ksܧ|��.�/4� @�14��y�ޓh�y0>�辠[�̧�}�ͰO�nRjg�����WO+>o���X�mx�&:j����/H�����"�n}dQ���X�ޥ���S�k^�F��*�^��n�����~is�now��u��L����6_v��s���8��;݅�+�t�a�ɴ�H�'/�ާ��Zgר��n-�ӟ@[:� ����և,7w7��������+��~v~}~��w<���[CW�ǥ�s��}������-������_,�_��[sǇU�n{��Հ�m�9cϗ��%sJA��ơy����i�9c��;o�DrRB˃�GQ)=~M}�d�uki��΢��!��LG���G`!�L$xNc{2��Qb�aE&^�O9�r��ٻ[�*�	�5%�A%'<)�I[D9뚆2	v&G9t��S#ճ)�����Ui�.�
�2ґ�*i�Αe]B]{q�b�ǡ�l�j���OMT�l����� P�� �)�eۜ�2En�@��ך�m#rњ�I��B9��%����b����L��JCh�&h
�1��P���J7��:�t4~��F�+�E���!є��,]-�%��z�G�i@`?I�_��7��t���X!�������B��V9�V��)&s�MM�ѱur�m1�o�S�5�%�� �넃OG�(MS]�ZT4��B�!F����)S;fdN4�\��-�uT�U=�������D<Z�Ǆ{��S@����Эu�8�Y��Z�o�k�^�L�C��<�]'�xc5^*=.�v����$��ߥ��u�{�����|����ϟ�����م/0���:����޿scs���/�=z��`o������f�<�\��y���lg�?v��G?8���o/^�\����>}u��챯����?W~z�k��\�[��[���5mZ��m���<��f�{Bq ���l�3�rP��>��9wl����ױ@�<�c���h��6J��!���QGG��4uh
�H�����2�ꁆKa5#*�\>�:�Цr!#�D�g����d-��q�W+����׏9~�|)�������{�rH1Q�~x�i�B��:jBVa�: �q �V�����!VL!4�MCLC�H���u�m�|���T-+f���q*=�8�g�?p�@Z���Ljx_ce{떦�ml�O?)~Sc!�6����C���t�s�tp<"hr<�k>�'���,5)p>0ߔSt����E{ֶ�r�B��sIrY����X�Ꝅ�,�)�@�����AuU��f��;�d�&�̔�	���W R3^h���`�N_E8ML-y2���Y]���8�bhD���u����������W��Y����ݝ����;6v������^n�\������������[7[O>�x���G����ݯ�������g��ٿ�����=�/O߼�zsz}��������?.�<;y�Ҿ_����=>9��`-�ӿ�����\]hjV�!�r�{,��+�L�G�`Y���(K���F��R��o��a�.E.��\�=�GO�u��L�ƒ�7�ڐEߘB���Th"�&RVBi�n7 �1M�� b�	�k�� ���'ĀƊV�I���f"�@P"�&
�C���t�sXR�y�S���:^h�C�P�E�/�>�u.K��l�ꦫd>�rJ�Ô� �8CX�`�3�wD|����0��rTl^.�i~��␕�x�ZE��?�La��S��%�9���Ac�M9�!�6⛖%aA��ɩ["l�rR�R�U�N�&����B�:�So@LSc�8�'��	$e9��D�Ù)�+�'���q�r9L	cc�D���v�BV�3\���B���^�zFR4���� Í�s�Yx�Le��Ea�K�a2��Yz��8���v�ZE)XEYp�>C�*�7N:���!����hr��bdE�s ��3`���3Ǳ0�Ug6�H�1��qRk]����|)�:�qǟg��ܤg-~�I �[#��M4} ����7`uM������4L�YB�~:�z��T��u�ý��+D��S��5���i�T��08!h��I���/k���Tq�I��ݮD#+a]qf��G��
�O���4�X�ٞ�#�bY!�V�cĔ���z���|#5Y�)�gR��7Vt*Sk"t��i6�a�Y�	�g)�g?N�x��
�Q+$?��������ܴޒ�7~Rґ��\���D'_���E3e���2.�QKԒ��0~�N���\�R�'��tJ�I��7�� Dr�e���B��)���ɇ�Un)� �A,j��Nk)]b��:GN�6E�2�1�"Cz�B0�ԉi�qX"�Me�45�>�b�m�����1S�`u��M�t�#��&75&X���8u�J$w�2��^TJ[Q�pd=�D���'U��4��H���$�&�Z�^o)��"SK�Ojz��T��%�\g5~K�)�Sz�|�Q�m�l��&%W��_�ڲ�M���W}��B��僗�'.�q���Ùw��m.}2�$=F�g_�����%}���q�ssm��>�D�\�s���ҹo�}����m����m�Њl�~�_!;�q�Wڮy���G��ݮ����Ź���xZÿr����d�3~2T17OGz�Q����V����pl��}�q�4�n>2��еM��ݯZ?��:��{wrs���H�k5�~�s�G:Ǖp_���}q鎥�����M��i����.?�ϧn�"iz�Qeu�Qg�؜�cFz�����pᶺ-����q2̱���w�� Kdp�I�����(Ec����y��
Ն(X	|Q ��X��e9���/g���1*�U K_b)�89d�����OJԦ���Ç�5�������*���C��y=D����|Q����Y.��Q]S�E��R��6��\m@�h������VR��gQ�P�R6&����u�V���m�6��*�Ig�����֥U=hR���t�=;���Z���5CО���G�.ARS-Ȑqt8V�:�[V��_�PE�u�a@6�����Ԍ�!����-���&?���E��1-��懔��Ig�H�q�d4H��6��Y�I�Yj�ҷi��S�TLR�4;�B�ˏ>\ᢟh-Q�fn�Q��rF�!��F^	�*ֳ���喭�����g3z���r{FP��ʃ��a��t B�Ś�=�6�|��5U�{�1v⺊MT&Ĳ��ZJ�c|`�9��d�Z
�T���"��x9a6�%�Z�
A�z�ip��ێ����v��`����������ߜ?�{h�.N6����nno������GO�={��y����y�Yϻ��ׯo|����������/_�������.�7��|�郍������J�%{9�� �����n:���l���@�,�>i�:�l�|ƴ�٭��ϱu�76'�u������v@F3��ƾ-���e�����9�ĩ�*�L	`�
=Kj��g��ԃi)*R0M��	G#�Z�ɪ1%��#Á4��"
4ҁpX:�L�͇T.�؞L�B���R��gS�H�2j[J4�B�@D
���N�5P��|4�\H&���z���)���9��~]��)ue��,Ω1	ҧ��;�)U�J��S���
v*��۶��G�{�	�U�dM�c�K�M��r�~�\8�����)ѻ>Z����r���)�Od�-S�Ǧ��΁��5#�oViȐ�i� r�u��B�#"�%N�B�9���dc^E�CT�OF=sD����d�_	�=%�"�ͼ�(͗��L�HT�/K�p�8�TZ-O>@���"�l���֮z-t�2�Ã��G|������x�mm���a�r�_�=��_}��Ϗ��×��`^�_�z��?~�����?��}p�ɳ�G�k�����o~:}��_�������g�/��O�����9��ӛý���7�6�x諗O�}����7_}7���+Xdu����W_}e�{z�X�U3;c��m�7�[�-j�@k�LV;�.A:ж�l�i��]Tۈ�,Ŗb��w�c���R5#�[K��&�h�29�!+E�j�
�����7�2	qʪmN�p�o�H�(��D��W.:Z6B0[HR��sQ��p��D�B|L>GEQ�(��h=��rX��8s��4#p�$�(���19�1�������Ψ)I$A�����jK|�h)���,�qV�JGpފ�Hk)%)�(>+�i#Ο�&9<�MUD�CN��9�p�{J��Q3�&���K����R��UtnZ��Y.dvȯd��R�#G9E�,
)�=���~4�L�V�Y�q:���=����n끲��]l��!��-��q�s���6�hL}���	\��%��BjpE|�Q9#!}~��eiF�f�p�2M�	�^p��Xn��rE�&��#Ԟ�q,�ϙ%��s�3�qV��N>�)+1&5�Q�|��!ued���PW�%��:��e��4u,�r(�ȏ�cԃP��qʂ�^NY�b* L}���(�з�����A��C��
2�+AQ��1���<}!����FULk�����#k�L��ޖ"��8�d�!�hJy�MV4SQR�Y��q8�RK�	���C�tuCLg]NK��ʖ(To)�v8"W4�H�[H�W�N�6"�-B"�v^��1���Y��������:R��H͈YE�5E�#��1!S�GA�,I�ؘ�N���*�_VOV3��xjь�4'�H2	*
� �h�LLx��
d�X�9r��6����(!�������x\3c��(���Ym���@>��@�I�NUd!K��1��SJ�d#Wz�GhD�q�eAڜg'�Y�#˘SW��2�\�d�TT�� %����O�k�7���[�hvuV7�4]��ߠ��BmK�.���k����jUTnk�gMkR{F�F��M�.��>SH��{3�B+Bhu9�����*��Z�_�3���}�d��yS��~��[����s�r�R�K�>�9B����� ��c��9}�����s-Ets�ngs�������>�owe��Zt�:�MP߿炇.�9�w7}����5�|���כw�~C�������������__��w,��o��L�⼰��ʸ�8�6���]���8=ݵ�A��Kмy��=������.��n���y��[���/ߜ�n^�m]�h�ͺ/�;��沎���wQIn�ϫ.?f�@��Sѫ���2>��l�ؚ�F/���ߦ=��v���΁h��2'��ީe�t��c���ހ��X��,���=�ZQ>.?g�($Tq��h/��V��-V�D��S���U?��A��U�6��Y�tU�_n��x\����mJ�E�؇����D8�GK���(
�xoU'H�a4��[OSp�A�#KD{�h��D���h��O �� q k�|H�6t�jAb��\����]IS�����A�dSK�QV�r9��)t"8m�k\��L�H��>'�V��w��<yBA��8�B�qtщi����9h�����q���DR�D�VE'�Js0���@joUD���R����S!jq���
]�"�ˊ�0!0S��.�1#+�1�9��>;X�?���K%2�8Q��)�Y���b���jr�y��d8�۟��;�;i�h�O\|���|����#����A� ��=d��L����W�)��*��b=k;��d[�Sƹ�
�2�F!���Ho�Ԟ4��X�]����������+���.Rl��˻�qxܜt6�k���+���`a�����n���#�ؼ�a��oFo����O<z�|�f{ck�З>�t�ys��������_|y�����W�6.�9{u���7//�6��A������suy~�p����>K�5����kuF˷u��}iN˷d��� -О�L��u���l:]����dq�"Hʎ�v�>�&��N�*�#�*@~m��A4SVK|L|��x�QN�t��.I�:��Ħ�O�O��2���b@%mfU���e��9B6P	!d!���-�p���%S��t:�ҧ0�v�A*�Z�����^�)+2[MQ��a��9��V�1e����P��Y4AL`%�gωLK�C�?9��VEg!�Mq~#|Ґ��V�_�E�BSM�ԯ�q��W"�D�{R�u>�eaN\�?��@`�K������F�֪)�!�+ǩ�@>�
	�b],#�S�Q!|'v�q��</�F��J"�W�Ӿ�(��R��    IDAT��K���A�/�`
h�F<!�P҃�co.��tK?�t�5�2�FdL�t����e~A����N!�\�[�^�m�m�n�_���n�<<|�������?�������������������gO?�?��ݯ�|uq���?;�胫��ݽ�Ͻ|�쓏����b�y���w�w�g[�7�������8<��5��'�ׅ�Op�{�w<����V}���܋�
/�F��9�΢,�­�'v!{����|�Τ ���B�PX�bl ��i��FD�Շ�*B�_��"+����5����U�sj���(TuQ6����_(fc��8���HL������m�H��~8��P�T45>����^�Q��,�fʓcW�cF��).Y�N��4�EE�A&<3�=��T:�#��j�<��3=#K�iZB
�_��!p q����CR�ȉ �eB���mӪ�ҩ��m�3�Mg	�r��,g��ә�q�
�]�IA�aM���@cG�L��1C�8Q�bq�B�S0;әBY�B��:�
�2��T)*�&7�`�p�E)3��m�\Q���� |��Pmg��D
��Sb;�oCB*��R�HJ�-E� )��[{M!��ьtZ�$��Ő����{�@�Y�l�+�̵�Qmh�ᘝ�)�䰪��',�~V�gQ4�9�ʔ���bÁ�A�3Sc��Ul-��c�Bh��h� ��}!���৉�55�N�P)I%�X�rK���L�C�����3!�F>������O�'���
�5@����d���NG�r���#XQ>}#�,c��3�T���s���I�,��6T���,Z3�3%~c �QP+>��k)"�A��Z��j4kf�Hnlu|�����Y�@(w�8�ω��Qz`~��3rqN��YW����,��E��T*�`�ɕ�|�����O�줬�2Vخ��W^-�NT�6A�5�42:��r�ԛQ2��s�!�jh�8��S�a
�A��Y��3Q
&��Mj�5-Zb%ڊ�!��X,�H
�>f�B�b�Ҍ���4)p��Q.�X֬�6�C�V���z�av�Lm�)�2F��Or���51�ϟ�Y�F��2�,�^K�v�TNg�Ka�ƺ2^���MK�x匌r
���9@��Y6`@L�5�2��>�� D�"_:P�^t�3V4�Z훐=�m!���7��|CE��ru�i��o��񵨊����ξ�o�2�ǹg
 ��tU�W�]t̙1��+i�gQ�����9�к�7>v9��g�����n��<Kcy���i	?ω��ܸ[���#�~ӻ_|tu髙��'HO.n..��}�ޝ��us��[߽g�n���2����㣑�v��H��ޞ�`����W���u��"�hf{yn[����qU_H+��'}]�O��>�nm�[��l߭�m��>��'0>����;��W�׮W{��o~}\�w�����|j�ʽT��a��������|�jG�2:�f'��w�($Bg��.���"MEI�%*�PF	~o�5�	���HH����;��t��íTb:�D4`�� #d| ���A�@S��+��1N#�ej�*��I�0��hGb� ��G� �Su���_�a8��^!�;��ŪeJ�=*]��D@f�1 �(����X���Z��e1�M%���F#�\�ji�tNY
��ꭢ�ެEEQ���Q�J�T��|`���Թ�lY�8m�������h8L:}��i>�Y�8��Q4_�1�#�l�_|���D�?I����(����3��b�ӟ#gZ����p�J�)���'��cB�4�^JGk�R�1!|)"h��y�T#���c:��,�,V{��!w�y�k�j���^�܄�qg�X�-nu��̴�
A%4@��U픖k՘�KDS1k��B|��Bh�pYV��i;���SL�>��3��ꫯ�}M�3}0=A䣦�|�(i�`l���r#����";R<��r��v������rz{!6�N�m��'9��{.w"�X�W]��+_v������wW'�;kO�]]޽}��M��<����Ç�E�<}��ɿ��?��s�y�����������������hwn���w?�/?;���O�=����O�{q;_�rrhٽ��.��k����2e�eK��BY���4���� H�;o��Egp�;T�8L�s�t��&�Iw
:~�Y �W.�/dt�T�(pк��	K-x�B؁Ԫi"5�2#S65�Us��L�Ң���,ScG
�?��h�v'�(�ڶQՊ��Vsp��(�tb�3�oL'DW�JP�P��9�@�j���p�r���)Y�Z�)NƗ���-�5Y�t|L�
_�3��$�:rN:%�Y�@J	�b�F���[2��,�fY���� �8�H	M)�zC�)�1Z���q*����q�M!�Q%�F`N�	�5�|h��$�q�L���h���Rꍣa^bZ�|�G�֕f���dZ�h�h�`��C3_��y"R�S�~<G1�g�z�5P-Uzh�H��eҋe����|�2�5#����r�q�`TbĄ�!**���%�ZU�k'���~������%��~����h�{u�e��GO��?=>����������7�Tu�j�p�����������{;O>�|w�~����������?}p|x����9�x�{���ݏ?���`�7��l\�m����P?����E�\��z�u������}���$����믿��v��4o!��Z���=�"S���֡,��h��,5������}[��_m$�P�����}���#3Sׁf�O��KD�cQ�S->'��5FF �����YU�!��;�@#�z+4ӏ�f��D3�n��gl��,��%�c�Of99����c|��9h�Ԅ��ƙQ80�5�**H���g	xʥ���,儌�,�D�D�!�ɩOS8C �q�8j�*eNK��tL�����E��ᬢ���E��B����*Wt6�Ё��2�˚
Y
���-�H�V�%6
�)ku���f�V�V�L'?54��6��S$P�Ʀh4e��7�	6�SP�89Bɚ��fJ��!�M3�����m`��a--I����M'�#R�M�ԇSo88��8)��,��c6�-�JaM���0Q��T2��;=8!�qѾ?.�!B
'M�*�Ӹhju���BJo�B���N�Y
B�Wu�8�(f��*"�Nl9|)BM9)�r�tȶRQ��Q�S�D����M��4�d"�h���G��);�V��>eA��
��o���YQ�Z|"aMeQ��hf"�'1��O����j��Z�����(�Կ��s�!����1eLN��i�)j��p4#K3M�F&7B����2�,M�!�����
I4m]S�I2e�Ƨ��ac)3J��)�U���J�!R(��1B�&�PԔ	e�φ�rb�"�ȇTE�I�����$�a���t�2U40i�����1��PkJ$���C�K���|�$��ƑbTq��5VȔ�1�I�c'�T85�3�հt����L�hZ?FVŖ��L�)e2���R��@��Q���	�U�Bq�8Y�_gF��U!�B��s�� �n��~I�	>DJ4k�����(����?�2�M�)^J=�M��r����w�"t���)�O�nJ���)Ͱ� ��Z�2��B#|N�҆�ր*D�7j�����]X������w �d���ߦ�{�z��$̝�ѳ��_֫��y�(��t'����|F�U0���ť�����g��������wuw��s��bTa��M�5|�3��9ʻ��M��s��K�r������nl���]����y~��r����rZ��}��V��%�5�?�9>Zꎨ��I��������J˟b���[~�fk���D7�U�^<����gv�����f�Oo^�����-\ߠl1W:[w+v��59�/�.�6��u�ƽ��c��Utή�m)Y��c-4�>;�L��Pr�=�f����:��`:��;�].���Bc�(����:1��%Yc�)t2P-QR�9�"�P�&���I?_n�M�j�Lh��4�I���(ך(3!��kG��.7�M�#%��sVOA����zi�FG��׳f �@��t�P�s��[�9�JS��%"��%����+-|c�C)����V e]�CVT�(��Sn����J�ҕ�5�oj������[KU�qR�_E� #s�E�?#�׸0�Q�\�aԈG�CP�d9��B�,��od1g��1"��9�#��B����=�I	U8k�i��#my5���`Q�
1M�*	t�!;̺*7��p�C贖zH�J����g���SCc�9@
i	���:^��UDn	9��*��'E��D���1�*u�1�RiY,��ly�g��L���h^�F�Ɵ*(@�P�:r�U��G���A[
�]p2A8J��XO�
|fM�Ɨ�߹9~PӍD�Hk������x�X��/0��Iz7��2��p�z}w��'>��B��;=9zz䣞��������������w�;�۾��Ϟ�퍛����_�>����ѻ���k�~@��'y���;$w
w��O}Q��Dj�]��~ñiW���u�Fkgv�f����� �l����I����_W�Ϟ���>��^��G�Pb9�<�tT׆���45<N�3;�������>�ON��`%�l!�q@ *�B� L��t!�B����8�f��8�&�f"�����t�%�vI�jU:)!=�mQ���)�Sυ�M���u;{��B89��%r�-!� ���NR�6"C8��L����/+����ʁ;g���e�F�F
f{@��f9a&3��#�&H����S�U5��4�/+�dN)F�F�&1Egc:8B��TYM��α��oD+K"'��w�w<�`*�q��s��HXB�Z��{���D���V�[fi^�<k�v;F�Tԓ g������N 8��1���,�?|�X���E�Fͳ�rJ0"=��9��T֋���ЉCA�n���� GQ7���'RR
駖�3Q�ӓ���,
�@������I�����;�u,��<�w��=B1h�V
��������(��V���I1����;�����D���a�m���fvxx�C�������˿���q����?_��]l�m�(}�䛯...��o?>�{��A�3������럿���_|���������՗�����������3���������+�O?�ܽ{ru�ӻ[�>}�U1A�~<D�
���͚���z`O�m��je��=Y^)����Z"^F�(�	i���(V� #��C:���ڠJj�H1���>�
Ї̞�&Dc T-���p��"ySNd�l�Zj\��HdfT�\͑�l�������R�IMy&!˕&>�>r`}3�5��ŠP��N���_R��fR��zL!��	o%�%���lH�A�.W�!��D��
�Gi��.�(L:�R�A��<���"�M�2�\B���+��٭d��jy�\�I��pA���D���5DK�!�،��A|����\Ԕ�Y�8~�Yj�7r�z�R�+��2�r�%���hޔ;~���1�8M�P5�)�yr�k�J"���k�.�ئ ���~�crM��h%-c�8����N2�C2�Ȟ�Z1`F�������\lH:�4dw��q�?h}��2��U��,�D8�j@��	V@�|��*���iw��h���5�!�<�(L<r���
�!s	��}đ���}�����B�,K�HA.䊔�͘ C�\���Y\ YL���6��\ՀI��Ŗ�PxH��Y��Id?E6�EH�R���c��R#�5 )M�j��X=�p�\Cv�ȕnȕ��ι;��`j�È �� �
��2��%�� �� c o�@}e �̼�@��J�E���cB�p�����|g�Y��&
�!����V)�A�\M��� K�*j-��gЇk�c�{�G�w2��)�[�M'0�h��N��RC����,C+�ެqJ7���pG ��c�����*C`��XI�!)a��Q��`�14j�@�!�e/2c/�T�@R���f^��)=M�D�Z���������5d̞[ϕw� ��.0&�1�U��K#(J,;�(��������=���/BӉ&�Q
8���Q��1��8��������KQ�����EU!>��ܩIV��p�*o��q�"�`��A4F�&�v_Il�@v���r��[��䑻
y���C����A���s��a�܇�KG�7��]���#]f<p��㔏^d������k��㶶~�����`�ù�˓��ə�.��B�SŦ��.WU��)�6N�.j.2�6�ctku]'<��&����ٸ���({<SҲ��c��R;^�z��Y6��<��a���Z�f%��qK���ַ0ww[_�t�h��Z������+s}2�-�?����ǃ�%�5����p3w�u����ܗH�5|�j�Ou�Ö��n5.��9۔��6��b������p�m�me��mbݶ��g��iN�5�.�1RC�'��e�aD���p=L��4gTC�TL����̅�W-;���6WQȳ 6��gkB}���˂���Z�e����ǲb4�+@|C����	��]#B�K
���ِ-����Y�IG��^��>ڮN"�py�jN�E���`O�����\l�/;�>BU)�@=��&\%bc"�PF����1
gP�c&%��C4� &Lv/r��Ŗ���V
�t
.��!\@|�Ȗ�ls,P
L�Y-;5�Yd�B`��80\T $Y�����U�bF���@C@C��CxS3�2�2�Bo'�'D�}�t��]�'G�pC�(hY�����@��ԄhB0-rg�b�,v�bV'�P?R\���b �V�]���\p�4s��Pc$�.�E�PM��2�W�^����8� ��2���&q9�x;��a�3�rIl� �Eh�����8OBJ��.g�gǳ����õ��=��~��~}��Ci�����������/?{�۹1��o^|����������޼>9ܞ�z�O�{������7_��0���}\��N���{��-��ۺ��x�ޜ~��k�8[�w�KǏ�`er��9@��g�����lL�v����r�7��V�є-�ri�1��a�<7�p�L�B9��(���v�!��mU�M�Ʊ�Bz �U�ŧO���ڵ@�@���׌iȘB�.�*��b�����Yvyy3�����K1ή���dc2 z�M��� ��Dƥ�h�1�B��/ġ#P��L~^=��A��%b�pf��
Ψ��a�-���\����OD�����^C�9����rM�������*#C����a�|�U���R��NJ_�@mFsM�4���j��	����+ƅS%8��Ȏ�02Y�fͤ��D��Ԁ^9M/Z`�V�"�:�SK�@Q�H�٩��h�2fU!�N��j&p�z*@Y��.mR�e!��2&�3I^RR8AQn�z'-5!NVI��� �[�`h^p�:ו�T�¤<��h#�v+��
�/?r�o������idws鵓K����������ę���ݍ{�����SSq��h�}{�ө?�ᣧ���f�a��~�������������?J�x�z���_�������_}�_���ݛ_ܺ�{������~:���w�>jq֟~���ݷo���tzt�{��$
�cϏ��>,:>e{0~��4���X��=j�L�R�r��h�HY�6��9�q�!Ñt�sS�U��5�
������8-@�j�k��`�4��&4����ԄK�_T=d&eD�)0���
���5DKG�9�}<M�!�f]OXyD���2��e8�ԐK¦��gCJ!�E����g��(�f�1#�ۑd��eD`4���<c[^�X���Ӕ�Ø46B�� ��P�8VI"e�ES�� j�4!bC�MJ�&VFy�v�t��)�#;<qB#I)�["`j��3ऴ*a��+�H)�(FS�&�&
A���y���h���dy����Q�r1��	��)�+g    IDATG̲���'�-�YWF.��S1zv)�f�O�8�aY��I��ǩ�V��L9��,�������S�,*�eӌ#\lv���08�C�k��T�'���f����\E�z�*oK��ǜ�q�Ţiz5L�^T�����3��1٭��!�E��̮��*I$o�"h�ȩ�h@��a���ǉ�fh�H����S@��;f�e^�4eC4H}:s� y�I���!oe��X.`��,]�qB�,~�̅ւ��)$o�@M��,��+�=�O�2��gj^���35ܰ@��*���&�2搑�T���0�Cf��^�X�>,�� S����l
���bѨ��7!\�=�J��1S�шG�7�ҕ���P:`4C4M�];2&C_m��΍�_�Y��Z�Z`�+oǞDd�՗7}L�X��B"T9{�.��n���B��V�Lx��W "�"�`� P�\�##$��4���	z&�:�r�5�R�;��Ŗt"gy\�d�Z��d˩�i�>iiB�Q}��~U�U[�d"$��xH�EH�����-
�T:V�� ڻl��-''��u�HM,���D�
a�9w9P�\yhI1�C�A
�������� �5����,{l(�R�~�!&A骤���6��ވ���/�� �����è����4�k1dͰ�RhBhVy%�C�@n"!��7�;�|�Ы4oa�{�����/�ج�ޣ�G�n�ȸ��J>8�MJ�&���7�}�;�������X9�����?�\̣�g7].�ި���E���'G��~+W �mvG����o�ܻ�q�V?�i/�����G_��t�`'I������v�:���p����VGk�IV�r1r�����`�]o_�U��歟������c}ws�1�wVww'��@����>�,��������d}y�}z�:>9;X���S����w�����k���u�/���;/�-���ՃK����w��s��Լ�j/�T�;�����-��	l��ӎ}G�-�� ;��v�;�����*�h�����=^�-�xgx� �*��Q^�a"c�&|"�
F`hpC�R�iX_me��j��=F��%� �a`vCHRn��zpd��4d��Z-ܲ�v��nX:j&�<
��̷��D�jL��/�K�e�l�%�e�)�B�RŲ��x�\l`x�Q"��4�TE֛i@L��)�bL�&�p�벜��d�p�8ER�
))/A}k�)/�W^�h��-�D���H +�GF�]�!q���(�a�E��֤	�B�lF����?�U@���F�ԇ��n����%m-N�����G�k���J �'��&FK�R��}BؚDC��h#T���I
G���j��&H
����(FS��Y�?L�OAߦ;de��pl�=[F�@�Ȉ��M�XG�������k��$�����r[J�� u�\r 	i�K��W�ƈɠ��Y6c<���:���/B�og����|��C`�fK�K�kO,�����q��95����M<�"�\�����ݝ������������o��|~����|�z.NG㊦>@��N:��zܜx�9=xu~��ŋW_�|�ͻ�ݻ�����ݑ�
|�]��'��N�9���x2;}v:ni8�B@㖢�YUKd�2Z�V�ry�8fm���, ��hѸ:3����(x����h;��[J�N�RXy��E"͐ln��5���[
 �p;^@

�R`�(}�YR��0G�
h��k���[���h=\O���)�P���!��+iڌ��+�b�󲁕�H�S�] ������C&(�a���֬sj8p�b�T*&\,{�ť��:3�,*�5ąP��zvI�
�� ;@Ŀ���ɥ��Y�1�ZH���`}���Iř^C�v�].H�r��s1�"�;	��OVo�����!���r�v+�3��-�ı�@!�SF�(`��/��/��2�+@_���=^I5v�����D�k|�n��j��ς��s�1;dj�1%*�@��
Cg'���8o�;���A�A� 5�@C�dv/�:������*R ��tl�1[4j�+~NcեV�����h�w���x$=��Lw�9�rC
?�����xu|�2�g'g�S?�|su}u{����rƟk����}kӻ�㪤{ќ~����g�<����|{��������������������OO�^��|���������wW?_+�KCG�C�EY7+������W��5q�-�����y�5���ķ\z:\zd
��FMsz�;p^4�!��J��vA�I�W,���ήx�X��˨UB�!��"K�!/<{�ZQ)H��O����dT��<�M)8od={�%>�'�zsLV�����3Jͥ#3(@q���J�n���T���^�a^ò֦HsǤl��%�7���Z���,��*T	[�^���+�XLjz9o���C�q�pC����;nؼ�Jh^l!��1���V=�@���N�0BSӓ��O��k��� �2�)��t�8��>]�f4�\d DUև1�����!��h��y�>o
�\���]�jČ�U^^���/Z
���kj�Ҕ%W�@H��aH/k�L"�z��8@�f�-�i�gU��s�hR$�
�|C�a+�0J\2vކ��cI�Ѥf���țB��CĆ�E@�O�����ѐo��ڬ9)�|�	A(��RT�(8^l�=%E6BI��\^x)THM�l��±n�4H�h�� 5�r	o�P13�X�0B� #~�0�Wp�H*�*)�p o��S1!�R�b����+i�I��+0�@
�6\S�,�!��p��>�ʠ/��@���.DkfU�h��0S��%t�5IG��&�̀�a�!�)Qd�����Y"����8�+C��MK��~��CrMre�5-W=�Է�[H=��"�a���ɫ-�D:����r���Q�r"�����T�~+�L�a��z"r��w���)�5��|�AT+c�V��0�8�gH��c�URϋ_���ᱟ]ޔ�hp�&BA3��j� �M�4Գ30a�d�{M��o���:L�g�,��և����ҙ!U��y�&�h�U��j(�f�R�3�MO��m�פP[��\<��f���Fs�Y�ɇ�G��4�zu"��C0{h#����H9>��?j���MS��un����畢!o��,��J0��-Y��Sp��	�>���6���3�vur��V?ّ�K_w�W
���(�x�\:W�܋������3O| �ЏEښW�\e<�ۍ������i.WRp-�r�ٱ�f�:�ܮ�(�ճ������ݍb�{���z�.��5��룗��ǳ?v����|q�{'~,�گo��K���w���S~�l�埫����D��w���z/dq�G��x��u���<]��k����K��"X�������;�o.�N�'�Oi�]��m�x�n�\�7 ������c���޷�) �uO�Q�������}|���
+���W���|?~j������MZ�/��� �xۼ�#D6Ԥ��=�}��7�������O\:o�8�R�g���H�UF��G�pF��*�N)�z!pF�|  ËՋ�0�{C��Z��)�-$w=4��i�C�Y�,Ԏ�&����&�Oؖ���#Ք)$�I	^ &���4B���5��^˞�W�,D4HKD�]�aKQ�|{/��#�\�_.50 �+ ACYJ$��H@�e@�T�(æ�N��Jī/;)!�����#0(�$ZӤ	���.�9�2
G�3�hE%>�%�q�0'Gx.��*/j�[Bp��!�G^�ae0Cf@v�b�H�z�$V�X50�B[�V	�Yg��Ch}�Ii��*�sMX"���">$Y}�\l�!#��H��V2�J�K*�7:֡��`hǽ��)��a��������eN�"�u��M�<`\9s��"��tD�
Qr�"��7yCMYzj���Z���C�g����ۓ#���F`�ow2����v{����.."l�K������ ?������ʇb�\����������z<��7/^��O7�;��@��x�4�i���r�x�Y#Oև�����[�z&~�ŗ/O�����������#CB}5���3�Sۻݨhu���;?�����UM�큷g�؂�mkYp�����`Za��v:vʳ��I�Y��B )Kw����()�ڨp�˘��X"�R�\d��Z���R���{����4� 5�l��2�LA�148o��z:z��8�\��p.H60f�@�aR�Q7敝WT!���q4:\�nXIM�\ȆS���?��0�u¥� ��x�V�Z���Ը���4F��Z.i?�zb���#O�j�u�BJQ.éoٹ�hz��p`R���,D�l��X���(���	7Y ��K�װ���i�?��Ґ5d`!sM�5WCyۣ�8�!Sa�<�TC��� 8z6\Od"�)8{�=l=B��]j�p|}���"n[m��%�-):�.ʉ�sGϬG��U32��֪Y����.g|Q8\
��|1U�L!P=���]U��m���x?��g�??;]y:sw�Ϟ?{z��\���\��镏������������O��׻��oV��}��~��/�>=;?M�����'��qvz���_����]<�aǓ�O^�x��'O��go�/�~|��|��7���������oO�����o~wy��K>����Ŏ�c!�%�y�Vl�0}'d��Κ���h}�U��L��bS`��.ͳ<>e���٪��dTO%aVϲ�㡍3i�k��hz�%�Y�*i8�R(�2�a�sU�$�ЈL#Z��F
!��>�ÆB���!��Q|��1	�⑉T�,������La�N
X`�D���D��I-�F�}���\*� t�Sg�x���4~R���L��8��)�5uNqC�*gdW[..��4*{δ	���wx0�1��'��͚#G��f���s��2��0�ƾ8��>#�^���!A�\��k�Z�hS��aX��(Wm+�eX&<��8�
�t2[���%+�Ӱ5D�P��QS�
�G��h45d4W��h����0��
�:Ȧɕ`Rb˅Y�aLoM�V�hr���ǿ�r>���BYF�B��ݬ��@��d�jj@��k�$�N��4[��@���4��hrD�rAh�`Ȧ��q��+�0M|ubN}��:��%EY�Bg"6�(.�!��N��S�k*WI�P q��"�m�J��X���1,2�����v�e�)����q��!�\�����a �5M�b!��K��UF���-�S���S-Z:b-r��T@��VRYH�Ѫ�-v��a�2dd�&!� Y�@#�`X����d_��3�*�>o3
�����r1*�`6<�4�-��!��eI�����/QH/�"L)����T�E%E�1���s���g[ʢjpF^�-D,p*'%�;��F�Lg�����\�Ef����a�2o��gv��iy+^Uq�eL�,����T$UlQz!b�)�eܯ��\8l"*#�^Ƽ\�p�ɲK���N<#�\�d�O��jB�*�ϋP���0�DNAo�RL>B-2<}"z5��Q��)�15!8�\zH��(�N���zxQB��p4
Cz���,�@�bټfgXv�l�K'��x�^C1�)�p`�Kα�d/�{7o˜���#~���������z9�\�sf�s��P�h�1I�s���/t�l���劣���q�Y���ˇ-���O��u����YZ���U�w��*9/��cx�e�g��S?��d�x����?���>z����é�i|��ƍm�o�ua����v��V��������͒�]�6�w�r�l}��O�r=��;~���WI�����c���c/��pw�>��'��?�3=?=��Ξ.0Y*��}�����z'��ֵXKjm�3&h�|9�=�C}�9�f����T�����~~8��6�Z�k��+�e�P���}
��6���Ey7 ���-\�=��V�����o g��[岼�m^���j4��5�j(D����x5�f��dK*�!�����2
i��'��3�>�Y�
5�i�I"��궴��H��l�Y4��$���\&�	T�@(\�7�z��v�K��!)Gl�yت��6���X!n�a%��P�&D/�x�sT��X��MP�m��q@.;HM��+J�2b�	d�r%�nq���e8�	�Z���)�7�ĉ��2ZL�&\kM��+@��.��\�(�D��H6&���K�-d�X�]3�N�8t�(�S^�C���\�	���$�πϤ.?[C|{*]˨4`F�aY�3D���i[(
�%.��*�T����f��Av�L��}$@Z�j�l@��
�,P7��fF=@�U�Ǉ'�/�2�,★Õ�)���AG��)��#�믿��_�ڗ�]ݔ��yV�s��t�T�� Q�r���5L�&YG._)��#~�{��y������;(gN�;z����f���]�ܞ}<	:��eo|���_��������t����Ó�Jm��������ݐ:]���qK�X�y2�]ix�^y"�A�������'�/?��ޮ/|������=�)��S���n7~���X�/�z���Z�K�&evQ�fm ��Z+۩�ӊ!�o%�����z��a�-);��eR�]��'+EG5� ���\6bY��u�N\H{�cH�"a�CY�t�1�b��hdR��k���W�T@(6/�!T�����
Z���P&��/)��]�e������Q0d�����֙���*{6�p}̡��$<��3J!)�(8'� �\yl�΀�d/�>LX��A3��ΪI�bk�.c#2�R��J� �M'Y=�h�e�j���d�	)��7B
̛ �@��K�CH�P��� a�=�_F�Pٌ
��&���PFC4�UU8&��@򪊷��`j�s��R`�V��t&�d�R���d� �2�K�E� |�'(�Oi��Y��sZ�J�Aơ	gwNP�9:�Y�t�����SWE�D��!n�zo���O�M�Y��حkΟl\q}z~�x|����}�]����E�Ob������=sv~P����3���G��6_|���3�j}�/�>������q㖇����˻�w�__<~�f�����������`������6��r����^��js���aw��諚>g��2ɓ�WI�����/z����¶���l)�\6�E��8Z�I�"/�ތ�n�m�ؔ	2�Q�rd.P=v��o7��҄�;4v�!bg��Cqi!�ؘl�ɦ������V�u�`��L��xKgj��\^��h�+�p&b7D����B�j"�!��J�r�� NB"����(5���u6,5N�8� _#�Y�B��൙���!�kQ�p�bs�P�!H݁W%���k&�G�7w�Y��R�ǲ��	�5�U2�Ją��B53 �(b�&PH�����Ѥp��Z"�cǙȦ�Gn�+�ԉ�e"!�U%;�P���@5TLC��<KR�8e�c"�E1�65�ɗ(o�ͫ��t����- ���(�AZZ��r���'MFH
͋lL��K�z*���qe�3�Nٰp�Fg�\!���!�2&3�����;��H���UvF�%^ޢJ��r�
�\:|�&�	�%sq�y��!P+5�����B�'G���>m8����y)�M`�^ßR��a�����f:�s5dI0���Y?az#��5�8f6��l�6�1�O`�J����6cU�3m�ƥ�N�8��r80���!"P��S���l�@}Q=�����'��><�a���5A=����s	��ID����0�{A�+DoX�@���.!).�I��2��Q6CX"H��
ġ��1��b��ؚ(X�!��B���&���n�1��~�
44�Yd"� ��!��K�n���n$�xf 䪗B��Jjh@��U�h������ᜩ�+�f4�@CSc"Tɬ0�,�Zo�Ⓣ���KT.!��'��b���ό�q���&ˋS��]C`@"�1�TE�
�    IDAT$�ea��Kc  �S���U��0���zBĢ�T>'k̻�>0q*���c��O����w��L����.SS��h�R�B�����BY��zC�@���0������xK'ȫ���p�p�E�J=�rE��5^��@(֥�\���UAQv�K6���p��q%s�+��>U�z�ѕJW3]|�뎲G'�s���|��y�������78����\DT�tc�۝T�k�����]�\���g��O�^�z~w��S����<9���z��~�ۺ *����#�]}<X��;�;89��o�n�'�.m��J6�0�8�,�/�>z�o�yYo�]e��2�3��⊦_�;|rp�6���u�]WeO�VϞ�zC��q}�b|���`s|�k2ח7����Z���թ�.�ا-O��~4�<�e3��c��N��ꬍB��,�8fx;��MJ/
���#��^z�'*�ѣ��q������S�S�q��x.﮸�c�G�H�J@�ג��J�!�IQ%),�lS><)�58fQ������Z�lCM�b�&C�hSS��w<�)�5H��7�A�Fop��(.v���HYJ4��Y�=����"U�Z�C��ڂ�D�z��(L��R�ըYp!�D���\Z�h:�D�A�!؊�b��J���U�����W��֪RB��Z�����X5��3�
FӸ�hDl��+���E�5���Ov
1)�����b��~���5�UbX���Τ�~5�
�Q	CxbXyf�ꛯs�_or��3�N�c��s���'ȨH�B̆z���P�^C�Ya���� ۝�S��1��%o�ͽ���ƠbxI)	�r��V��@��܁��3�:�Ł�.�)��N��;þ�)�2z�m�cqV.�y�;j���E��VMU�ВIŕh�k��,.��5m����#�AG��5�3̎�1/;��3�����������xGzs��no�����O��?����O����oߜ]��>|��we|�b��0ZG�[�d�a�5�'<5?k���<��49jY������'�W��n\9��&_O\��Wn�>�ܯo=)��iOz��m�N���,��*[��������04.[a�]o��6�ݵt�V����u�<��)"l!�����QdOeDS@�*��)�"W�h|t �N����
Υ� q�e�`(AK�����10����-��\�38�@v!*���"<:j��R��-$edC�z�ꤹ_0Z�ٳ6`x�lQse������Ѱ(:�\�X=��
N�"��{�]��hs��D��8)4��qr)�D�Vys��P_��E!�edS��2����0t�ǩWF=sJ��9΂[�h�������7YZH���K'��>C �~�\�Dm� -�t�=$��r���#�TYr!��BD�gQa� P� ���jњ�sWO$�y�E��4mփ��I�)�&����x\�!�>�%�D�7�IT���	E_%�5O4��m!���ai��'��44'R�o^���ś?�yt��bwx����>�\�󻷾v隆�<���/./~��۟�/�؝m}��GYw�������?{v>��x��՛�O^�|>�3��W��1/~���_�����_�l�_~��_����n^��������cG�������O���^�xz�r���v�_�4q��Z����,&e鬆�[@�������\C�cxK�`˥����5��[@F�p�	Sc'�߯_%��[I�l`h!�d@0����6�i�0�؟��)�Q=�Q!�,/�H�]�4���1��@4H��x%��:oC�H��qE(�:r�Ґ�*�3?Fx�;�b5���0!p�4㷞5�g3�ڗ%2
Zdy�ȉfD�3)6C���/�g8o�x|=$B�s��d���GK9F���jB�v�5���24�4˃[�Qcp� ��!zHmN�5/A#�S�%�Ȯ�"^2N}C^ M���"T D�z`�8�N2��&�PO<|�y�[�%�8�
7d7(�-{H�p�Ł��\,e�䣵Y\�f�a���~R�:)�SR\��#JH���"\v���Nnz'F`�pe�K`+�ljRZQ�8��D�2Ը�H�a�ܹ�Du�b�M�J��F�H�%�C 5��b�3��:�Ky��g[C4y-�p�r�Y:�͝�[�T۟��d�.�ZR4gal8~��%W3JR8C����!�i*2>����cRXy�ɛ&p�̼��k3���b�5ޢ�h����&'Z�
CÁ��R���ŧ��3���q4�Q�ǒ�x�/C�aX,��lF��V<od"VX��E0��WRu��]/��f�Ob��e O[����X�>���Jm��5Km8�"jl
ڤX��U��3x!�ˎ��%Rߔ��Yc"�U��k��!Y �\K�c�T�`�R0,$��?�DGƘ��'h8��gț�(V�5ԫA�B`�n�6�\�f����৙=5���[%L���4��U���װ�30B�[[��TX�鳧H6�͎��@�9�8E�E��bj��r�ù��W<Y��1��Ȣ4HY�(��7����]���Xr�+c�����x�'��g ���s��^l���R��*x�l8��J�$�����6M��3D=8�fQ��ʂ\T	N��F`�z��Ad��1��nt�6}�r|��K�?�n�d\�t�����F�"�S�@�^��.���}G�n��n���M��A ^��>�����5ޑ�?�?�)����z�j���ڷ�v>�m�<����7b�3V�ރ�f������v��������D�.��+�+G˝�9[w�_Xa9f�R,�x�� {��/tZˍK����"���=7.�Һ?|�������5����Se=]�)�����nW����ћ��������wP���������n���}�3>�y{���oP[j��u����n��3[�kq�a;�↎��\@�\�rlx#%����:¹���HnX�l=)}ǌo�R@��(�D��.
^��Տ<ˋ�ϋ��������4����GH!e:ar�h��z� ��p�6�z���(�d��_�b��e�h2���6G!�d���j7��%�('3RN���J�BǪ���̧�&*2��l'4��zw�����i:�V�T�M�wx���5�ZFم(�A*�,i_Z��K�t��zrR��@�;�)���Z��]�O�P"gh.����#c
��]8� �B�nHj_���&�:����H:h@C��e������by�H�w0��V��)2(atX:��3���2�] A��L�Pٕ�����g���E�e���K��Ѧ �~�D�j��5�0'Y��-N^�: L���S��ty�EM�6�rQ�]����OBX���qͬ+���)Z�)%���+�WS�GP��=����;,��1�=-?9�+����S�k����>�7^�H�Y����js������k��7�&vO����Ż��f���~x}���Uܻ�����j�nn���?�����kw��������G��u��Ϋ�����'~S�uN���O>_�����~���G�gCwZ�%����x�����qKmw}�n	�gO�/�z�j����?���5�˲��bo;suX4�no|�i��B���[4[�b���c"���1X|���@Y|ِ"w��A��!�*�����r1�SAF3b4̦ �͐��� j���G��.�K�\	��,�D�1c�S(c'�\�ɏ	)����a|�D��Z�X����椦8�ar
��\rAN#����p��]kyK��q�'���T����b��9�d
�$Km?��[y��y�y�d��%��6��
+��l}��#'ESfL�!af�/
�g�8�H"�����j\Sg���Wkv����me|4�^1� �c(\F^&�ԲEq� �8*<�@�r99�y��ȫ�����P.��:������_TNSNk%�#�F��6)�s�LЙG�����+�8΄�Jm�l����t��g�^��t�>����7_�៞�~����O?~�?��ow�.[~����w{��Ѽ�:�t��V�=^=n������ן����_��������"/W�]�tk���������듃����E�ן<;���׏~�mnׯ_<y�U�w켦<r�����O1��=}xr�p�>tկG���{�8\ͥ-�CՎ�2W���ڦ�
8Zd�\�@�˥'.�Bi�2,��|���©E`WM:z͎����*IF[�G�c������ݰD)Jͮ��8ȼ*76C����5�3����:!�t&.�2A �\lL�ԁ�B���\��8�q��8�f��]��Z���3�UW��l+S�0GL�tҡ���C��KD�!f5�g+Τa�%�b����z���y+)Z��˨G�i(��9�g�8ir�h�0�w.N
�1C��Q�B���9�y�	VC

�C�Zԧ�?�q���;E�d$X֓NQ�7��»��8�H0�l�}۲ #o|�$M����h��!���xv��e�<�Q�G2#c����Y�,A���$oy٭3S0���؊�O��H.}��\3д�b�3��_S�\z��\��FV�B�O
Gϥ)��n�[gL�9��r�.��F��w���� M����q2�%ԏ�lC4Yd7G��\�#��C��l.��������E�f"v��(\Ur5�T��f���S�ڦK��D��h�.
M����G1ԗ������7� N6��K,8аf��C��҂���GدAU�����r	i����L'q`j�8U�5����8E�ɦVH�'�T�*���H�v%���VasM
A��hԈ �B8B��2�� b�+�NSh(V�/���h�z�&�+��,�S.*�)b
��A�F��C.�0�^$Cj��������\��E���1M}-�)̂�Rf��}�Y����xa��@v|�Ԇ�=|����@aN'�~��\���8�d7L��V�S%����Q�f����l�m�F���N�?��C�5�KVߡ(*�fdX��ԦT��46����z8P˫��e�ò ۗ�B�b�^� {�����-KG:!�E��,�+�, $��K9A.��0ۯVI8Ps�5|o��C1}��HV���̘xف�(��s�2y�<���m��v��;\�s7L;�o���q��kO"��{���ʥ��/#.>��Wӎ ��ε���]>5-���Nx�K�Ǔ}t|��e���Í��������oI^]��o������~�
p-�{�㛦�w�T2�]����"�����a�z�M�5Nߧ\�O�A쨁|<˪��[�� w��{��=���a��/m>>��>�f�|�����~�f�v6ݵ��FO��6�燻��?�ܝ=�on�6����a�ܽ��Ɲr����8�n���oU�9<;ٚ��#��o�z��-����Y{
W������X��q�e�1=��8~���1��	��e)�O�H6���k�aj@	p��å	�$s���B�O����R�8���e��]��J��*I'%���W�|�S��v�jKD�K�^�y��)»�䊀�x�B�4.��-w�����K'�8N��	R��7�G�n@dog)�\4jͅ��U�VRHE
G&���2o�*A����� a��V�:]���-��*H⤐[+��p���pQP)�Bɠ�ZY��:��#P3�\���!?�{x�\.�5�B��
6�%&[lm�"+ț�!P3��>�Ѽ��@̼��p!sX�!�)wx4AW�h�'�F��T��V�Z�C �]&e��fQ�r�$��^,�ji6�����GY��I1JgX.!@� ʰY�heD3o�Z
�\!��pz-�ԭ;���Or]�o�ql����nN;�J�Z�^"Xb�lTi�d�H�s�ʪ&C.�M�q�.���2��ZK3fc����5:��U������y�&������J��������-i�O�߽���_�훿�n����/|���~���x��٬֫��;?6}}��٩���/n��߾;����������}������¯��O��ɧ��\�􅞕;������X��\=u��M��������{�>�|�����t�M�l^J7�ks�Pf�f�-H��`a;��6R_H�Y'�#\�(�P�)�"pC}�NB���,>�3�s�����Y�#&K��h��)C6�b�g0�2�1�Ly3�@���	p3*��g���+��+)��5��!�W	�P������č�,/��.ܐ�eT�2�O�W�ꓒښ&��c�L-����ግO�1ɛN��Vl��&���Ȥ��q�R�D��y32���%J�`>w��h38��i��׸&�B=q�f�����7}��q�*�!<.9~� q���%�$�&0��-#W�����,�,G����Ac����)���v���>rb*@RY���Q:R����,�I��t�
/�1QLY(�j|�d�c"���2:��#T�@��\j��]���Od>�����O~��;�_>?���yx������⻿�]}���ŕ��\�����҇���ƹ��q�0>CZ��ɠ�������o���}�c~������������Od�p�r�S:��Xz=�x}w��7�w�
�C���i�_~q��<�_^��l��p|�u9Z�1���m�N���v��q�1�eC�Jd^=/��$2���S�/�Kd[�E� �Y�4�d�p4^u�2�DF^@�0S��F��\�H�)��=5�Z��*55H���8�#�tIS/�,�k!��ň)��)��t lM��_~6����p F���W�)��'8up"��&�aO��mRp=)�Zv ���L��J
ԗ�QT�S�P%�g�j��MCM��l��54"�\�[�T�'��%Dl��EQ����9G��)�#f�&Nj�N����	O��@RD���Xn ��չ7\���^x6��ɥ/#c�C[�\Jb�� =����8�!\F�R�X`'a&ek�̿C�ÑKѰ!���1��9��~Qم7����(*Y}g�VC?���6i��q���-���z�M@!@�(G�\�Bʎ0r|\�Dn�{�T����G^��	f e�!�dCd7Ԓ��BC=~��ZRlF+�m�Q���߲VR5�2�
W�J�S�B����U��ټ���֊M-/AC���i��5��y=#�V?)�!o�a���!�
!��Nj쩉��"O�p}.����*a�]��ڌ-�aSkX�>e!��G����c#YFMl��tD��4��)`*X�mBʫg#�bK]��R�J_.�ROW
q('+�pjB�� �������3)�,�W��P͆ҕ���Q��J��(ƴ�D���0xeW��BK�3�p�ֶ�D��*I�U"`
����f���Zm�X��Me���/Kk^���	�U$�1�詉bhbUh(j�l�s%Ŧ��V�1���fߋ#!�RƜ��kF��1}����:��!�AAT�v�A$��!)���@4��&e�!�V~�BN%A$š)�����p�bg��UU�"��!�>�(df�c��>R�y+3A=&ٲ�����j�N|����{F�/DlxLCKT�p"�Y*[�F-�WO+��G��PC�-��Ř�^���fǌǛ�H8�o!Ж�*Ru�^+��h���ީ.������۔���Ũ/qz��3���Ρ`?v���}ץJϫx~|�W*W#ȵO{�O�����U	H/?<���V~�e\9=�nU7C��n|3�~�t�g^���K.�����=���\��xS�sI5=�z!mv35�`�@qH���&�"e
�t�L�q3~@�WJ=N|[�����wo}5����.��|rz��>}��������������5Ue���8�m����7��m �n�w���_NsY�l��^�y����=_��;۫���0;5wDu<��m%�W��#��ٰ��)�!�.;�p4�ֱ�$��]�mg�(oG��Q���z���"��S�?f�a2��    IDAT�/����5G6��A0�@�ey�oM�jy�e�Pc��+��p��R-�#�傰���'�#9&B5x���ژ��'�iP梀I-Z_,��TP=�z7FR���9E�#0/��l\͑j��k7�+��@����5�55 5�3U[��r	�ˈ��WR!l.LjlI�!>��d�%�f����
d`�*]"eD�[o3V��1�������\x1���=��l=�������#�U^�fȫ1�m(Vc�x)煴�� ��(���E9��i����#���b���95�Vo��-�AHߐM=Dq2�5"�Sʐ��Xe�d�k��lg]�.#�(��G��`SC`ﲷ�g���2\�&@�8����矻/-Q	,����Q($��c,��	�t��b���	*W��q��hC�mƚ����Ԅ�m��κ����ix:�޾;�3h��6{x⋓O�r���������ps��?}��tu��=s�q狋�ƽ�.�����������O��}�����ѯ��Ϟ?����n������؜>m��4�,wW?~������s��x.�M�X��r�׽۟�+}܋���~�s9���E���R��-�- <���m�����/�
��M���!H���e���v�s;V$¡`�-2;$2�F���NQ� �)��
$�ɝNL
���Y�C�L�A�O��ԁz4�FP���7�I3)����Lj���58;��a'�h�e$2]坫�0��� �Z�ZR՟&NT�(C!y	2���ƟHy��ڌ
�P�R�iR@��U°�1EQ(^l=B"S*94-Z}e;N-Z٣�>��0 Y�L��!���Fm�����x��1 ����j��#�<WIv�S�\
#�eR�U[..�Ѧ�&D3�R��a�����A�쬂�l�,(ӃZ��ݯ� 2_�_�*%VZ�*��=�a��\�p���\�S@�Y�C�毱�,��&��'*!I!�m����@���S�\�g�^���x^<�<y��O?9Z]~��on��~����\��߿�����5��K�b�I�����I��ȥ��}�����f����w����;�C�n5�9>9�:?��������?�\���W}�����l^�|z����ٙ�:�^�^m�}<f�e�?�<_����닻����B*T]�c���`;�llGx���D�V���zC��->�7�m˨![j4�����1�d�<�Pn��Y4"�T�qA����ЙՆ�q��C0��Ԅ4y�����br�Z�@���Z!�L�1FY����ԉ�GR����.\�HD����L�7#x���Z|�p-�>��@��1��S�WORlH�e,K"��)�s�҇ ���s}0�����I��k	���)��?�d�/{��WXR<p�4Uhk��K=��E��OZYf,f�E�E�a��I���a�g�83����a(��S��ߧ���z�%�ˆDK��k����Uy�d_$?<NS(*Qs%g:!y�RO>�rU�X�z�Z�e�!�ɋ&���7�d�+��S�:�V��	1�-���#�g�*�h*�����g�
�b�ɕ�B ����L.�lٛ�!��[�f���#��0Y���BQ�f�,��)�����#��T��/����܊aV�!�B)��E�FnF1���g 4/���g.�W=h��']w�#I�e���5��ܗ�ZX]��p0�ÀC� _���D�$��ê����ɪ�Υ"c��|�O��!m�J&$��{�WD���TM��T6���bk�*6P��J')�6�⭀b��eG0$_O0Y�� ����!l�VyyE!������2�Y�_c#+i�B��ֻ��48�!�䰁�U�7$h.ф�1g=)�[�6�� .@ѿ�+D�s�XH)p��
��ն�ߋ���^��R�v
�pM�-�x�*���px�r�6��b�Ր!pr�^��֫r�2��4U����UR���~��0� �Ɔ���2�3ԓ1��~%�2D3\O��x�,A��GY�y�J�+\�V ��*^x`��6��I��Ջ*�2���<��*�͘Q��q��[��/<r.���
Tsv�h��ˎl;Fk(\
`C��&�o4Y"�3sA�4�R�g����R����I��\�Ԭ���{)�KA
�G?�0�7}2J�|���
4h^�g4e����V����z�\l��܌2z�$嘃\�L�P��(�����j�rIΛ'E�'86os���|D�x�:�^�}_?�y#��`����9��ģ�|!x�c��}�q��8{8�G���x�k�}\��u`l���ԖL#l��Z� ���D���������x���y뢥���c�����͛+'S��x�?>wsu����݃���˝�;������/Wկ�u��ǚ�Є�+���?n=u	�c���y������U�ʪ����c����2��o6n��v|���<pjw�v�����͓��ýq��z�m�.ɺ�s�����L#f���\������h����G`��aԷ���`ۚ��*��n�fǷ�8�=gl�w�r66$A�}��K��p��p͐�ޥ�O?���#<D�X�6��|�,���-�D��,{%�7C��f24HQj�bbʈ	i�FHP�1���J	n���b�I�l�u��m��]����,�'���闩u�`[�.J�#�H Ѵ�齜y-�ted�R��p��^s�Dv��f7�ӑW��*85=!��H�HJmld��a���8���t��R0�[�b�5^�����J�%�`�C+/�PkM;��/iQI%��d�4.�&�h+��ȈY����T��4�pUA4��LK�!#-P8Ôy�B4�L�� �f��.)�J�p�!HĐ�ް�����l��*����l��B-f�y�����q�o�X��єB����ՓW�,^8Dҁ��15C�me���bMN�d5���?������Դ���)��́*��eB5��
uM&ZE4Q��EMYH8�/�����!?g9Vw�^��}:_��u���ʗ�6|�f��xs��ށg��Y����p>��>~������������{�g0������:�x�vu~��d�����������'Vu���7���\���{{�u�d�����㍇{~���r\��t��'	�]�m��������96���qr{�z��q��.��?. ���b�k�-�f���[F5����8(����~yØ��po<hb뭤&�a��:������/E��_sqېWo�4�R	�@;�7<�<�\��m�nR\���/E��ghp��t�Hu�H?��䭇�e7l�!\��¤1��z4C�#�H4�@=��E��\�Z��?/�B�B*5���՗��5�z��:s��	��d�Wژ��kH/��tpr1"�/���ajlQ�2qQ
H�	����3��@�b�«*q�R#�#g�h�[C�!۲M�h.\�&�ʋ)�L�%;\Ŧɫ��h�a�7T�zHs��'[��U^v4�+Ne���;�7��r/y�5Q�W�f(�r�l�R�x�h��7t����84��N�����!ZB�ّu�h�
�H8���U�X�fʥ���p��g�4��m(�@Q�2�lƦo���w����l���އl}�����/�����?�뻛���������y4��nz���x ���������l�gϾ����ιo����#!�/NN.l����g�|���5�>���s�;�w��Ci�t��G�/�����Ǉ�[O��짯~���������k߮ww��nv�<`�Xfdeئ����R�:��QD�&�ǒZdv��-H�[l|���Ϊ�5!6A�*��7 :��}cfIJ=�%PIh���D�d���bJ�x}4��B ��*Kç�*�V�!��>���K=9��p~DVy�)�d��S ���BPd����Y}�?�zd�DQfk�4 �t��h�*��P�^=8\����M��lw�$�����#ML���Y1\h.�~�� C�e�=�f�"����S�8z��ylt�	�ԌY���K��/�Y?o�R����������m���ݞm� k������ o.y�k�6�b�h�
,o:\�p��Ŋ
�a����N��>p:�� �-��*��P��_��af�5�A�/ja�k�`XvvC�t���
kRI��N�ȕ�V$Nk.�+�G�eG��ٍ��-���'������;+�a7d'�X��d)'�&�\
0,��gv"�r���2��KS��h�`D[�j�-���`o%��ՙ�:����0��MP3�҉�"LHQIrA�Mx��˛~���, A��5�D$��=5���S�a8qٲ��lF�񫹤%B�����S������O��ĳS�T�~.r��!�f�"o� ��D4F�K1���xv�z)e�kB����N�	���M�!}C�F-D/�^k�\��4����X��i
Y�{���2B*,[TŔ�S��*��>\ ٤��I�FGOD:8��ņg� ������3�\E1Գ5ʭ���tp�6:A�+&eA#��1�y�����F֐q�q���i�JBc��\h�
k}���[�����E�w΢���-a������րD lF5�<�1�Sh.�d2 ұ5��4_�g#h�5��������,r.l��,�b�*>Pc�Uj�����},��_�B�'J}�Bx5d�V䔪�@���'°R����L�'e�UU.��ڟ���g�9j�9�Q@�T��*�5�ODv%�zΜ�΍�7�$�L�PzN�_|��Y�|��E8��2��\�}φ����q��t��:ll�dw�y哪K�������W%�O6��s:��[�u���>�`'����y}�}w�*������������ó��ͻϞ�����Q������y��ѓݣ��g�N�.�F2~�RFՎ�L幽rB�ޯr��ݸ�TUۻn�tA��h�#�t��ҕ��b<ЅGgo7��};���ȯ���89}�z����gw�?ڿ�S�OV��^�6������ۭ���W�g�H�3�}�D��o�6+�<�x$�׫����o¹Mm5v����mG.���jmVC5Qv�
�_P�Yb�FC`5�Xϐ��;��8�+�ؑ�Kd�v�a�3i�D8�ts�{�g�z��~�U�KScO5�4��Jj�1�ǲ���(�����;�r�����kl�!�5g�����N����δc�����iv�uo�Ry��p	��/��F�a¥Ƨ'�� ^.���q�&��4\w@V0D YLʕ��S@����󆗈8�
�CZ"'��G��Q�P� �@4��F(;�\���5"�Й�&�ᘼ��pv���P�dz��1�5�)9�a]��z�e��:��5k��)hkڂ�Z48C�XpC�N��B�a��p��em��;�(
���A�%��գ�D�Ǯ�Ĭ$8'lgvnVH�%�D&VR6h[�>���TmӔE��=ːTv|.d�z�����R��7�q�L
:k=��1k�A�xR(6	�D��E�b�!$�R5�+7�����N_1Ƌ�g�.7���Ǜ�X��jA?m�jw����Ww�8��ۓ�ݍ�n��:�9~�ӟ��o~��k~����?xxx2~H���˓�k��{�Q�O_<�͗�?�f�����ӛO���^�:�|�ѓ���S���l�)�훫���\�Σ���20���;�h��]�S`�^�^g�_��ƺ�i�pl�� ֧m o1,&���nSu]ӲSt��p��}ȶ�����Y����	�z��6@V��S�������g���i��C\�v�e.�`oR[�m!��zC�R&���G��l����2�z�Z"���;oCR8@�8၆�\!q���f��t�j��/ߤ�ʁe�6�&DR�zay�yK�0����9^�XF�EQ �#W��
\v9x����,�X��(Y�)�1�R)k�����	��Dx1٥kX��]Ka�m�S���@jbq�����k)�R��� 6�Oe`���u.�2��s��A3L�!E��٦�4��pz!�ԻH۴�m����ȼD���z��gW��IC�'V��!�?�/��&�Y��?;�!�r��kBԦb"�lj�� ����p�%���ih456�V�C��r�<|s:~3�͛����/��O��=�>pvyv�g��3t�m��ً��=���+�m�l�޺;����,/��pr�ȯ���o^�\_�_��������o=?��豩]�y������ݫ��������V�9�@㣦�`�������|v��ϗ�oz���J�۷g�q,5)}�4;Қ���o$Eô��[{�U"�ȉ�(�'e^͟P�8-2q`{)dR�����"���2f,��������g7Dh#V�Y��A�7dse��"6���pL-�.��(�4�P�:3�b��p�8�P3ęQ�`��zLHM������$nc�ы-�\Iyjpv���GD0�7w;F�\��3>�ƕ�a�@�z-�ar�Yď�R!�Ԑc]�a���) M��`C�jN�0ٲ�iӄW?/P՚�D0�Ϲ 4�5�4d�*�(ei3#$2;�@�s
�4�#$���n
:ꧠ!���aH,�,|���\�v|}� 
�!X�#u���kI5
k"�4}L}Q1�-����c���ȆqM��b
��kᒎ�_�xS�W�ݯ��$�Dl����Ԛ&�A�ˈPIl�Dq
��ȉ�I� �\7^C=�9"h)��"ռ����q���r���.�p�8��\%1ٌ�Y�ጲ)����*\�)���ґ&�.��˼
�,r.�t��B��J��s���bz��f=��u
4d�K��;��U$#>�jg"Cv
�k��$B���9W+S_v{c��/��ԧ#�@{nنt�38m!Z�zd�SˀhC�!��[@%�Z��g8�B�`�2,<e^R��+I��f[p�0�Y3���p���fH�����sih�\zR^��%���'���W��f30�!0��uA�^m��E 8���Lp�� S$��kt�pM�XSN��Kk��K!&LC�w1�3c��r����* º]���ֳ\���W9[�V�y!�+�ά0�ɏ�l
zd�f-��Z�v�z��O3�NR+/�f��Z6YL��&
�t���e7RFFN���j�N3b*���
��l`��'����jKԚظ8j�el���pHk��<:�W�X���C���>���UԔ����e���An3�$��&6*������w���}7q�U%����n���� =gU���=>pEr��W��/�7�g�~����Z\o��c�nߢݸ�jU�s�Љ^Oj��0�t�i]^��񻜞p7Ξ��zჸ����@<w4��}���u�_�ںr-�pwo߇�q��ަ_ń�>����5LG �]D�Z��4eO�sau\`��o��븮���˝~�E��;����qq�ֽ�G��!������s�d��u��ݮ��o] u��";	~����;�n56Q�)Q��&�]3������[O��v���1M����Vfl��i�osXv4�vapi��R��۲�h�F�/0o��Q���KD�:����`BLSo������Ԫ�Xv�2	@)�dGf(#r^���g�̆g�k���J��e���e�ƾ�ܦ儒.�gLӂ0��_�aj֖���t�Dx��N�(��,m�R�ESC5SА1�0�G��W?�B(�%��p�)�W�z�h4[
qjJņh�f��q�&�2��j�S�)� �hi6���]Ƞ�Ff�O_:�զ�U�3W*7Y+V�֭,I����F��T/PT�U��#�4��L�����QI�Aj3��}�C�LG��o[��xi����֐�LmH[�1
�bmSj@�ԧ�&�s��� ��V�-��S���]Lo+�n�U����D���ѷM
dM8}FS�7)F)p�8B�45�z�LYv�%�Y{E��믿6dC39�"    IDATr��/��q�O 	;6!�xr����By5d��h̒Ec������<��r.oO���K.�y�\.vR�0��{ޓ�O�\��w��<�����ç����/������������>���7W׫��������������?���7���v��o~�}������?����������'Ox�����(��{Lh���#w�θ��͌n|���r�+�W�G�＇y�K�t�o�X&k֚Y���ű���V������?u�6��-�+���ۺdmr������V�漘��!z�����D1ѐ5
�h�8l��n�`��R�D��lR����x=�b ZE2D���MA��oH�jy�Z!�q �VBG�n"hZ
�3��!���aY��3�T+�+ټ�V�$�dK+>ۏb�fWaH�)
�d[U������m�~3�4��r1�'<�^��k���Wg4/vÌ9YCRB³��֯�(̦�1\�^�����pi�S_��-|���Z������|'B�0��v�6�b��[�)�7Mv^��R��,ǡ�K�^����C�E�q	��'[���1g%��ӮBVCs�t�As�h�\�t,���Nz�}]����L��C���b��� ��MOͰ����ZP^��\��~��w7�ar��*��y�������7�.�3��OZ��|�{��G�~���7���G/�.=�ǵԱ}|�eӯl�0+?z{�k(��w���l\���yrz~t���J��~���l��|���w�ӛ�_}����/=&����>|���zu����_*�~����~t��˗�~�l��fw�s	|�rA�Y�EĶ��0A�l�z���\��e}���@�wd[M�YO64돯�#�>D�}��l���.�7^P��h�m�j���,Rh��� ����W����Y��g@L���N�}R��Ub
/�3BH��]S��������ھS����h��0H�!��T)R`�3��1��bF��7C���j�t��!N
qxi�ف�d����x�ˈ����(A�HF���ځ����a�z=D�!�3{�����oχ�L3��WS����	1Ԅ����N���ؑ13 b� �ڰ�Q��=�5C=�,+#\�z��P�3b��Q��8�Gc�����e�̋��Sx�I��e�p�SGv^}��b�[.6�Y#�A�c�F�(}j�� ^������w��Q�E���P�&����a 4���.�(�65��X�%�ȕ��B�b�6�x1D�4 ��5�
��n�	LM/����'.D".ʥ�3��)v�_h�$�7�ɨ��7���6t���b�_R�gT�D2ʵ����)��!�2F�4����;���9�t��y-�-HDkF���z!�l=5�%np�%�1�TCd=$�Y[`|2f��&d=WP�)���/fy���@C�!z-��2('�g��'��D�I�E^��m �V2�#�t|�o�:��U=��lF��*lڭC)�)cj�N8Z}��~�R�U������h�}�3Z:f�8�T��3�L$\�8���f��!�D^>�^��3�0(h�A����
Ѹ M�N-D8#d��Z�@�D��H��`QSM`!3��j����jy�e����N��f
���D5�d�+p_�Hk�F\��gj`��k��C*o���dgX�);ë���2Rk8��J���
�Yͥ��ht:��(��,�"��E`����U>�Y��"C|&�����!vfH������d;�+�w^�j�����e��q��2������1���3�6�/-�JD�)R��!�<�v<E�jܸ4x��긘�ɸ�皠g܍KwV�=��y��&!O#b����Y���ripܝ��G���j�[Bn�Ы��q�qܭⲫF.�[����W;��k_���tIt���s�//W~,����}�w�:!�Lo�NL�;8�7(��ES7p���屸�1W_W��u�K��7c�q9tw\][j����w��7��{>�������g?x+��7_��z��zuzwy����K�F��q�.py�qr��A�ݴy~�����y���������ҩ�i�^
��3�v��+���������^vW;	ͼ��3�����!Z۝��~��ݗ��M�.�B��sG�*[H�%�踴��@C�����#�9А1��J��n"��aK�U���@���vҩ�si:D�V�!а�G��|8o
���M�*K'o)D9	C9�fԖ���{�) ��%B&U.
�ʓH���G ��r)5 CdC6���(C^���c���@8����T����EM���L�lk��x�Rmr	4D�k�zCd��Dn.s�YR.�X�4�p��x�W�a�h�b�ɲSH9����Wv`�g���2
i�7t���s�?��
q��b'�\��0�t�/��u���x�Q�p��N�/��򫯾�?��/BۮWA���x5'��mviٽ����~投J�4)�2j�H��QC\��S�z�:����+K�G�.�)�w����t�ɪ��0��r�*%��^����3�Sʪl\f��-�B��7v� ��7�eS#.�9퉳N����7Ic\�<���@᎗�����vW�n��ӫգ��C/����/�����|�p����g����~����w��.<Wp��ޭ�/�N�}{q��Ͽ�?n�����O����G�^�_��}�?�i����������������_�9tH�{x���-�_�e�p]\�wUt�}0.M/Ss7k�B�5ˢYIo!����կl'k�5}[�u6d�l�^4)�"1�(����\���=/�ǚ���|KH�P�����f���ڔ���}��XY
�C���k��&E�uZQR��1�'˫q�7�-E�`, Zʆ<JZO�,��:�a5�n�>	�@���k@F�h��-(��B4��#odF{C� 
��"P�Z�\v'^�m�����
�ϗ3��
8mH�hM�T2A�����tR ذ�0ܰV�4�C ��7#а:˘�+oj��f5�	����Y}��M�!�"�q�tB�����9��m8/�Pq/U�އ�T���Z�.��[x��*
(B��d@�Sy�B��� ׄ�T����m��wm��(4���K�-x�b3�v?y5�j���q@���%r����@=����=z�|���ѭ��͆�Y��C���ŋg/O��r������8�r福\������_�=���Ń'>�-�<pvۻ��ً�������]^��p�ݣ��>:�Q�bso����|�����>{{~r�:~���O>�z�#�މ�|��z廪�۹|��[���|򳟟��?�9;�Y�p����W{<�'������aSq4��`�m8��=���Ӗm�,`�Ɛ��}�Vkτ�!4��m�lQd�$1�A��(���(�!�j�5.=d�u7�K�x {*�
$B��F���/)�(C.�^���2D^����35M��3ث25�p�^���k��AAc��o��X��K��CC�P�!��
΋I�M�n�fR�*�F�1gyD�x�i���>WYF�Қ#�)��#��%��:�{�cE����(�p�yᤀ�Y����/D�Am�!�@8��S��%"X=�������z��P��Q��+DO�\�m�8gv.vC�b(B*���4��5��E���e��e_'WC��'XAd8��!����U%�)4�ʀH���������L)`��rIW ��!�L�`���xy���H��C��xE��2�BcD��D�p�%��л�ܵ�sN��)����C<}=�Oq��X�֎Z��ri��/�4S/�8!�xшO�J�m��;���z-���P�s���v�%��8���>o��T�Lr|���%0<��Bڻ�/DO����9�t"���f�&����P`8L!��zZ���S9�![mU�pf�3������LT:���	�S���z��s���\��Rlep�E⊇p!�t�����������
3&Ͱ����zn,��K��wQ�2���p�V~��d+!<���$�Ѫ�z�ނ4�t�
�b��ڢ4^�l^_`�pR�ʋ���)]uN�Q�� ����7��M9�(FS��,�$��Q�����45�
�k$"谦��)R~�8CnĤ`"��Ex(##�a	e �{���&E$e�6�!��^V ����O��k]�B=_�6��7Hm6 �FA�UxL�����"
a��Z���	���f�����2H'2>�(��X|Fe�ǈ �����Z�CO����¡��Ԣ�cU���u������Ħ�N�-����Y=MD
Ϟ�q6�J{иg��(-o��!%�[J����:%�>�������z|#oǷr]5��|�u*w԰��AzC���6����2��?���\����z���j�|w��r��*�[V\��C,�ҍ���jr�O�W��S7�ƹs����v�<u�]=Oo������ǲ,Oĵ;~���{A��i��{������[�e^��y����qlk�<�	V���>�����]\�\�~yu����B� gw�'חo7W�ۧ���w`ܘ�����Źk�7W�^bn����۹�4�k��\�{H������x���m�	�g�+��׉h�4
M��`���7��rИ;�ؠK�'���B����&��G��֦�,Sa
* �\M���'2|�\d���8s�]`
&��<5�T���4���yZ�q>J��I�@��3H�a�[%V��V���˥�R+�e��Ѻ��)������/;P��^A�Z��4����cT��
áM
"����L�zx;�a$�%�P6�φ��7RaZ4}3-!c�͈N���0�MB�M���D��{{Ⲥ��8KrE^�T*�f�Z)ʘ�jd��;C��Ia�FIC��'�І軷�&�7�6H���qE�O>�L�y�{o%e�5�Væ���mP��йӒZ�>Z���Bϟ��������-B:�[C����Rv�yn�.9z��N�^�Y"��W	0qM���R��?�+(򌕚K
�7�|����^}�g�}�"���*?��Ϝ��6񤗀
�
C/�a�(�ںX�Y�$��ZU�2�/��g��& ��;�m���!��v��ڤ���7,�}�����|���Ėߗg�NVo�����'�|�s}��ų�|~�w��Ǉ�����O=��ۓo�޽��r�Ce���F�a�w�G6�ܺ�|o�����W77�x�����.^}���}��������~z���0z��ZWG=���������'x��z����x�
�������O7��n;Ya{��}��[����l���[+��mׁ�eK��`��r@�+� 0\D��K��,�� �Rh��!�\^	�l�bI��������l�3B(3(Gf3p �
�USs�
�	Ѧ8005���^����ڸ����gp1�\�f_`����r�!\ϥ�ӒE��d��ZsQ�0���1A�g��6��}ì�5�^��o��
0_Q���e���he�ނ-#ou�T�\���c�]�)Uy���6�B���o���C:2�4�ŏiXxC6���q��� [�^���_��dY����������0=�������td��B���KgP0�W�)�*�0�kZ��9�h8l8[vM^�f��p��B1�$��C�T�J�:I!�ՠ0�Ws��5��/�K^jh�J��%��=Q��=y��3�n�<X�sr������'�_l�8u����Vʷ_{����3?�|��}{�*�Ǝ_Q��p�{V����-�u��Ý�7���͓������������tpt�����7�����=��ϟ?x�����~�OJ�Qsv~��:���:x����W���8~��'K߃u��펯y�u�T3�VL?f����V���|��Tl&[ͺ�[=���H���
��Ӵ�b��I��ڣ��._��eG0��Z

K�AY��)���q��H"�����z8�l�=C2��
�;9��5"�𖫂�B^x�Y*�$e(�]�yA��7�i�W���ᔈ�Q��e	[ �}�d�0�@:g��9���h���zysj�����Tm'�a�XKdMf���Ӭ��[�+\+0>!@^��lF�lF����E*��p`Rf
��`�l^�=]^b����g��
��H�!OD"v#��\h5^
��D���U�?l"IUsaW�t)Dn��?�p4y'��!C�K�Ey�+����E�j3x��f�e��U D�\��Y=�p���O.��&o�cCp 8�������� eQa����Sf�iE1Is�7) ��!������X�VIl"��M������]j#/PTE��V�t��4�#�� $Aü՜��k��F� �$0p�d�Z!ed7�w��ה�@jy�A��(Wʘ��5̤0!\�l����g�D�6MU'���I��ۆ8b��E�)�D��gx�>��1�=�]HO!�6P�g�XͰ�mXl�p�&<^���ϰ�@jB�Q��y�Ē.E=#�p}8}{ce��3f�Ș��.��g)�f���|���3���3Q̦����+{���G8�X��l�K�d�m}�!�!!��!W��@��ِ��X�de�ʞ&�;u�)��0����*E|�D����o�ȨH����5�0�X�,����@k��bO~
�hZ"�!�#B����6�G�D��J�9�,�N,�)2�^e�TI.��UeOΈ�7�K�=�r�by��nrAh�q ��\��
�S����#�ǌ��Q.M ����9�(�d4/!s��ri	
'���^,�4=2���yKd�;2��g��{N���G�S���񍍠Q NP�4�D2�8f
H%�'����km�|�>\�[I4�D�\d�Н�V�qs��65�3�-���n�/J:��l�3뎯�nm_ݸ�S1� µQWUM���z���KȥM�i��m�㹮��	E۾��ݭx��ٸ���$,}�ʅT��s˩��+Ϗ�����T����i<*�R��N��*mw���fv���m�[;�;��#���y������q�'8ݸ��h����볓�����\OT��ʶ�:9�y}z}���5��+w�xȂ�L��V6�Uq���^ƫd�o�e[�sŪ�vVu.��6J��a#�bέ�e��C�׋�b�-z#]v;��S���p�q8[
����N�9X�iҙA�ʢj@=�A3{�fm%�[�!I%��l���U"�ڲ��z:5����yrbe�#{�1̱W���L" qQhC B��I��Y/.�ea���/�ŇW?�\�Z=r�g  7�T�i�����U!D:G������ì���K��J�n��� �!���ZI[[{�R��(�/\��%5�E����g):&�8�5ip-D��4и&'�Ѭy1���I�Ojz3��M"J�Ed6 ��jv�Sv2��m�+X@6AYra�fFC�e�&@Bӌ*^FH�ˎ�W��h�a{?r���K�E$/�٤�R ��.gS� �	�<0����(�'h(
�N��@�^J.=o'�yC�$kF��~��_�8%�ӟ��JZO�&�:;ViV�y�v�����s>�\���ؤ�ʢ8닓K/�~���㲦�8"\�I���\��<����՜�qy�G���p~���g[Wj��X��7�ӗ����COp�دO���O��V�Ϸ�������?^��������M�B8��s��Vw���ӟo����l���z���<op�`kﳟ|��������
�?��_��?r \��;H��k�_}�������\�G9�:_v���Ifm�!6 �9z[�/�xlӶP6R"p���uȰ��]���I�����è�\�'�֙��>!5���,�ֶa��W�3چ����m>
p�̀ϫ�DƖ|����X�lB���5C�}6͡��`"՟W�4��LK�,d]��g�k���E$oL:���^��y�0�ҫX/d�`�m�)ׇ�g�ة���U�cȎ�P�g�e���    IDAT7�So�$��l"� v"�!�@JZʐ})ʥ/�����,l�h&+SϞ��� ��xY�2sR���v�)R�d��x��� �)|6�*���5��'(ҺUU"@.k�U������+�e�
b��V��E]%4���	�,\��m��!R(IϦ�Y�u>o:�9r�-�F��qL����d7_LG�J�,܌Z|�\��c��]o�fG����ꭵo��tf�v_u������?����ߟ_��y򝘽c� ����9z�������/7��ݎy{�����sx����7B�����������W�@�s�wu�v���ٷ������'�����px5��zso|��{����\�;9y��Ưy<=��|�����c����3��4|䳽��iF�DFg�����?WY&ޖ����A�x�q�᪒�[���G�5&��x|����e����|�e3�M�	6����OG=�n:��)��O}dHR8pv��l�u�	r�=)VI�)@I��z�-�!#dc�ri�6�h�yۇS8k�]׉,�i*8�~�#��l�\�);�fL5
Z��b�s���(��5�V��a�!D쟁����'�!Dϛ�@�)7,*�\��FJ ;m2{)%��f�@�֖ʨ<�0�ʘŔ%�\������x���R�z��B;'.�Q���a)�hS9W`�1�f1�s1��g%�M��S�=�\E�S�֕�����ox��g�B"�?[��5#�f(V���'���'>� ��7Ch���q[O��&W���3!K�BA�!<2�,����#�!��(�\U�D�,�xR�U���˅	� ְ��"�>�D�_��Y��hO�UHWYF��7MF6���R�΋��8�!��Ҷ� �\
`�� �W��z��b�z`Y����QƩ���H�V�Z�,�Y����GK��z��V ;<}�[C8N=e����!#5`{P�,��K�O'[/Q�1�'��Q�	�/C���7$XK��Glv���E���|���	��(P!�ʈ�k���!ZKZ8�lLvFL��8W�BA4e�4;+a�8q�L�����O'Y
s4�T//�&V��×�=2�p��xS3��)��t��o��'��d���٢�yi�WRL^�{S!���4��(!��T0�ڴ�1�"�N�RT���S�PCFh�b�M?5q���Y�µ�A+��+0��+Q����J������#�����ke�#�ZO�<0f�޳f�>��0۔l�b����	����3���;��@�0��a!��K9�Z����gjFQ�����N�\���8R���g��ܜ��Y@��U�Q�B��wI�"�ʝ��e7k���g�.;�Ϯ��CW5]h��).Q^���S�l�}��hќ��v�qsc�^QW�ƽ��o|]��]_���8���O�Q�֒����;�>^��Y���Qx�}�;.���M��?�i6���n=���~����wNپ�ٵn"���Ce�n91&k�(��ź������S�RrYb��z�޵�˞���˞o+�+���/���z���@�u��p��$�l������l����G���ua�tG�n�����S7l��r-�i��K����-v'���"����}�!� "\�{��6�z�>�P_^�M��%ٹ�O?�ԉe��8A��-�K�̫�꬇�!C�z�
��ևԏla2�+D����Q�pm"��	��avhE��n�3�-J_ٌ��a�a^.R�l�s-�f�EG�-���/Kk��Q�#0��S�6G3""/As�Ԇ��o�Ef���3�u/���"s�)�	J��(�[�̥�2��J��Ţ1�ou�,se�(@�_k!�����r|�
CLP%?b�����!��p�)Q��XN[$��*��_�̀��M� � 3@̿R�!��R�dk�c{e�SCc�7�R-u�p�BZ:�!D�m=�MJl�f%-�}@/�9���.%����lG{�3��.uu��R�i���d蹄땁���W�JJgHM� F{_"W��a����|�;�Av��&g���?��9c̔MX����$n&f�kXK�r�@�]�p;y4n��Ø��e<���OI��{v�y��������/~�ů>{|����?�nm���y�:�|���������?<���f�����'0ܬ��=y��?�o=�;���￿����OoN.ow7���^���/���_>��ӏ?}��'�?�xo����o���^���l�<�o�۾��h{��!�y�����i��?A�{7��mYӷ⭆�lCZ"��l�h3��Rl!hB
����w.Kg�~�1��w" �6��x�;/���F�_R�@mY|J��MF:Z􉣕�M�t4UQP���^�8N[��@�ә6���R<Y�jZ�Ĺ���BT"
��\zA�B�Rv!����YyK�(#��'�&o������4���೙��ұ��:��D��O6�h��ժ�_�1#5�O�HG-�^=z}��)WL�{r���&bwBָ�ad�N}v���_�	�\U+İ����-�����0�+�(`���t��pF"���G�/dڼ�z�&d�����- �����j�^���4�W+����q<�2"��Z%#�Ը�(�ʆk}Z7� d��T*C
�T��[�@�/;�J��f����a.�lX��v�_�Ƿ@.��V
WQ���S�_k�ڽ�`�{�w�;�w7�G���ۯnn��uuys���'?�����nxD����ʋ������;�{�ؿ����/nO7/_���{s��>�[ԏ�~�_���?��總#wr^����wku���m>z�t{ӧ���G7��޾~�������������<y������ͭӛ���������b�T+�^�,�o�B̗׊Ysˢ�Ѭp�Ik�'�G�qT�0IipM߫����h�3ޤ�ky�+)[�FǦ�v!�@c�K�Ȗ���b*��OM����C~G+D
I�b�Z��u�fxQ�A7�If�=��EI�(��2ɒ[�k�Pc�48�:�g��z^8>�\� �A�`��d��(�ݐovU�8�R�R�W �m}8�FX�Q�Ckmõ�\���i�Q���X4F'�����1d'B9Y���y!3�Ax%���ɖ��_82���b�� �k38�L���NM�\@�U�"$�!&Z�fRCx���t�2�e�F���1l%��M�����W
�T
S-�,3�Բ���ު��n�������ib�瘗@��-/P�K+DxX�JE�Ŕ�7�2
��+8���l��I�z↓�`�ZHEB�UXh͝7<��R�2�^��Z�RT|Y0��,UX,D9�-c�D����3����J�D���RGƱ��р��t zi�	�W��8p��3H-͹�$������o"��\LR��9����K-�A2AH���O
�i�@Va3�=4�8�W�B=j+c"��\���A�ZU ~�X�+>�(.H+P�����R�	L'�83�.0��ڍ!��c� ��������Q���aQzj�6�2��\��>c!�!Lh�4/�T6�TF��q���6M^
8�2f�\�H�.�3d�8/��4g�p��t�a�˕���`K�/pH"����>�,fYͫ2�����oFl��@�����z�
���L�M)j/��� v���&K)<�98�l���/0Z�bfpIm�����E�h�z`�ːH�!��ШeW�a��l�E��Č a�)�!M��͚������x.����dTSk8Nd�ٳtp ��4�Z8��OQ��meI���R �lʅ�  C�\T��J�G$�v"���d�V�>���@ʥ����]_^���r������ )���z�����H���L�J�x��9�wK����h�&��G_wR���i[;̦/���-�2��.j.yz�릓���"��������/v^os���顈w��O�vu{�qp����Ƹ[�W�}�޽��bϠ���7wn|���B��uy�f{ٗ�3���k��x歃��o^ݽ~qr�r���j�]{���xz펛j�:�q"���з��ho���Ý}�N��/��ܮv7���l|��8�������=yw��uq�����Y�ۺ�߾�j�J�,����nO��5�t�F*�h��=�.������4M�X�e?d�";�=e=P�;s	������mn:{c?���#9��"A��BSU̔���,�M�8���p�_k�L3d.m�
7DP���5dsU$[ �E�^��2�6Y6�Bq1&X����0��]R��oۨj�
�O<�B��ճL_�l}�ة/��>�%gp���a�[g"��*���h(0e}OS��`�0	��Z���C,�8�R#7�K��B"k�4�'��U�x����� ėky�}hE�o��������z-�k���ԖM֐�\zHk����ر�)�ҫ![,o���ȼRāKӂ<}��d�*�3�=Z�0�d��#��7d����B�*�pYO�O�ͷN hh��N�"��R�(���QRdͩK�I���#%��0�5}�f�<��R�3#L�ʋc�;����_����A��C�;H|��?Y���h����D��PB�r�h^y���)�u�[n�����K��1�%�����������NL��|�����?���t������7_����lm�۟���>���Η�rW'�ׇG�GǏ6��=:||�q~�R�уÇ���{n�y����k7�<}��h����ѓ����~���ᛋ��=�8��Zs��=�}J��W�go=�����㧏��z�I�^>�ݺ;�߳�:����)�<�-�}?��6s�f��l�[:���/-�1�g�?ںRX^��&�es���`P�Sh#2�"/�QhY��!k@�aS�sq^[�6�Y��%�V�O�l
yg��#��Iњj���l��D�"��ZQV�����â ���B��?c@=\8�,l=[+�ٕE/���-6\�XF��\@�ڏ����1�v�&o!��X޹���z���ڽ�RX��f�/>���ä L�\f����K�aA���=v!�1
�.
-.�� �`�ky����M0fv"��h*�å�o(v*d��K�hB2
4�^G�#h	6�8����:�8 ��i�鵉���g�ﻏ[�;���HE�z؎-R��M�q�ZQ�QHT��y�@��4�Qͻ��\��A�٥o����R;$�:��_��b��KRk�)���,<����87o.ߜ�`�>~o{k߷P���}bۺ�-�O={���㕯�>{��������˘n�3�OJ�#������͉on���:�}��f���Ǜ�����ԃǏ>��铧G'o<�|lM_X��|p|�t��>�W��h�o����~�����ƕ��/|���ٛo.�,��g����S�4#ke�c��6�<-o.|�->�(��eX[��8�VR/#ڈY�Ig������������Ĭ�������h�S�yɚBrәC�i'h,�X �!�,�^_���ӡ0����WZh��8P+0;g���1�j�	�`+3�(���d1ęE�m2Cd}�U�-d�xw� ��5��D��1ԣ�6�a@���J0MU)>A�t���o:B"@���+�����vE H3��&ת���B�ѸjpF}!8Z���҇3D�	���l�"��M�!��ʻ�b�	���4SC�u�ZCRN�E~�\�x�h�W�՗�l�H��m�T��[�8�!8����PC�8�"k@/��b3jU�L����iHH-�jHٮ�ц�"��'�q���C��{�N^ޡ��LgD��`VC�#3��B杯��'͑`)�j�#���)B�lYC��O��~
���ɮl}��TLL����gmeTO��/uv
ّ'b�!O�ZA����p��%j:��f�ۣ�I��OC�h�`������K?s��GЀ��4�B�^G^��S�O;M4
��+�)�L}�����׸6�QÁh\t*�W+�>}��M9W��C4����Ή�y�*U�����&R.�DqUj!�8� �����Z�9,�-�@�P)�y7Ը��K�����q�qBpj� � ��/_��RH�4dL���(62�=�\�1�e"�e,��
����Z�������g�p^�>J +�����υY�޹���S�M'��z�~Tj,$2p�3D��'�g��/�i�'�f�M�(
W%��f,αV�6��J	4D��oA�s�XT�fGH�Q3$g��adI��W�^�E���ȕj(
R���_��M����96��Eô](�W�DK��]1��RlF[�.
���)T�@Q���!���.B��~ˠ��3�4!ȪE.�AH.�@����e �䅆︯�����1L��5^�j�'s�0>8P��r�g�>���˚����Tջ�M�Ar["cO�n��u5�r#H��#e_��;����=�l8��ǻ=_���0�������G֝�H�d�~�̈�k��e����J�] \�^H�B ���Z�� ^��!�g.{z��ZrόL���Y�@��mu�9�y�1s������T>~�yzxu�wi4�M�NJk��|z����I���_?�{�W�o��?�^�x��ˊ.����;Na���j��ރ[�n�6�~z���=f����ʅ��C?��u��nu�{�7���o���on������ON�O7G뽳�~��Ә�����7O֛O�8�d��r}}q}q���컾q�&�uޱ<����@��vlpY�}�8�6���u$����	��ز6� }��W��O�p��}�&[/���?�i��X;�>�D���/<����_~�,��e�x���&�PHepi�$�v�������Z�b�?B� y�akh*��5�f��=?�1D� ������?�BV4v��DY(:��)83��pL�q�ؐ�q̢ڪ°��ә.d�>AF)	"K��WR5̌,/o�[S95ù�hJ����`�Bָ��撚]:�$T�,\��P"�&#&\��5ӧ���@���ιT)�aR�%�)_�U��(��B�E��d��5Cs���l-e�e�|��Iq�tz�7eC_2hq��k��z��6��b c2��)�ڸ�)k�I��m��E�鋍���f��U��B�U*�&�(5�8�H���r��͎���X�3M���)x�n����O�;�c�f���w�.����2i�#*k��K.�W)�si�i�1�(�Û�u������w�5��ۘ��~P���.z>�Y�Y�	�����x����ٿ�������ާgW�ow><�5�q�T?켸oT.,�v���W�{��gޯ6�����\-�|�n�9����g�ӳO>�h���[	=|��z����}������ݎ�{�+��Y�n�0�����W��ov��rs���o���u�7{@�g�:>ZKa%-��b��\��V�nd�Z@L��hż��]�pB�l�	j1{�������p�Ҷ�(L!m���D$bK���v!��*��F�P�z"�����!�hp�e?����A�\��Dél�l��
ˋ@98�#�ns�p��M�t~����%�S/�A���C��Rn�k�b�
($5�4
�&jf��)�4}y!q��Z�J���(�'���v�4��/M`8���D$��E^�K��#�Z�zRH��x!�����#��I!K�`jsC��P��o󊢃��-���2�8&ج��#$%<��S!������?����ʛ5�I��8XC�^�S���a�u����A�D.�z�8�p�7��Y������� ���\�u����?\ �8@1�yQK���7@�Q:-������gr�|�����.�v.���_<�{�˃ͻ�������՛��?�=�?�xsw�-��q|tt}~�$���Y�>e]]�������/~x~��ᇾO���k/��O�}xp�љ'O����y�'�O�������{�x������k�0�ݷ�Y��x��h��    IDAT������}�K8����[���A��F8�Ӽ���j+�e5���\V�VnmC�t�� ҞS�)� �v�Q�� l�4�T��̀�e��� ��n�(�j�0���~��T�!^�	��X����3�+�O-W:4�y��,���鵐G=Sߐ����%*o�/���O�
�a�V��s��+�$�H:�-q�a�O��ŪS[�ƙ���e/jR0��T`3b�� �-��j!&�F���D�٪p����*]!��Ưdv�h�c�.���PRʘ��S���'�mX3)͘z6�6M��$0脤�M W-�rA���;�y�"T�~)��8U�8~�#�m����a�a��\�u�E띥X�)K����G�0ڟ��y�;ڰ) �!�Z����H���ѶNvN�!�[�����C�fL�BpZ
FT��B��A��B|�Yϫ1�u��/jzg�)�'>��0�U��Ӝ)��O��칊��)W��UH.'2�S"=d�0��p�����ٔ��D�b�1��3qjm�B�K�x/n:<��!Mv������t$b�6�/>M��6�-)FY5Qe�:p��b�[F����2�,��\۹�2�OA^޲0��V;���\�������	�QU�6��\h͋]1"Ajy㫍Q1ȼ)0�G�P �P��z4�p�]�ّ�ȥ�V
ÔϨA�.���M'ù�
�Ivᐩ`�B=�^�OTF+P�mq���Q`%I4� �� ��Ћ-{�
�O��/KNhx�B��[��r����������l^��q�������=��%�B�1ę�y''e���jm�ȣ��)��K����� )/$<r������Cx!���e�g�]�<xa��ޢp�m�vNSO�\���0�|��ϰ]�x8\B�U�Z`8fR�}��j�z�wt����U�t����g�-�@���e���9}Qͅ|������.?��-]h4?o�eR�&�Y��k������y�O��*݋��n��	��,�EP{ƚ}�^�V��`���t���b�Yϑ��V����O�tǽa��{��-�ˏn����8�{pv{s�|�/���b�n9���rX���1�D�
ힴ����q�w\���3'dŏ�x�-r7(sd��K?W�H�����m�/S��W��z����9�;_7vH��L{�ͅ,��do�Y�'���T�������8}vr��w_^�q�&f��#6}�;�@}��r�x�G+7�n�w�Y������;�n��`�K���T�0���;7�zlD�� z�=�=6��bl��#,�G�!YL{E�[闎�\����4}I�%".!����(~)�
�d�K�=A��K1�{MM>��Bǐ]��l����Z�@C=)-�u�v��Yq��	��(����D�L����q�ނ8��;��8WV=�%��G�%5M+���)T�ses��ߖ�A�~B=8�����n�Кi��N���A�����wp'�ZҩN�͑W�nX���O��H48[��W�DcǩRh�6r�����Z|8Cô��撇4�(�pd6��.#��W�,VL���Ь0v����٘!��A�Ό�����0BD`Cx�!���� -��b kt��g���.�a�����Ϧ�-�%<q.jeI��H�z��R+&�!qx��&{E2����i��si��ԀO��cO�b�֮�lX%^����J7GM.�!N���B�kE�҂�喵��D�~�᢫*Q�HD�|�p/�����.pQ�w���9{�k(��4�ٝ��>xv��{��?��_�.�\�N��n��>}:�~u���\���ݏח�Ǉ6����W��vu�ns���ų�~��S�{W{�˳��_y����?>~񱻯�~���v��O��v��Н�wN�_�_���#r�wޯx�w|3�_�g�9�z����7��cc-�]��$����N�t���+ǖ��ZC��Φ)�R8�Zj�	"�e���O�BY^�Y|ۈ�]�˕�H������-��j5v������`{��N����"\�Ia�\����4y�( s�q�5^
��T��Ȍm��@m�⢜~���;�sq�٢���B��bV�_�!���F�>B�U�3�ЀS3�Ne��b�G 2$�xij-We#Ts.6��[��k\�5�\!�[1^��/�!<�a
q�0���
 R�L�(Yl&6���MO�B��3��8k#�j�!�j�_HQ��M)�OȆjNy���p���'�ނɥO6ċ��\q�m;�:�ͳ��yŧ��Dy)�wi�(�������q����(�%H<Y�j������AC,AoH�<��(`�#��/�(��JR��~���'>c{�(�e\�|����{��߮W'���ݝ�_~����W�~7B��d�2����s�Օ�G��8pg��	�V��������ߟ�ݼx~t�ڷ�yd����O��O���>��/�����������cƝW��>���t|�ԏ:�<�����ꍻ����j��o�;\��<q�r���aԷK��aA��cy���ʚ�2��{[�&��Pc��-;ͤ-ײ&��`�0�Z:�K٪�5�B �a��AU�D�Gn7�5/�!P:`!�h�<�8Z�Bʆt�	;�=�I�D���,\��(d�S(��gl+7��lh.RQe!�3������X!�J��bE�!��)�i"4�/�񗽖f/�IQnȘH��t�HgV� &8E�p�,l�![��R����;�ʫת�+oF[Y CR.B�b�J�,�d�J�ǬFn�B��+eC [��Mc���R ð��Ed���
/j���R dT��TL��«h��K�a�9,V?[���)_����oh�j�YTۂ=��0D`Q�)���Bf1�������4M_lYl�۸Ł�6/WE�i6������Y�W�()�ˈ\�l74mfL
�(�t����o�%m��c�30�j��j@k�sR������8�l�Y@JĘ��+l�ǁ�l��MH!\R��!h���q��N0����Z��"|
��
��g��);����e�.c:�^=l��!�fy3 ���Z�D?����/c_���Z�t�����?���04LQ\z`"��[=�+��@˞�j���hGr)E�S��� ��K1x'2u�1�R�U���B�`�V������\(��6.�GƤ�u���`2Dũ7L�0�ꏙr� 8Z�z�,�y)��0�-�������a4�9��-�@��Y��jn�֓!��=�IP�1'n��I�]���� �#3fy���*C��8�&+]�����Gc�\\�+���AN$�a���h�*Rp�D���΂��T��(j��1d�a,p�?r�����qi�V!�(�������hB�2� ՐZ��#�������r��\8��P���F�s��$EY+��ڰ�3VV��+ؐ��Ov����+V��BDE#�!.�i�.��8�vu��յ�u�}�-R�Vү.������ȭ��D�\�\�1`�����ʎ�B>8!�6wP�N~h��+G��y�fT����D�C5�#����2=d�|}𽻼�u�v�XgT�_�K%�W�G������P�E�>�/�︺�{Is�=j�]Z}��c7����}���f�#{k7��-]u״G��=^���
$5?2����-��|з�]ܼq׽��''�"˷Zyj�������˓�7�V����S�n=��h<i�F�#���+��i���!m<�F����ظ6�t���5�K��J����Ч~=r��A���ɝB�	�y3�&��Ȓy����!��3D)��$iv��A���.V_�Cs�&;��2;E�B"�;��	*#~ų�R����7�4)�v��yu�l�"D3S'���j+X|-��!�6D�����T"�
�`�*IvLQ�# 	�r�&Yy��Y�ج��@� "��DM�8/��D��No8Mx=uRָ4g�
/�(�,���U�'��\l4 �V �t*/q >N�=�������R����E�z��w��� ���0���ѐ5�V2GaE������s�Vy��4)PV��D�ٕ�ЀsH�MJ���]sI
�I%UF�fg����8B���Y"˫B����8�,j���\�hNq�b�(q�/\�N&�MV����zQ�(�0�L޿�1IY
M^�8�8���j��9�O?����ꯜ(����7^Ծ�aߐ�Y�j�,�PWQCWA�w�K5~�	���bJ��[�j�k�-�[!xq���04=)_�Y"�m���#�/��>�˻ݍo�|��g����W_���������z���zuq����n��x�du�����������Wߟ=9���_���7>w�����������N>�l��d�s��z���7�^��	���kwx������lv}��[��k���C���׫��������q�/ś���ŵl��ֲi�M����lB����cAk�,�U���mi��CK�W�ބld��ܒ���t�Kv>�!/嚡�,��&�F�e���~R��K�,R30�h��&R1&�����L�I�2
��� ٹ�7�d�QT�
�啨��R��Y���s��"h�D���&�W������/|Jm��h1"�r��֫9N�Clb�L�Jv�)�@p��N˰���^: M6C��Z�!n%є��05���֙`.4;�p�K�>/��^6z�B|���J!�(n	WI���UF9!���,q�Z�z�p���N�� ę����J� GFӄ�CJ4m|ŗ��%iF�p��N��N�2:&88x�p�� by�h4;bP+
�N�� �{g�#mdQ�\4��ẕ,RwxD(eL��E
��+E�ςkR��Cm�������_��/~��Wo�:{�+5�<�O��ON>|zr���wO���8��������9�0�˄W>����ͮOn>FIh������gG�_����������w�OwW>���^����=��>yz��8��:��۫�w+_�::}���O._����W_��Gw��9���4�=c�,�V��kZKa�ltC�e=w0�o+[FᘽY��B���}��H�>55�j}�I
o:��vo3���gK� �P��rs�"�8�XCv!3�3M6����M$N
\�t�+Fo�	�Jа�s�P��`*rV��i�%�hM��<���44})�eā� ��\�!/[�H��x6�l�qRn�SNdd}���G��Ƿ�4��AK���V:��H����	޿W
A(')��K_"���d��Vp��	��I������0���젔�X�K���4�(R3'P�東�q	�h�;9���M���َJ29l��F| �j�_�I�,P=��hp��>�(�>NA��B�3/p��:���S^���E�NDX}�F�m5�D��Bh�u"��7�ʅ)��-HH��5��[ ���q�-b�c�0����2�_?�����%��ڸ�h��%20-[������ �Ֆl�h�#����o��D�r��Hj{H���6��Q<��#�p.v�͂=A�O�8���l��ѩ�R%%�o��\���DA(�IM��Y� �dh�W�[T�z
��d�{֣T���qA���p��ə��!�B��@�2������XƄHg�������W?���k3u��%��^C���1�&.�a��r�5jz%�Լ�R7kP[Tu�J�MPk�J�+�%>+!���o���m�7W�\�R�KT=����8��p�M�aB�^M���x��J��!����%��>��5�����"4�6g�5Ae0��1COG��N���Op�ʥ_4;�z��Ua�	VX�����y�PٓY���b��b�,�)��̪�hr��5�V����%�G.��*}��Q��p�xH%�g��k�+ȫ5#.HR��!�G�-^3�2�5���7�I��댰5�4��c�l�@��h�9��0;����f,[
�z���X�
���6\��_M��l���O��@!գ���[1t(�B5x���{/�ˌ.��^on����KƇƱ��쁚;㇍���_��@�3�旐���9�<�J�,���)���d�8�a��V���n	;\^J��w���*��/T|wx}p�浸�y��}��I�B=J�/-�����H��wC�uE���{�����|��]f�DԞ`l
���Av�z�	�����H��鏥�,_/^sL}�����z?�t�q��������w��7��*����lVG��˻��g�}sy~q�2��չ������=f�yi?�ܘ�ݎ�A��:� ��Xj/�)�V����X��d
53�}��V���O����W� ���^�g�;ce�P��=��������_��s���ص��\1�#h8wxvCsA�^ä�d5^̔�"�D�P
�4���p}R��!y%�B~��_����5�V&�(a��i4Y�okŮ64�F(8���sFpL}�^��-��[\��:_���l.G�&�DM��
�������?�&��@ 2Da�"���L�sw�%����S=��d�ːM���u�R��m�a4�1��DN��0
Zd}\h�C�j��p139�@��M�$��\)T����Y�m�)Ϋq八\lӡ ����Ξ��\�DR��m^��a@"SH°�Κ�Ț%el�1T�\4��HI͛fQ� ��zvQe,\osi�i;Ô��i茢;����������x��!���Ͱ�2��ٞ�6ٿ�ۿu��;��#�_c�/0ӖO�/������8u�Q�bf2L-N��bJ���%`��`�����w��n����0�I�=�M�ט�;<�ه�������������Ӄ����?����?�N���/_���ϟ�A�ۿ�&�z�w�|�z>z��>��+y�~��~�w��8��������+7(��읃��󓛻w�����ݛ#o��7��ݛ�����z�����r��_���g���św���c�\���[C�}���qȖ2��y��,���n�uw`�ĖCscFL�6l5�����m�XR���)����)�3�-�岙�m���/e�&ʶ���eygv���ij�W�1��RN4�h�ؘM�hXCcD�f��� �-\3/W��ε�����h��t��E��8@=��Y	PC�hf1̞޲���a����5C��+D
��M��!��e���[�@!������=����[�vK �f��?�M!-)�z�,X%��pBMo:���Y��\�A��#0j\����1Z"٢B�À��"�
)�~�@�'��MP�!A�����f�hہ���ىn'-o�\e	1L���Ew��*ָ�U�e��&�����+DFC�F�Pa!��T�aӤ��H�H� �����j�Yb�%��Ť,Jv���2r�V��CdY��q���s;�{�C������_En޺=̑��xt�s��ǖNv�	��O��r��WՇ듧�wW{���;���|�n}�z��X������g����?�x��Wo��ϓ�S�P�Ah���C7xry������o�O��~��;�������޾:�a�c�P&/��uT��l*�fz��<�`�E��c��%`1�8Vئa�����E�����^��v������o5	I��4۬tD�]�UL�@�� cV%YU�A-B����'8�%6��3dr����
��p)* �`Ӈ'UFC��đ{M�	�ʈ�͵���n-A�\zʆr�S�:\@-��*4L'M|}e3x54�F|zc�I���א�Ly�Z��&�&�*AF(�6Z�l��kh����NʹЀM�]8W6��m��`��Ԁ�c���k-�F�0�\������m'�Z��\qAR������!�̂Ƅ�"d���24
��)�T [㚫QaȕN"�hU�WjC�FGϦ�]v
��bӉ��6jZ��-c�G��g���jf�$��jȦ3e�������
ch���Ј�N��l.=/��3��)K[rr    IDATU��5S�EԒmtŊҦ�BH�!���S���/}Cxv�r��7�DL?9�f�赙Y�Q�>ХQ� 
�7�� 琗����P����b���P#��`��4]�ޝ˸]N�^��RO� �tq�T�fXΤm�x�h�&�B^}3��A�a�:S 
�z��x�e��f�P1l`��UmF�+	!�����,B �M؞&\�e.$}4�B�窇6"�e%���[�Sa����v�w"D��xv���P�ԫ����!��0���E.�Ѱp!�Z��5Ԧ~��W�A��ŘU��g�V"��Yg��8F4�e4��Pm���j��V�NASdC�j�;H�*�ؙ�)�1��-�͑?�yq	�W%�M)+3�*D@�B��ە��r�!�њ�\��ތ��0Ј���ShA�M��������lѸf.���Jb�9A�Y�̅�41�if�BF�\����M=�����.W4�,�A�zf�lI�p?�B��!fd���V�ShC@�ɅY�t�;`�A3�1
�i���t~����p~Բ�4R�nR�5䢣1����=eW�מ79�*�yL������^���Ea�]"��_E�J�ɘ4]ĳ#q���p[�%�}o��{��vs#����{<6���Oѻ��7������wv��|���5ǯ*��K�{�M����͎������+~��s�����x�&k��~O���q�[�<����؟�&����������w�c��r�j��������2Wn|;�|���d,�u_�5���Ϟ<=\н��9�}8;�;����f>=zr}q�����̓9\���\ܾy{�Ai�{u�wqu{���{���7��{i<�����SUc�;�?�=Y�6�������2�B��Vΰ�p�+�ٍW���;�`�H�oi?�lXKVO��Go(ʞdk��B��-50�
f3���s)9�B�#l#�
�/���f�sjhUΛ,�b20�*܅�]����^��s�D�A��gv'إ�H^}�i�(5��)LD.R�|����,>\�&ؐ-Px� +~4�Qj�#���-�0�jcw嵂�^��2�EU�T4N&�y���QzY$�jDd�e�D ��2j����S�Q����,�ly�B�����TS�!D/��kx�Ļ�%VF �F�N�bٲ��b6)C��JdJe$�\��B����0m}-�6����j�A�ah8B�ZR6��M�ͥ�i�#@��)d���
��2ZI�y�����[ ;C�l��b�ժ���^M~<�Bq	�_cw�c؋Z"6.Da�g�����������URC����5n�@p���!M)~��✋��Xq�gH����U��o��hJiz����N��xҳ1�B$���Yۙ���m��)�O1w��x��/����o��׎��G�ׯ�{us����?�����N��o\�Vxwu9!�2�d<r�}�}���j������ɇ���ߜ�m�n�vν�7��+�OO�W��a<��~����a|ݯyV;G�?�x�>:9~�yv~���fow<��}V{ONN�]�IYS0��9�/��:wܑԖ :~�ݢ�����)���ZL�8�i�!�;� ��h��>��2��q���m�4��I�,��mwC^��)5|6^6o��!�B�ڣв#�������L�y�.��=OeL����Ϯ�4����z�Ħ63V�vI2�E�L��>����V3,��h�*�������5{��SC���u���ǰ����ry��W/�b�����d24
v�&��n��j�XdM�U�f�zR�eN�w�������0�h!��gO&�L�"!V�
����k��S1�y� K��r�g e�yi��8��y!Ӌ��K�,	Ό�!�`�m`mA��w{Z�;�� 'E�p�[`d^4!� �E����m�����4���D\������ 7@ȿJ��>��:$6/�����hp�W�}�����vϮn־�����^����.7���J���bs�r�5T�3?:y��X�f�����*�wϙ���=8yzx���_�>9��g�;7w�w�ח;O�x���o�z�ݟn.���m�9��{���]�#��M<y鷟����||Z�]\|�9<"}x�������x�9��h�*v uh�h-��6�W��5��4V�u�\��-��(i�ْ� ����
L��ȿ�� ¹������`�d׈�߼�	De�֓��"��0�������l�Q�1��Ei�7cf,<P�0����䪷>�*���E0�V����4�E�_�zx1U�%��*6����D��k\��M*�C��g8�Y$P3�.�)R���k�)�0��)�gp̈��hy��,p�%0\�c+T��i�2-���W�̂	D�N1�5^�I�k"�1����3��m�MHY
�V�~��Ti�ֶ`r�S�VT��@���O�I�AhI�=r|�D�cj��$�OA }=D��V'�άG�m{�p�\�4q�K����z��p�թ��m�ĉ���y)�e�5L�8�.f�8i)6>�֌y�$$0|�װ,�������C���0jM|�͵���X={�-W���x	2��-D��sEېAp[C.HQ����ls�/K��g.!����p��5k���k70d+U,)���sYަ^8\��fXU��.��UҌ�)�{v5���p�j��h��(���ri�u�ԧ���B* �]א���V��7�r��g�D����p|}L=��L��ʷ�e!�N�jHm΅���|C4�ZC4vxR�g�l��L��B+�F��g�諐1[Qz�(]�>�N�	�1ʈ\
}���8l4�9d�y5G�p4.���_"���Q͉����i�$�%����z`;9?ex�4	F��hpM�f
����z�������'"��p�G� ���*�g�f5�Lr��W��މh6�v�yKm�>@'C Bu�1S���(m����8��,����.c��l^1���z /r�����*k^�3�$÷`ˈcH�׿��ϒ�n�"J�+`��A� ��zC[�笶�
��1���\yI�(��l�ps$����u��,��p4�5`�2�ݛ;ϔT�����������[~���c#����g�l�35�<�O��}�--�R��
��[��[ȯA���맚�|���>J?��/���u��/5�o�������۞�����q��egP�xފ_Z�3�������}<lV���X��F��G��ˇ���SP�Mj\p5R��T���	4YۡT�Ͳ\�[p����qS\�&���x�����'��wW�]��=(�������������t燝۳���w/��7��7���^�c�����ܺ�զ�<���l�,�{隡���uT�&[^�c�m8v�Ӷ�-�U �Yh�v!���n��~��Nq|�B������� �@C�TL{�^�!0�f$�X�Ɉ&��"��%M*��0�J���a���0r����&���`�6x5��l��W���ǽIڼ�%��z
�
�!���!�Ev����"g,e�8�A�"ÁS�>����y�2�I���]����~g:%�D�l�!ŢT0}C.M=.�0{����b�_�h�DYL�jfDH�W�����@h��ਪps�`6Gv.f|���S�85�T|逩UC?AC��>/C,��,8 .����/KRہ�;D�:lW�mD�&["}����-E�O۫+���dR�*��'�Z�ƶ�����2�)P���TG#�lS`D�b+��r.o�4� XRCL65��
@h?TF����߹����{�R�\�leƪ����_�u8�N�3qK�>�\VYQ��"򖕫=�t��a<��rL�1E)����޹��QG_y�����o���߼��o�����ã�_>���ӏ�����_|��GP��L���ӣc��q�Cog�_{��;*��إҝ�������5��{X�l��tu�M��}u�����S�?�s��z�m�͙����~u���{_�w�_�����^�-˘Ųӛ��k2�|9��T��S��i���\�b�ޙ�6y�l��XaY,�XC�2�Xa�W�e�_�҉B j�h�l.�z):��J�0Ge(	߰(����֌xف*4���],�ԓ�HuFȎ@����[P�q�=�Kd� �C����=��e&�5�A���Uh�������53�"Q��
�����H�J���λX.�O��bL�W7)���_MG���_��mU5Y|.�!��Q �+ì)KU	�14��2 zͰ�cF�$B
b���1Z�2�!I�2�4) �cC��7ĉ�NV�oXTY�!a;��R�2�DcC�QT���jn�8I�q,;[��Ƌ�\�b��Ѧ��mўcI�!pG��8��q�:�!���5�ih��m�#��(�J�t��`7�c��}՞iO�ځ���_�ve!ڒslSQl�fT#eߏY�ܭ��^]�^�_�[��]�>����վ������ջ��'��2f�ٖ��Ev������]��cV{�O�|��{���]���#��|�����������廛O��t��$��n��|��]]��=��g��3�t�˫���x;������ƃ�}b���ʗq���5U°8�Z�O��b���0�D^��j���<�"��%hh��6V�z�5��EN�V�4)^��B@�}�P+�W���&;$q6�6%���.N�٘ڬ0�>C o6;�2¥k�5�S�p�v@Q�����ƛ�t��Y����H
��!h@s�����0�!�Z�Lv[*MH�(W���J�h���L��+PvhH�,�6�4���R��$|��Ŋ���[s�4��p���`� D�!���B�[��P�
+5�$�esg�34�@-��6#;f:8-/W�B�gcH/�8�b��SpQ�Y3��!�)��G��Հ�!D�6�5��Ԭ�����0 ����*'fu����x�1*)��'["��8{WjR(�L2q|M=)#Ӂ��d��M$�!�0�˅�Q����"�����8_x�ԈH]x�Ȇl�a�E��ך���s݈�*��y��$'��VO���3;Z��`���rU{./��)ϐj+�M9M4�O��J�Ȭ6Y��t3�ڢүNA��r������q4��U�z!zAߔ�%]�F|vs1�/]!�Ct�-�+P_"ʉ��!D�e7,u�pQ��#����V@�Chk3�G�g��Ɩ4��S�\Ce��\F�[�P��J]�8e��!]e����fT��v�Ov/-5�v����@�
Ì �h�1d�;�z쟀�T����-А~ʭg��� �h��� �4�$��G�g��y��WO�-���Q��7;���Z|k�x�7�ˋ�H��D~��.4�lC
m�y� -���6�Z�#B53 �$�vid�p Nd[p�c�	��5�\yI!4S���!�H�Q�R^)��4�\(�/�%��v���B�qR��ؼ��
l�����*�H:41g1P�/i�@�@g-|&�<��j��pIj8��ʈ_=4{m��7,�)������1�pmfb��,WQ�>pA4�6�X)؉@D� �5�D��x�f�s����.W�7�7��J����9eHʦuZ�n<f�#.��=��{}6�n���\;��y\���kL��rw{�j���ٛ��OׇϏ�l���-�	���&*�s)�5��qw�.�t>�O��Z���fqt�����p�����E���WYowo���O	��▛ܚ���8
sSڽ�)����<��k��员���r��]���w��7{W=%�xw7Τ�=����������I�=�~]-u]7��ݬ�Y�ag���|��}�\�Ĳ�c?g��*����ǫJ������ � [�����o8q4S���$�����5ñ�;N�ĥ�z\����vR��Ǟ�n�������W�2�m{"��`�p��D�J�>?���"$���J&Ra3<)��ȋB`�(��-#W��MD�3TI��٦ә+�hbM�`C^:b��@5@4���6\+��BC�0f�A3��%���Ugǫ*��/f�m���ZP��1���tҁ�B�ϩ5�N�[.����G�/.}�wV�P�h����o+
�e�ҔG�8ͤ�@=�����n������Z!�����!��)�M+o|�V�����z&�1Nk���h��4^�bMl��f�[:��IBJȠ&0���!�"B_��&�-�F#.W�i.�j�� ��z. e�+[F^8�B����
���m�5����k�AXJ/i��Qc7C	�8�ٚ���!U���%Y5A&���vi���[�xxs"�
�۸_�y�����N=�޼�������ݕ۵��_��߬N>��������_�^ݾ�����p�������J�6��
ޯ�s����{!�Vg��Xɧ/�ԛ�3���Y=���?ݽ��&{���P���������w^��wO��vw���w{���ꝵ{(эn�����{M�����dm�m��m����[ծkv�@v�Y���d}�ĒRe��f��j�9��ꈋ-5f�KNG� 3H�Xd�Z.��@dL����y�l��}F�pj)�ӌC���G�>h�B�m��Ȇ��h��!�!���
A�.��=T޷26eHǐ���+5�풐k*)�X=�(!�H[�\1���F��n��I����d���8�V��Ǳ� z��&/\����/_�Ű�?����Wjx�����������@�8��LQUΨ=ċ"�ܑ��2x54���h�3S���8����*��18�a
z.�y�H:S��/�!����.Jc�s) U�D�	��PԬ�p��DcX��l)^����6=����Z�\%M�&W`�YX�vo���mh%�����P��U��^�%�u �͊`�����Q}�ÛA��*O8���/�f�\���e��ƛ���ߚ9��P��|�>~�l�9�;�[z���r��+O�N��p�Yp�y����?�z�b���O^��G)�\����[��|������w_����?}���g������pp�v���_���Rzq}���[��7���g�_>�����~���?~��7o}���"���]o�n��i�_|������bq����W��h!m��Y����V�Um�)h-�X4�Ck=5�=>�t��X�����R� ������+�jD�q�ZQ���v^���[��b#�ԑ��+BH�!C�����_��1Hm���S.�J�	�J�Ë��빐)�4N�J�dI�R�5"��6W &e�(�G�А���Tv�_�֧@���EVF٧挒K#�O�!��4�򎊗	�r�0��r�e�K��m.��r��FX8�+Z���gR8�"��f�_+�'�rÔ��#c�pS��R?��-)#Y��%c"dC�ٳ�)ל2�%
1�p3�PR��+f�*Z�7)�Y9�a)�i.z��d�k(�s���ᵐz��®�� i�qZ��/{��5^�O
(m�<�H�r^�
�vC!I�~�C}�jV��1�&�t�0�Dʈ@��_1)���� ,0r�س06Y�n8E�UOjz�m\�fT�>���+�ƕ�B�0�mM8C�*��Jlt�ޘ;��ҧ/5C��,Đ���/ e��9ĉ�h�e!;�q�RI�d�YFk�fئ��15W�\���R�D�ժXU���R�f4C
�`��B�@m�����'X��).�����hM��a����������W�>a�ΥO��\�y�=
�~�8E�G��q�O����?B!h@}8�V��� ���PP�@�P�]�!�!c�Z?'H*�͘5��/���W�5u0�ˎ�Fp�[����c�e��I�kUj}�Gl�B:�µ�z=喫!B!\�D�p2���ءX8Dm��5.�ہ����j�O�!6AP3̦L��ȅ_:�I+$M`��E���C&3�!e��̟�V���+�����Ғ�k@�\hl^6�]����wd�5|�6M    IDAT#x���س�4!%����O
l�����5`�`�p��!z�� �#��T�V�<��K/<}���*��[�8�ӟ�?{\�ѱ����[y�ʜ�����G' ��i.?�ѷl�$�ε�b����;�6?�T���W��m���Pk<sux}{������c/�#��j���#����ᾋ��8�Lh�9K���s�#���v���m�[��K�����#w]r���;�s��j|�x����'+�槣��;�;��åR�6��d9�u�نCY�����������z��c�v�������������|�w}�Z�Q��%O輻=w�v|��y_H�쇚6��-M���^��=�i�s[²���e��|�6�;VtzĐ���hv����,B�3�.g���(��v�2/�v�D�H!�$7�NQ�f=��&DO$Y�69�F�~8��M��)^�ra�bp5�#P��^z!�f��L4g�(X@5��m�f�l:Z��t���P+_,M�8���u�a��XVC^Lm$X�CMI�,&�!��*[����i��ė�p�ʠٌ\)�xL���L���_ƹ>�B(� y�*xe��@�JM!Ry���k��v�Bꉷ��f�D����E�[p^�W��eā���k���_4w���va�@hFI2�!�[��i�n���2���n��b:\-YS�Ŭ66�B�y�ٝ�5��ωl5�d}���5����5[�mtu���ag(���S%.=0����E���~�a���$oy���Ɣ����z����y�8�캦i`��E��VJ{�W���:W3L�B����v'[s0ǷZܸ��e��Z$��&P�o�xC��W��N���Q�=�yo��v���O>9<=�[_��y�r��p�o�]��3��W�^�n���G���v�x����Q���������������ݭo��cds����sx����۫��7���B�ܷ�,F��k9ӽst�ψ�{���3L�YY��a�y���Ԭ�Yn$(X�Ԭ �M8Ц��P��[g�,�m<풒%���/�cmIA��ᲰK� �U@Y�]���AU��� Q�tl�z!�S�`X^CF���0gxC�kC���� �ajB�������p�mq�F� 
�m��X��f��۔�l�D��$����d8^�z{n��3�^����Bޫ��Zo3s�oj#뒈PM�ˮ%E[�Q��&����^$Ȱߪ�1�L���Z���^s���bL����z�l.��f�+�To��\�\C1��>�,�Ф�%bT�!N����b+�G3D��>�ұEm���Έ��P�	��&����h�0L�l�"��7�b�$qHI�������-K�l���h=[I"`�� `Z.�N���͖e�)���B�Q��&� ����aur�9��Dvx;�����j4�<�M�(x�~���>�n���"�W���vN�}Z�vݏ���y��%?�������/��������Az��swu���2��X��m.7�=I��ĝh>8��ӟ�ܽ9z�������w��黯�׫�^~�5�E���8��g|�t���������?}��7�o�=�!{|z�[��O�X���x�ZLkT�U�-8��M�W��l��Yy'������m�^�mG�6Ck�EQ6���^�\��K��	լ�K�}�� �LI饋S����G���hY�3;�I�J��b�V�\J�K,�,�)��3 ��Q��v~8ļ"��W���g��p��9��\hN>2<���j
j���HbȨ͉����*oC��i�װYOM�4�EѬ�DT�=̛��YO�����Y�|M�Vgk��GT.����U�9^ͼ1�K7Ł��i{�'�߲ā؅����u��'��t8�F��
��g�"cjEM{2�����a)JMDCh`C�~/��F�U6���6��%�!nA4|��'��>B^Q�)�Q?C舒��ؔ�j�����������z��bk3�{���`X
"�a̙.�\��e�6V���&2gQB.��RTUp;��2�jl|�z���P3�a̤��z��)��o��7~C6#pN��HNM/)q+6������pn2!���Z��4����]�?.TQ�@=�����UN�M�-���װ�Rn1�� h��D0��a���N��ȕ��xk3!�-05}����B�L�ز��B��pfL'�M���a$-<��4D�9E��Pl}��b��->o4�����ν����ƙBߐ1�aF��8SD(��e���ˮxQ��z�b�p���=���#��� ^3L���5�s��&��UE��3׌��Ł��F`7��f�Bne�d�"P���S
 4l��
R�
H��PK*���h���Ȇk�!��h!oKA$o%!�Bj��^/E
�<�\����R�r��Ap�g�����j�%�`X��0���#��AC."}�zL�/|Tt>$��
�����e�;O��E�mq���8D�+J�ʨ��[�2�)j"���}��eG0�Z�� �Z���d���������i$/��"��O�9�wE�>o��;��~��y��zuyv�oIƏ;~���k~���#6������r�S��+��7�R�.�G~�ヷgU�ZjX������p�5AGoǽn7��=)�f�燒cm�C36�~	z}���l��r�/!�hk�����d�ew�S@�_�)ݽ�>>Dm.a�XH~��Cw�t�fe���o}���;�b�8�՟����:1m[{���S>��^����Bǵ�#��t���^n�0Y]_y|�Q����N�
5����K@�.,u�H���&�[��Pj��ێ#h9iƀ���".�h`6�NQ�M^�heLF"z�B����;�U�MQ����ct�sU��C4C}�Vr���\#��=��f�,�55qr1H��G����@�G "*�ӛ�	1�yEDj|�j��/E=��5��'�v�LljN�`�"�@�=$���|�Rcc�άĐN٧>��
!H���*����2l�V�RBp������Dҏ�x��9Z�Jժ��p��JњPP��t��&�N*'D��OOǔ��Q)(>��Le��d�fRC�Dؤ*2�^k�K����j��Ьes�3��&h�m�֍T}�6!�C1,���Ѐ��@�7,���bh-8/�R�L�����"1K�7�M��	^.���(by����ȉb�\oǼ�:L1lw�q��p/OQ��˿�c*�L]����/�����K�$T���ߤb2iG�ָ!�%hś!�q�݆`�������n'`��u�I^���=�����}������>�ٿ�~2ޡ�-�����\�_�lV�����_�x����ۛ�kϸ��/�]�z�<�����O֝59v\��/�<��nJ"5�e)��;����^��u��-K�S"��]3
�����΃C'���zֳVfn ������7�D�^>�{����WW�G�S��yp:���r����O.�.�ַ�����Z{U��7^aݒ�M�O��z�zͷ�^���;�Y1����u0yd�� �[�p���gY`+fS햽.��%��)�np���h
�A@����\z͚��D�h�zSo޼�zO2��R���$FxGH)�«�`�̨���S`�g�L�f��b� �!�0��@�M��N�+ZQ��s.SǂKT�?qL�-��_�P^�f�wTp�+#5=����Ԑ]�������I�����+�X
���Y;^3ġ浄mˈ�դT4�ܕ%�(���v�*ň"KFR���iA��4:��A͑� ��
�רBm[""��ek�;t�+/ZaDS�4����
C�I�͂��Z8İ��-��#K�O�!*�Y`j���#�gԤ@��b��Ѽ�q�3�e�Q�YWv3J�#5�Gh)x���S��"�V�W�h-�"K�l� �`��#�PT5�5�H� >Ns���3��6Q�\2�W����ˑ+��̢!cj�nh��R������������bu��p�z���-���|Bu���]n�����Ϟ�����߬���H�����j��]�Eك�p}��������/�`�Å�!_�\�Q������?�������������ҶO�����W�����7'g^��&�ٞ�ݯ_�|������W�q���LU�	j���[o���45I�d�VÚX����Qks�,Q[
A�AZ�����	���1-5\��\���phJ��rA:H���g��.m���e��صhM�P!�
Ȑԑ�d/����l����J�P0����P��[@xLHx�/��H��,ְ,�왫��)�1��''�D����Z��Jꩆ梪�m��ađ�N}S0D�e��4!�ȥ�֤���M�Mgz�cH.{'����l�ʘ2)����g�9
p�^y���O����>;�e�+6f�h1�>o����04`=`Q0�P���.{�(m�a�Ql���E����3
ד��K���P?r/+ɞ��(F
��o%aV�>�P��V
ұQ.Qb��[��[7��ks�
^����V�Ȇ�8�qi���5!��@�JG:Cd�f�m�,��6C�~oQ�!���!Z1���ʞ#)=�)0���-��]x��xj�ڜ#N�@4dޤ�[�%h�G�)0�%��9V	rE�:+ 3�B �JQR�͎Q�i ��!n�e�Ӥ���*�U�C�q
�A�W����D͂H� 
P1IS�2~�b+ �!�a�:!�I	I�T o��g�p���8����[�\�f��s1
iX��	l
�R�3v�3V <�4�R@+��i��J�L�C+�����J� P`y�Yv�z`ہ�6��5���!N"�%��j.W�D���(fU��gЏ\�����;������)$2�m��K
l^��2�El��C0����pV:�8p�+CHv!�"d��ǩͭ1��������ЀU�Q�⍠OaWB	�x#��ƈ��i*���Vx=� �R�\��h��P8D=e�CZ���p�F$Z�e�C�q�X��,�Wk� ��<��8���G��B��@����7�fvdH f��3/#Y����ɩ������ɋ�x�/�l��6C.|�
��(��|��.R8���6��t�Cػ+l�9�QmcJKj�j 0+�]�^��V�����[���7�.�6N�ӚJ=�U�����
ܸ,��1:�\�s����e�V�6q�8��T|�[e^b]@�W���}���<�����_��˕�������=����=��⒥̺e+]7}=�w���i��w���t�S���'oD}��W"}�r��=���z�#�E:��~N�]��G�Ų�;���3��u�up/'����˟*}�K�.5�@�X�{�?���z<yp����f�x��}q��N��G��� ��߃k���;U�}����o��?�}��ǧ�#oE77�������x��a�s��U;�|7���~����ᬑ�Z��rZG#�F;l�/��K[φ�m%~� #�KK�_�"!��_�@}�4gr
�,�q��2}��׼�I
G#�oHg�߭'2���3
�^�y!=���a_\F�n8!\�F�҄TR�zR�f��;P�'{�X!���tn���VO���z���ݥa�O����8�8\�=R�Q3���!�H����9^Q*��o�J!�C��R�F����Q�(L�bT�>$��KȖ�2��E�&����M�����e�Gfk�bi�E9�$5�A���Ԛ���Ǜ!����+�P=ڜQQMa�-B"JC�'k�^��נ�����S_��h�sU��{�d�b�T,)����а�J�8����
Rv�j�M
�v2nyp�n�����ؘ\�	:0�"�j�Y^L��ﵭy��z�f�I�ä�b֮F�~���
�X�<�����Obw9��uem�	�˪��Q�!�))E#a2���pd�XAh�ǅ`������� �by�3�k����5/dZ�T�["��oW��'>�c)������?�4���~x���~����Ojz%��~��Y?�x��|��Gs�����l뗳�n߿���셻Bl��ޝ\�_���ˣ�sr�ԙ峳����ó˳~��_�}�hN(��*+��ZS3���s�u�8�jX�D��D�[6 �p�B&�@ahM0��me8[OSR!8�!#d��r��/��lC!~^�p�cB��]�c�g?���	>f��5Q�zI�p=�^�*v$[vX�������ጚ5!R��	,c.d"�$��3]�KAdn���)8]�%���f�Uϐȕ>��B|;���BD9x�����i���s�%h
�F8�-+5H5+�-3�
�g��a�@��斎@C�ӤD��2h�
�C��-�^��6�Γ��9A�d]���=k��l�,��С<'"�d!pyq({3Q�!��aV�R�X.
��x^�!��>WvI���&����MO6�4Kd��Չ	)*C
��v��BS���)u�3E3��%JPA���p��R�&:��U-�V,2���W��nH����(�^����J���M+ܒ�㼢���q�9�oAC�������Ҫv�5�	���{�x��!�ӳg�n#��^;�]���V�Ǘg>�s耼�K��{��in2���O�Ǉ�ޫן��w�_�j�>v�����v����^8ƫ�c�����}�^���g/^��NJ)����~Idk�������������ͽ7C��o�|����F`�O�~<�ʹeaX({��[p�9�w��ű���S�%��[4�U�Ѐ�L0�^ B)�"��-���O����0ô���K+p�`�6/;Mᳶ���5|Y;N0�!��	��1{.!��"�CZ���|�r|`�r!��Bf�y��&��c�3x5QZ���v3DY�z�C����R�"<����+ q0�ΰ��@;�s	�W��W� �5�Nʐ�Qa4�p4�JJmj&��#��>��q�si��8�h8�"����H�.*;���R�w��� �|��W�,��͐�4̓]?j�iz|QZ�K���4�B��B���#��~lh^ r:l�����,@�և�����jӋ�f�X:�#l�c���nF`
��5�8p5xn�u���L��&�N�@�)�����p�q�����ո0�@Cv�2����-�	���&�N�z:�f'^8�����T -Y=��B�#C*�&D��E�7Ծg�%���p ��L��'Z�8�lR�"k��`�SU�2���(A��>e�V�N�?�#���kSЪ'o|�(p�u��>�ttx+)�FD�R�OW�~�'�j`��x+V=ld���dCj�֫'ڬ�B��^d'� ��uY�)K��R�b$����ʓm��&29bK�~�E�1dkM2,.���(��@3���[��XlK�S_���%E��J��XZ��#q}��-�ؐw9���0�Ũ$Q�M��yA�U�.�j!�j��6|C-MI[��?C ��;\��x[1�Z��y��>��rU�����͞�̒s����ːB����-{f�R�@H�D�!�!��3j杹�U��B4�o46���\�^k� �+�L�1�p�j4��r��Jdd�7�Q)㋭��B����Sk��P���3#������a8��M�n��M%5QUR�%
�����!���x���.!�WLǆ@
��(ei�1(�;'&�j#%�8/2��oXm��Q�ë�j���J�p�w^f��^ä"d�|h5>�ڡ�n�|�ܷ���4��R�;�n�*����/����zts,�w�~Z�p�vomӽ�?��'��f��󫜾A鄐�s�*u1�%Os�<�{��6���|n����3Ǒ�w�:�31n��䮹k7�u��UHo;��i�\?Z�Ó���θ#�	8Z�;��?��<��0 *�`�Y�	��mK8�{�l�Q�-������������볋cw��[�/�mO/�^<g�no��nVg���)��͚��P���X:�ut���9;?���G� �_*sE� ��Y��
�l�R���A�v����P|{:m�eqr�V~|,#.�}x~`8�������C�    IDAT����)D_v�^������ ZYD��&ؒ�.�P��Xx�Y7�c�&�m�0��"�!�e�"b=��tH5MgP4S��u^OH� �ܭ#�
��ٌ�YR���Ә?��O�,��d�p,~u���p!M��U��������L�W�:�';�)�ͥ�0;�����;'�e'��E�2T�L_1z��� �xKiAЬ*�)i"���W3P�����Ș���Ҁ5KmY�N�;Y�8G[��x��'e�C-������L9&#{�<m�%z��Ǆ�Oo.x4���l����m1%R�T�\.kC\Z��sAF�DlC,C�b����%�Ũ��qS�AH�W f�l�X�rC}^ �� �ƅ_=z����*��,���N[+_�������I�xA���C>�shj�"�;|�j�+Z6-F+H��V�y�����K���L�M_xt1��Ŏ[��?�)2˱<��n�~<9�9���<���������]�Y?�|y��'�{?������|����f����G/�����q�������{������y���n�G@�˽�8O�5��g��oo�׻�����<<|�=�sq�(e{m���-2^Mͮ��s�wa-���f���ⴋ.�x�v@S@��P���t u���B��=��plM"8CIC���h%���������@���)��a3��>�sN��U�����"�5� �;�Q���4�v��+#��P�v}jEM>#���a��^�h�h%U�U.S�Z�����|��GD�=$54�De ��� ���zC }e�=�T�1��V�L��(��T�1n�?��/��B:WUK$J�jF#����*LF�a��j����U
��I=��=۰��i�!��I�!�~I��p� �0q3�(D�@�� d[18d5�yk�B^x)����P�@bR���[L�b��f�5�/0~���O~d��8�B��\x�R��鏹V�6��i�(hpK���O1�4\��2�'�+���]�WC"-���@ނ��pܾ3���w�Z���PE/˫�e�Ƴ�#Q��Ŏ�Hw7߽y8:~�G��{�l.N��V��򻿽���>���?������o���?�e}w��Iqo�h���w���1�����St}�fu�����}��������'�^>�*��?�����VGO�/���_.�R>�ytyy������G>��n���������W���Ͽ��O����&^Oܴv\'v��6��*���2Y�����&Doa�U�vL��>D�8���w��.�^���d����Ed����v����!;���/��N�T�4�孆
��YR,f�ݾ쐥���Da*��\�puJ^�\���b�S�s�s�&
^��z�>g"h��y����=$��U$N��5j@�����>`v�1Ii���Bo"�K���H��WGljɲEif����;W{��u���@.cR��a�s����y�Mg�b�	N��z�x���*��O��Al�1����2�K�D 5̔!��-2>�t�UO�l�Gꑋ�S�Rc �
Ѹ
j#~i��C���0�%�0Y8�j��w�_r��6�J�'�S�����O�tZχR(�^ &[����sѧ&��z�"#�C��8zC�hq���
	�U��	"#~y�iN���%Ma���T[c�x�t�&�k׋��Ec�Z�d{�)HA�筏V����Z���d˥�+O�0�l^=\�����@Y�\�
u2��JGxC}R�R��(e�P����t��c2 r�����%���:�g�4gU@�	
L�J��"�{�\�W���v�[+;�K�3�Jjq2����q�;�!l��R�!#�	�,�L���5d-C�&vꈅ���VI�E���~
S��\p!8U��b��>Y��@+۞�i�5�Ld�V�I�Tme ��!#~	����$B A@��a��7G��X"�������/�!0��@=<�!/�Dz6������U��PT%baǏ0S�kS6)^CF�M*����Hm�$������KH?<�f���v��g1�գ��%bL��pʻ �K\��b!\��ΐ�D+�t)�L�"����j��ir���[".H�)ԧ�&�� =���K$�t����>��֤�ja��-�X`��5��������;��w1D�O��+/���cM�/o^�:\!od�k��jHM�zᲗ���݌b�j�o�\T�k��J"� �g慣���Z=�\N�y�ϫ`�@	\tt��/�q��F��=���]�\@�K��EGo�}�s,�؀AQn�z�������d<.2:m��.w�� }'�぀���4�b����'�Ի��ps��*%�M��V�{n�亠���h�ڍ�+����噻�/���U'�GBmX.�v`[%C�cZ��p;�ҏY��n���ǟs��k�{��k�8�/.���k�g���^�z�����G�w�g'����{~m�����6+_����q�ڪ����׹kʵ�ʰ���n+pl��ϴr��@|C���A4Sӓգ�hlk�7}c>�l�����8w�LSyR8�3/N6objh��p)� K��_�3������i�ɲ5v|d�,�jS�D4�	�l������-�p�tz����D��1p�Tcq���GӸ�'��`/Vsˋ���B�P��"�t�JdH����7�Wm,
H�\�O��2��+[F=r��j�ed����N C�Jz���t���Ddv�*��4`%�X�z�!P�Hk���dG�"��d�=�@Z.�Ef��`�����JS_��'�@!�@C���,�8���Oְfؤ�)��*�Υ��H�*����B��ZϦiU�qM�(H��Pв�mYy���N�[m�"T0�� �O$��"�!�)Uab���b��Wc�E�G���P��C��o�ƥQ�[���+3N����.u�v��.U/����rk%AV_�5l��9����^0������8���ڋ�X���<�B�cE�W�{��<�?}���������`��x�G������o�O�O?�<~�Y;Q�o�����^��ݵ���/>�?xwr���|}w�5�����?<�z�]������:x�Acme�vh<�Gi�e��4Ǭ!��U;i},���P֓WH�E�x�çƛ����g��%�HJ��	QR"��1D�L�]Ʃ)d�ey��MJ��}�ķ��������u{������	�DeT�!�l�)�r*)C�8�d�p�6���Z�f��&c��5x���4!�BM����H�_Qj�W����\VI���v�D����R�~,ʫ,[嘡/Pk�<8�b�����Da
�B���d���9�)$B�� �c��pe�����c�����t3)5�!�㇬OR�e�կf'Ra�y�q�����0p@�'�2���� �!�*lep��5���|�ëD��41�]M�r�e��Kƅ8�"�$L��>:�Qǒ�ݰ�Bd)0e��g��Gk����Q�\�O#� @�-��mU���ի?5 ��F��tZ4"x"Eٸ��$%
�1P/6W/EȤ:�)���zz�+�75
Rck+���ϟ-׏����i�����{���1�����^��~��>}�7_?��
����qk���7g����_;VWoo�Vw>��w�ڷ�Ww�6<��J�5ܞ��^�88�{t[���7��~u��WO�>�{ώN}����)�p�Y_�;�>����x��흗#/z�t�=�����;W�D3�Y�dk=Û/9>[����`�Ze�)pQh[}Hӛa$����v���2�Xj��h4�|�M�b��g����c�RK_T^|�AA�����!2��Ɉ_m��)����(!>��P"�������q�-u��vɘZ!hqqr�� R����H�^�����[��.�pFlUw��[Ҋ� �B�[v�V^`I�2��E�9��
I͚�@F�!-���!L^��d�%�m����0$C/$��I��*�@Qy+���*ԗ�:�M�a�b#0:��D��@��2ZC�f�g?i�?é	�S�ͽ�c�B�-<[O<v�6iLG�A:l t��c9���_����l(�&C�����4S3S^C�i3�r��K�q��	1,�1�-����B��Xh�+E��Zd><��Ł`���J��j�\UH)��)�@C���:�x��S��F�l� /��f]ld�r;@|��g@TR1�MVa�s��!��pM���)oI�4�3�8@�m͌b���e�����j�Z(�S1L"�)��Q���f
,]}���R���a�1#5i��e����U2�3Z6A�8�W!$0�,%-�UB` C��PaiB
�=r��Mzx��zz4���Q��>�@4�i ����eT��eѷ��HJ,���&�R�S�nH��gK��5:�!34�~2 �X
�b��I�ݺ	O�s`K����raV*�&;W)�UѪ0ZI��Ѵjc@p��.�~��qB
4��S�f�^�*����.`�ٲ�� c��0���[%��4�e�WI>�%RI���D�]o(j�`@J��b�L�+PoH���!W��*߰�������e��1����GP��G�VXT��>MRm@4H^}����i(*�^3�x5C��0�������m�zd
ΓiB�է#ќ,o�+�'�����ǔ����
,����fT���(j���ow�8%�a#0�Q��/�ls�[�z"�j&X�t��5q��}W�T��ɩ�.\�})���ƸviI�6������*��b�Ȯ_���%K��RF��-g���w<��5ݞ�ܐֵ��S�N:<;8z8�O�2v�5O�zr�I��h�o[ZI7Cr��7)��{�{�//N�Ƴ���x�-��k_�<{>\W%�t��5��ß��:�d�sI���(ݽV�c�|�x���x�[��z�G��ا�>�|y��~�6}cӎ�{��ĺ7����έㆈ>�:_�[�nha�������;뚑��"��\�j��e/�K�6����&�c��).�Q���b�I�����k���8J�)5й��T���D*�>>{�dg�@����
1^ϥMC��@g<p�56�b^b�=@pe�G�eԚu!&Ճ9e��n�g�!~j�5:���M�ݎ�T���$�)�&;�؁�އOA���z��B32YQf*�c�`��F�{��� k��y�P����Z!����,\򒂋R�thy��+��	�A�*c�Y�W�����_|�ɟ��Z���!2VC^��~4x��#�!N60�������\���!=�8d���� ��z�V�"����2��~"z����!)оTg^' ��T��P�H�Q��	�U�@D�b��B���z8�>�M�א�PcDF��S���s�B��y���p w$x�����ޚ��;]kqN�IOrI�����D���
�R�MTS��3���r�|(�;�<�x��x��AЛ��u��=���t��'v��桟q�������~��O^�?;w��;t�Q����Ǿ������_|���,���z|�}z�<=\o7�n}����A֏��G>��]��ٻ�_=�<>�Y��#+��t�t�ۍwn��N^�����:�b�߂,�{i�L�е�h�4�i}�y��ą�-�=�V���l)��[�6��@9~j 8َ��Ȑ"P�B�J�s�K�=k(��6�_~���b�#K�*�
����
c8��@���+�`��^8�2���0��?���7������APY=��ַ�@.Yx٭$�F���[:0�s��)X!�����4my]x3��&�&���+v
z��_�ޟ =�)�w�@A����y�5�^�U1l��
�3���M�t��i���GSF�۟R㘈�S"��I֐�����k�bk"*�t)K�t4��*�z��@�J����2l�t4I!����5C�8ȶR�N���(�%��k�p=M�\�2��\!�j`��U >���k*@
O9N!��^ӡ�U���2��5�)t�lM:6�*��+�j����jF��S������D
�(��Ls���h�i"괉l�h�G`�V����򓟨S�}�K%�i��������>���rs{���n��v:��d����[/��A�է���Q���W߾��O��{??����������9>=Y?<n�?y�ɏ�7__������b�>�_���7o�����ڻ�9;~{xv�ʯy>7��G�9�QT���8:p���ʕV���vs�=����Mw]w8�����Z���dM�CƳ�E3M9�$��[����p�����ϥ��la�h
��G� W�\%������&b�b2�$�a=�X���`gP(��DΖ�z�w]�+	3�!��&�!�tD�Wy�fI!l^-}=���d�+��z�3\�ē�0��
4l�d�H{���K����;6��p��VF�d=$�
0�^���c��O$A~.!�� �!�zpQ.��04���/��������/��j��L��k�qY7��,�Q|/2��s�0�E%>{�\�c��H�S��בfؖA4L^��B�ywW�k�rC�o�J'0��6�bC(h����(��\��7Sve�i>>v*x"�֭CŐ2�&�|{f�'˥��RpMM�R`�!��I��_���+C/�K��S�̕>&�p"��oX��h�z.���J ��g����i��M9�hDf!S$c�hs������T�I��\L�a������a۬8e�U�k.�Ô1�����h�X��
ѐS@f��H� PHÙ�r^.��H����4�ƈ3+�T��V�J�EI7�s�>�j��w ���w7�0&B�z8�V q�Lo���'�{M\/#�P�&�Y��T{�_ü��IG�a���'��K4��!)�3qF�����ъ�8VU�B��2�2�����1)3�,QU�eȥ�T������BC|�3]5��^�����g�Dv�o�'�]����)�[F:����«�S� ������P��H��S�-;�D�����x�E����WY��8�
˰�)�EO!BGa��P�D�-�,�A�@.|��MM����0�<��!P�-����y
�EO�@6/�g���QF=��k���p֐�~��n%�y�Bd�
�A�M��@�\X.�@��,�@ e6)"s��!��ፌ�	��]-�QxQz�C����Q�Ҩ��0&���xce��ws�K�Gh���ȅ�,�Ɇ�/��Z|��CM �@� -�os���Úp�&m�]��ݸZ9�%s������]֤8��-�#jd��(&���������&�����p���Cb~|�f��^:��L���ѳqg<�+�5:�߻s��ѳ��ܿ;�UΣ�������_��/�����97��g���K�
33�+��g]�d�#m�T��v,�]y|<�8|X?���V�7s��{mo�G�oo7��ͧ��7n�7�w������#��6g��"�����~{}�w��s�ky�:t
����y�^�ks<���Rt�2ԩ�Jr�y����&Fn��|�G_j��c/���h-��05!����e:zEu9��#���';��J}�{{V2�
�5]��P�*Q��_�@j	�sMf��ژ��Ny��B�l4�[^s�Kj.x0����hB��L�eAhXyB0���M�1�lo�4�vF��R𪓦ʉ�U$B"8�v
"��p�@�sez�}ϛTʪ2D�B�м�:�f弳 M���ɔW��,>�
���ԔZv����] �>�8��b( �_� ��K.�\�(�����-C��4e6�~�D�me�K�@f%Dc�2r�-Α.N5�83d�ᔂ�	�z�l"�u�=�FM�8���B��e,��8�l��9�ێ^"�;�Q���S�VK��6U��:z�� �Iw|t��a^I�P��	���&\�S���!�������գQ�|��75����͗4<���@����r�k�H�S��`H�O>BҨ����qZA8Q�@Ṳᵍ�@    IDATUi��-�#�ԃ0>[4>u�qH�v'G�ӃӋ�����խ˔��tps���`s|t}��=���7����~�n��^����"��ˋ��¸��ߨv.۝����؞��/���g�S�T���t�wx��]{�?�=�Y��S_~���n���q+�8��6�y)��c���f���⛰V�m���lL���C`]���׬R�lq��8��s����P�^.�?��¥�d��Nٻ��(e�\C�+�����#VS9&�˫gS7��!�����B�"g�� Ѹ4�ɠ�n����`���\��Ë?�LhY��"-[`�eas�L��M���)/A��@��������10�jϚ�=��~j�ۤI��d�/R��A�VR�J��,�9*�)0����'� ��ܵF�m5�SP�_|a�8!���F
�'����ʥM"��XG��( -E�(�P���¼\%5������H��$����Q"�l�6A��+;��
&�+�FJT}:�@M\#�48�h@Q�l���؎�Y�����Z�µB���*��2�Bv�ٛQ��w�eI��«����HAF�%;B��5��E���J0�8t�r9n��]�t �l�ݤ`�e��z:
j(đ��KO�I��I%"��V�P����L�4��3���g����<�}��2��M���c���{���۫w����'Gϼ��"�Ǜ��fuoz>C�tt�v�wj5ܨ����������w�w�wbǧ�9�w�oN��n��ݮ����?��ű��oT�'H�'G������k?���������ߨ��#2{��S�ۣՑ��1������\d����.0,�Y���n�52&BK���ᅳ��e���4����R��m��6b�Bd�\b�#JD_����"�()32��f����\�'�]�� �5a��h5�V8�K����f��A���auf�$%p�`h!���!=�Z�
S3�*a��)6�����̙�t��UU��)��54F%�j�OY�f�o��J�g��p��eHM:v}F��9�a��Kk�4SKy�0��u�o��S��t،�'� �U��+�>ex��R��K���1�e��_8Y|xR1��������y��$rȜE�����T�e%�F��i3R�RM8�rՐ5�8�b:�w�b"��dT-�l-W}�L��H��h56��W��Dp ����z�l�jF��<F��x �s/�vjs�0Ѫ�A�]y����d�x`�l5{|�)��$�N�+�t���`�|���b	j�B��=��J���ë-D�,��mA���@S���j��*g�4&�YI�R赪ep	�.2�+\����5H����ũ6� �A��~`Cś���K-��Iڰ !�@�D�%�8А�D���)V�T��rI'��}|��h��S&���w�K/�j/��0( [�B��"0BI��h\�a"�S��aE�"�#6W
)#��ͨ�"���D��wJ�BO�,�yf�$:e�w���� J3��lH�ʨ�l5D0��Ȑb6����KPC(
'M��6�Mg��B���cV�d2 )ף��*��Ε=e�w����w���!TrIK��-2D�xk%|�|,���MDH}�b�bp���s�@�Zv4Q�l�S3YމL�e7,W
��s]o7�ů�����w�T	>Ψ�8Da:�45CM:���R �n^H�J�^H�45v#~)�S�p��B]Ų�*(
(i"�sRg�)X
}�>�+�P�r�r|�pʃy���y��;N�~Xj�.�Tk:cb�eBo�������DQ#����ɾ�Q
_Xt-�;Eg����+c�|9ҧ�W~����Zx'���,:ޮ��t�qsvq���Z�˰7�6o��|��T��gkbB�����X����fĵ���Y{]?8'�G���9q;&�j�N����?�}���7��[;�|�^�nO�{������������������ͻ����i�r��N�^��|���k7�=�z�=����q��#fNC���[���K��6ێh��x�]�A8zޞ����6�&&R�j�{Pp��S�"P���ڗ
J�v��)J�Yd���EeK�&2�]�l��J�l%�	dhB�),��'�� ��0��:�D�����R'\%&�\��K���o��h=�4�MG��](0�PY�)T��Łw��WF���D��v��I��������JJAI����1�W�(���i�+
�8�,��Q	N\OY".5hs�YR�����l^����	[��&D�xRpM�\�K�U=��X�c"���1Dy=y*C�p��b��h2B�����!��ِK���gϐ����l)l���x+�F0��Z}���ά��P"�eI�tȚ�;~��wvN��Ԁ��;co���2�4�V�@�� �~C8e�PsQ���Q��{!6/�qI䢘��,�Բ3Ȋb�e�H��P\�-��kW
�|aL1
C#��x��U���|뱅�5��y!ȹT 7��^oȶܖey���6������=��7�=��|��=����~�̋�O����'?|�٧g�/|��d����3�OO�/�ܷM}���%����9�٥�o�{�^�^����������������������]�Ni߬�6���p��u��_�n]�rnw���$�i���-�|-�kW��B��~&e�������Bzr���[
L5���g.:��K���l��9�d!Z��H�v�C�tJ��:R�����z�T�_�"�'%E��ήͫ ���J�t�f h)4����K�S���1ALv���'Y��\sȀ�5��
��ׂ͔p��G�YL��܂��!5N`��ҷ���_��3��'���M�.+Xv��,�����g������x-2�R�XB �)cK���L�s�B .��c	M���hz�G����"Um���������o�[����;��R��)�24t�>Y�h\M��i�NfY\b'�b�-#A%��fT�\&�fLe�0���d!������q�j� N�@C%�N2���Ed6c*TC.�e	��Sϛ���b� �05�p�6,/����fkt�BC��k�vVH�z6���;��D8����ґ����g?����#R.d�^R�&U�WS��Ж�ٚ78� �__<�ؿ;Z{;�I�7�}�t�ȡ|䃕�7�߭W�o������ѳ��ǻk�>�ݸ��zs�s�~Y�p�>���>l�N/N_������߸E�����w��믎N�}j������ϟ?;:x�z����߿�~vyy�������������fux�w�?���������j;���XU~xF�D�o��	��{�y �*�!�HvT�∵�ʐ�°�D���,�(��(�Al�ZF{���XϏ@�k�4��e�c��b=�#��D�g ��:�a���414;�K:]!��!�\���dL�������W�aD��gDȦwH��)�;�'����2O�S���q1pJ�t�D���E�A�l�<�bǄ0��LQ�]j�S|Ғj8eӬZ}Q��s��i���ʈ����F#�� ��dk���8?tq�#h��n�ҏ��A����=�Ӂ00��D��w&b@,Bj�mAxd"�YZ�ʨZ�(.���5��2�jɶ��v��,l!8��ΕT��p��.�e�pi:1!�
�l��نs�r`j�� ��,d��,g��4���!����k�*A�^vk��-��H��Hi
\Z!�!ā���R&�gC�>{�F��§�:�HƬJ�e�U��k6.W�R+�pf�c�G��U���~���2�0���S&X�I'��h�0�5Q[Ip�R`��"�8�����)�]���6Zx}�i�}�K�a�T1�UdU�B�sM��w3"�S_^�
���[Fê-v�b�S�CF%�.��!%n:�i�F����P���صRD�d�\l�c�U�fkR^^C��T�쳒��C�埼B����V��E#>5���!Z�Je�xRgF���P/��n"d��Y����۬���tU�~��)$��(�� ��V��UjdC�!f!�}�^Ң�7WS�L&�V
 ¬n��I�_��Z=����T�>r^���1]��mʬ_,\�����!�i�2*&$��G'X�D��Gc���i����~&e��M-r��D
i���\��yَ|!l������۹����fsVb�Dl��A�1$�j�<xC\1��D=b���ʥ
�O�K���&��
�8z�2���j�'����Ws}�*w)�y��q�q|n��HY���go8�w5��<5��,h=ϒ�d����_.���X�O����C��_�]����U�˃�q5�4�DN 8�u|t�0�n�����#g���WO75�?}��7H��>��˕Ӿ�ߙ�;�m�7^�R����;�˺y�5n�7n�7�@y�}3C��2�|Lmܐv���xA�s5�߾�n\����3̫�������t�%?�������o���6��$ī���>��|y��/̸������i{yx9n�k�����⢌���U"�v��Q����������Kы�S�x����C�Xͺy�v����xg�)�����t B$*Wes)�>�,%b����
,/d��r�_��D&A��U�L�y�a�D���e����i֓��,�|�O��<�8��Qւ�Q�kG �jl�ф����gip4&��@��9���n��N�R��*c�b�$P�g ��J�S.�Al4�'�D���<'Y�a���(3����|ٲp	��Lن���칺����K�aj�,�z:y��
)�=u�	��� ;�S@�	d��g8[�j�j� �fXC�Eҙ�8hIA�'ȰA��ģ�l�h�J\8�;���BJĴ��v�v�Gǉ��v*�(��ν�}4����15� ��N=U"�\�Y>:@A�=RA/IR����;�a�f��"�aR�	[="b���zt��65!.���hJdR����i�\�Cg9]?�(R1	�T$K�I�i�ϔ��8�bơ0�C�I�[�hKo��ژ��˗!�.J��ѝ7�]a܌�Y�}s}r��z�������ٗ��싿�����������7ߺNg�O/~�ُ���<��F�������k�������q��OY�J�ow>��F�Ëן���z}zw�<>��#���޼�^�b���);�r��]oF���b��a1]46�J��VƖ;�:�EP0�~�왷n/R�m��k��@sT�O�46M�&
GF��������������oQ�����+J"MFM��Np�2���)>XT�J�i�SL2�ig'��N"&X
}�2���o�a h��ڴ�N��d�q�t��\��q�b^�F+�����+l5���#ӣρ����/]�c�}Y�����ʨ<���gkp�	!��7l�T"Jx+��˥����N�_u�G�NY�Ɣ��WV�d;n�t�Y��Ө��J�􇸫�Ѥf{b���fF���] su�*�5^�HI-E�YF:@�vͰI�PIB��Z��)L!z4�e�a46#$�^&E��&�ސK+0��YpQk���N!C/v�M��51d;HʎFP���P��d�,d.C $q[f;�D�YIM8\rOw8]6�Ԧ#@x��zTE�W���O�9N�h�N��h�sU���pis���zW5~��}��M�w/�O>�關���� ���������׽9:}��O��f�=������ũ[�����ӣ��S���Ʒ��ܖ�����ǃgk�7X�=�Z���no7~LӇ��}�[�/���=}w������<?r�Uu�����շ�����2�ڻ�~뱻^������+_']��Za+�4����[^�[���k�a�o�0[̼�������d#H�Yyj�S�%�[`�"��k!�b�m����� z�H��a6���6�5��L<�P%�J��M�=Ɇ	NĐH��
��+à�M��y�"��Ţ�e	�Ulx|dC������X`���њ/���8�Z�GB.�/V�b
�A�2�a�E��5Edi.���������y�h�d��hڜ�b2�&9���f�E6�!�ޞfO�iL��xQ�o^	�{����%�D=�"�,�2�Ӑ����
lr�Cx��i��C46D�v��9ֶz�J��>��
�� 2�J�7Y^K���q5��F��҉Y��،�^R�tDE V��p� �3�!0q=�+�#��)�k3�Qͅ|���*)Q���qT+�.�0e���#c&l���G6$>����Ɉl����50��-��VLEgT\�yKWxj����,�?�Z8o��7����5��B��T��o1L��Y~8��M�Jx5!pvS0�؉�&�w,�c�Xx��##̐r!L#�!���3�U��b�ÌS�t,���"V_���p���,R)��4[44MH�SH��(F:��X���~JULR���f7�	�Ԇ�!>-C:!l�K��0��R.̼p�!�el�!�Tɔe@��q��:����Ԋ�O�DI%R1)Ԇ�Ǖd˨~!4e���7\B�a�aԚ�L�F� �:!)ScWL`�l�,! l�����.��[�-�J�5d.�3�0 ��X.Q�Ų���h"h"�K�N�q)�^kȘ�e�� ���_�2d�獠WC�^3��
1!���J�)ݮ7��%2+L-/��&��C�L����)���3��J0��2f��ӌ���1��S,NYʮW���X|x=�d���T eQ����/��*�k&eWA�XdR�T?'i�Ƨx?�e�����f{2�v������\�Gl}	���B�8;~��w*�:p����b���N��f���:��j�;m�1n�d��=iѷkW��i�m�վ����]����bup�����K�������������S?��\:\=wG>��u���}�s�����������X�l���h�N>��߳\�;~��ک�����]���O�<=�[��řq�t�b����M6s��p����5���r�?���^��=�,�_��%�'�[���O����q|qs����c�B�w�����)z�3�zۭ���WC!�$��+�aߗS�ljzA!;,�'�C�(4C����%.K��i�Q@���<�>6 d�26)�=^*=Z�dh��Ȇ��?�T�p��Ĕ��/�f������aǇ7�/JH��ꔈS��F&�0`ӡХ��%65�Д�3A|�U���ԀbU���҈��U0��;ȅHJ��?�z0e�`�-[�^F��-��� h���k�\�W��"�Z!�J���~�B�G���N`��4�(�: ��ӟ��Y,D"��F���gG`��v�83VR�\8y�����4�*X��e�@�VF��5�  [UQZUQ�[F ��M_y�pdq�IWK�/�"�,��uQ@�j��PN���G����l^g��Kq4J��/�y~��$D�q�c�T.�@�:A͆�r���1��d�ӡp����u-7����RR��?��������TDjD�'=u�h�6�6�f"^O�Q+%NG�Rfeo]E���b�8�;�#.8�5G��ø�Ԟl� ���<9�w�?�*�g���_~�������{���j�������ߧ����/����G��\"u?�ǭW���?<;��{w��܍V~7���O�=���y�>;v���K�������h�����M廨i�ͯ�1G35/��z�'A��E����	��V�3�G�e�2��7�!��n�)S��鴤Bj\�\�٤���,�*T��գTe��t:��u�ķ�
�9vji%�R@zC��%�r`5��sE�����i���r1��E��\lx���`�j�]A�Bpf#.�ئ/\��,�Ї���?�®�&��l�,l���W��A�@���A��n=V��.�C�w�dth����C¥�"u��4�MCA n�6�h
�w��R�3��yqŧ��x���bUj��/��pM\�}o�Ӝ��P�g+R��7    IDAT���izft@Ҥ��T�(y=��r����)�j��	��l�����	��Ei�I�4E�a`�n2��\=�5+����
�Q����:�2R�d
Z����%W������ڔ��>^���\8�2�t���V�9�p
ʳh�:�ʶ�@+�+���>��sj�(4ǰG����c^�ʥ���N���*�b��?l�isd�u�{ U���9���cK�,yv����a�_x�k�<ȦD��E�lv7�
���t�u����zֳV�
�w�*C^I�;	��9~���/f��O���]�|<}qp�9����p���g��_n��o|u��ᵏ��zN�|}�~o�����G����ON� \ow'�'�^����z�r���7���_���w|b�����jwz{py}�p������������>~y�<R�x��|�����W�������������'X��s[�@	>K�#7�N^&���Q̑�Nn�8o[Lk�Z4^�"X
�j�1��V\Ӷ�^;d(
��m�%��J:׼�� ^^.�'bX�"^mp!�v̲�ͷlDR�D�Z�@6�ROB�@�)����-�p:��	V�~�ņ#�ǐ���KWyl4xujµ���"��a�
��7,V�%��Cp���'!�Vc�[��ɧƶ3(F��ҥo�� �Z��o�
����������͈M>8}�ri�P�Ũ5)Qp�+&[�à<m���g���\+j�~PFPC=��q ��7[��V��ؐ�2��℘�6�(��鰫V�+;�@���������NxL�24L4��B:%*STQm����D������ڂ8^s�<+�+(KUۦq��Ӑ�f��5�E��0.�1�Ry{8WIc�zд�p!�@^:i1�?)d\U3����������r��ʌY#o� ���I���.��F�f:z-(D�����e�U�DS/#ZL�PÙ{$~{�3 ��|
d����UC��!�t8l�r���R���Dz�\z.!�ay�B��AG�~��$���7,u!��<b��� Z����é5̫�S�F�"�)�G"T��E-�< �@�2>p�36�@ä2�HRv8�-G Q3��BC-;)CF�@�&W��.U�U��&�D��l�13�i�^fes�!�Z��b�\Z�ad�>�d�-����j��ȥ�d�;��ˮ��˨o�1�ֲ�����-��lNvs_�Ǟ�:'X����H͌�q�}c�����&5Ҍ
��
A �����^Hń�3j�8�d�Ǝ�\�y۷+�WmN�f6B!!�<��Ld�Ťf�?2�aI,���D�]�����ț"D+V_�Y��fC4L
��)�(�DKǕrR)d���aB_�rEhDK�!�JW�fI\UX�gK�LDc����+���Qn(6�D५�+I,Z� 6\ߎOs&����zU�%�ͪ���V��hY7S�p���� ?�56)#���
�]�-<R�惫�G���C�Ia���ԣ&����w�N�(Ͻα۸/����u��km��D��?k9��g�򧎇C��~��Î�ɡ�[�6�~��#�=ҵo�󳔷���WW�n �O��޳���o9���{�����˪��|�oy�?�O.[���颭k���ಥ}�����Rl�F���>��w�j|������>ٳ��^�N�̺�>�ߗ�����=یo�}q�r�@s���~w�w�nn6��GW֫S����ݸ�9����ѧ�e�Њl�i�C۸m����f��D�&�׼�W��o+k4K����%�LG����B%ʞ4`x}!zySX�ǎ��ПH�4��"���\���z�ͼsȘ|^�z��e��e�����J��!�*�2BL�"D6T�+W���=�[�B�Hi]�U9�>A"�^���@uJM�ތJ���!���[dsqq���Q�*�R�x�ū�����I��%6Ќh���WgE��*Z�T�@�«�2�˳l"l5��#А�X:l
j�"Ce`�E�R�M)D��(��=\K�� G@���P%b�E��׋�Go�>�bX��U����c����6�'\�/Ŷ�S�M
��h�(�ZU?�&Į"����~�ͅ�UUb� �Km68��24|}�z;�'�|��>�+󼲸3b^��L��z�X2�fC&���^�����W�:Eّ~��y2�~��ԽK�v[��P���m��j%S�\8))���VVkJ�P�"��D6�p��͖CC+�W7/QnV�W�������~��������,݇<<~v{�q�?�v�5�Юp�.�vܒ|���[V7��o������������L�Ӂ'�ww�����V�q7կp��}��k_v@�ŷ<��Ds�:����g5}���vy��=�������f�`��?�#�6�;4fj���޲�M߶q_Go���w��������Q���su�Q(l�1�5�B���7ɼhE����+Ўb��H�"�4� ͹�yS�J��BIc�ύ�+#��!��\�h�����C�}B�R��񵆊�!8�JP��h8r1De�d
3���mWoh��tf>�����g����jG�i�R������w�ڱ�n�8}�2�D�� J������xu������ӆn�LN�Pc�.o�����`|C6�d�7)6�
� �������}�>l�G���O��Ox��R:Z@KGb�L_"|���l��%�i8�Tz�8ّb�����x����奃LP%bS�T�u�Y��y[dL����_O8p��X^����hdg,�\���Ԇ�qT;	!��B�&�lv���.�ȢWOk�H�4��b�W����m#M�un���L��!lj�֙��lo������>A:Z��6��y����A`̒�GX�����C�����f|n�����֏t<{�q�pr�����?�[�N_ߺ���i/*�w_��˭7=�~b���x�E�O{n�����x~�}�����4~�a����/��ܺs��=���Ͼ����n������L+��WlV7w��~�����?����;E�<�]�p�~u7�I^�
_g�t�S65�fX�&� ڷ��)�ߢi8�����!l����½�J_��o?1l�,W�F�d��f��ќ��2�ٶf�
���IfLC���t���3A
����8{�q�l���
D�yyѸ�Zƒ�dL�����h'�d��L�a��)'�f6�����(.v��d["���,��R��ҋ�O>Z��D����Dh)T�pC-��g���/d×̣B.v��z`x�h͝aF3�tpZ"�2F3KӎmC��
��/)f+6�iH�XF�^Lv5�;�	jJ�cX��h��ȅ��HJl�z��,{N�`���`�L\��p�F-��/Ȇ#kD����(�8)��Q�^�̞��ȉwX�Z_��,oY�.�:�5�s����Up
8�����fP�o
�&%v�3�8�D����Wg�1[g4�p|�^�1�B.�h��C�O�a��=����7)� ���2����c^y�M�D��]��0�m���:\Տϐk�si��8:�2��3$c��8�+#Q�)0�fT"�24 �&�P8�!'Q1�����gH��e�w�h�4!�jҕq�ˎ��1c�u�g�N�H����H���U�˞4:���\�%R��sU�a�!)�f��>;�^+#05��l�y�\嵥&m?�l+7Ge��e��A�SfCDɅ�^�W�U�B�'�[�"R�p��Sa!l!r��+WC4m�Ȫ22��n�:�dL|"�Od��aV0'�2r�$��(�B*��(#Z��KH�C��D�&$���1+��b���>$�$g�1AL`e�*>o�D�i��)*�!Z��8��a���p6p�M&C�*u	��9?�z4�ZA�>L!��4L4=��k߀��@ȫ7���\x!){WқJo�)h\��3�Z�X��C����b��W�T� $����l9u䍙�v�^"����e.�[7Y���b��0�{"�n5��5ko���L�c�����!3���i±�O;���/�]�/W.;�Ώd.�F}�,�o�77=��6����Nn�(M��M�p�¨yy��Ξ�����Y���s>z�g�ђ�1e��	�x��1P�G.�;ǥ��7�eٹ�꺽��4Ɖ˞>�|����fm�,�%r���ޥ]u��M�)���7'7s�_������Fw7��������a{�^��wMV��3��?q-�a�U�_?lyvp��t�0��#�W�k��C�>�s���2>|����������jp5^SL_���d��IڠzAC�L�CΆ��fؚ/dE%b�H�^�@�x�1v]�!U�IF[�F#B"����
�s�<��&*��e�)�%�7�[�~�VF�pv�UҼ�@H���sՎ�����&��)�7g�嵤35��g�KC�A��H�0OA�"��%>5��m��4,�l����n� �p�F���M�X���΄M�R!�T�C����K��-�/�,/0ܰ\����G�Myl.� -�J����1��1����b�6�?��?��_��k��+�54$���Խç�z�*,���(V����\l�)`J��7���!f�S_"���Њ��aXp`
le��"�j�񲹤�a[v��;z��܏g+5W��Q�d5Rl�6�����6��yրU�F��n��cµ��̘s�# !5�R.^��oM�|� �H��D�7/�O?�ԭ4.�5�h���vSS��n�p����7��D��CF`��z@�cӋ��z�����%��A;��'_�\����&_��;��������/�>ܜ�B��g�}�g3�_~����ً�g�ث�������������^�|��W���w�{��hu����f嫣�ˇ�si}�k�;盳g�ɯ���po�MP��\���M����ɔ
o;�/���w���gR.G6�v�MN������s��Ƴ&z�֊�Q
dn��Cb��Km㼃P:8B����ָ�����~���4�fs���NRj�S�R��1U�f�}� N��I�kJ��?�tک�� b��i�y�d�N\,�I1�\��eo���ās^�X�V�p=�E|k�~�-?Yo�;}$.��n��Ħtp���[�p�^F'�V�"[��Ϯ�WC��j5��l�lehd�2��p4�4�$���(^E���̀bźq�j�f�{)������裏���?������VU�Vf������h�hZ4gLY��{f4Ŷ��4���g.Y�CMB�e�{5!���r��7|�֤�q��z��}N��R��*��[3j��V�a"���qLA�e���[C4{����OY���]��!�U�Є[Fj�,4^�X�!�>oa��+)��,d+(��o�����7Ӧi����tD`�=�nC9W{Kt��|u��xK�9��χ��3��|\�{�>�?_�~�`v�C[^n�=�yvu{ྣ�_��#5���.��(���m�#_Zs鼢�˻�杓o���?~a�ٝ�����_����|<��jup���Zpv��f��3�}�ë���o���������{*o��nkl��o�4lKY�мƊ,mҬI������̀4�A�.��e���ض�n�B�۞�&Ycx�\,qC�fnML�J�"^���LV����>f{Dm��S���g��&��C:I�n�7�ѐ�;���P?�"N$2fkK��|��
��pR\l�Q%�q*H�Ko���K6�zʒ>�!AR=f!�
@��f�4F|�ʀ0��/i!Rk�p�H��9dD�/FTv٧Tٓ��e����Z�B�t�k�'~
\U[U�,*/[�6Պ5
A���i���W���8���U����f$�+$o��������������]���[R�a�x���jh�f��Ho"3�Q�Pd��S�i:��%j�����R���r��ɅSe�KPH�8u��\��]>$�8)7�<6�6���\o�z|=P
zH�x��HT��±�e�O�Y��%�D�gU�SM�R˨'n:���������Lg�p��˦�H�)Ր��I��>�)�	�n����G��^pG	��q*c�p�)�\x�����Ґ!8�7�5d=�����-2�A_gh�!54 ��L�P���CF�������C"�p��\�A=\����Y����4MJ����7�����}�ɠ��J=��Ҕ㳧N��6���!�
��� �a�@h�=$ͩVI8!	V���5�l�z��6��
��f..�h���i��K�+�1�JFFh��e���a��5y���B)ʢGX����V��0��5)�cS�@d/:!��75�p.d/���IC(/�?����h�G+u��~�e7�ӏϞF^=~�z��VR6��&2��4I\��G��1�J-������9~�d�՗��[{�L]:����=�������+��
��-�!q�քaC����Lo�15!���:+�\	R����RV����Ѐ�:������顑�������r����Hd�,�V=O�a�ua�󓮉z���%��ps����2��m�����c�ۧ������a|��75]^�E���vLg�t�8|�m��N��	�1#�&��~��}���U�m�H�%:^y��ĕ�q;q�s��k��9����5Ε�^�	�a��N�l���]��_�C��������W/���ۋ�ӳ��G�y~�
�������~�û���\������x�ŗ���{{��2��x�����+υ��x��|�x�䨌U;���9�[]�mG�A�c%�������S�ibh��L��1m4��+iP��Ȁ�7��8�~��,_���o�#M����厣�=�1g W)�ә4��	�)����kB��4sqй��B"�1�:	ܵDCdL������_-/��(���)���E�\ct$BM�BC�p��0��)�mC0整���UA^Spv�n:�ԉE�b�/#[�XR�ٵ������̫���Բ ��'H?R.�&[�R�z��UU�p�aKd^l���p:�Kg{٫}��:��DR@K�a�si1gO<GcScL~60���D�##<r�flx�&�,��[Ƣ<���_��D� �RvBo�%4�\m;^�(��������j61�A8���&7dW��(
���ԟNE�v���[��h@�@Ŕ�^"�M�2�[���e��LТY.C7��U��?����!�Z�����M���g=��GBzl�D�aWf;�U1id4UV\���\&��8hڲ��=����˄�/��K���ױ{I[�zn����y��2�:x�^]^��s5��{j����ܜl�4�x}��}��ɡ�5w7ۗo.�Ou�N_\y�&���~����p�s����Cɹz������+x9����׽h�]7�Ƨ��V7�1Z��7S� ���3��d{��vzQ�>��-����bn$XU�Z��ąClC�z�%e����>A6<&C+���	�`[��б�ۤW�������Z�ǩ�p
�����Ѐ�U%���#�5�8�h����d���T�(�DR�Z����y���l(�2&M /�2Jj����E!hՉ��g��'�n�O8h-��G���P���Ue{��ف�|�;��hs[|"b��ZÎ[
��gpUؘ�r:6M|�MSS��e�fRv9�JVߒ�hd�ih��4�d�ySN�tE��Df�S�\v{
���Φgo���A��O?�Y��@��b������V,�K�s��^��)W5��X>9b��n�f.1e�)�*����D�2�f�h�k�8�K
 ���ىd�SF����}����dT����Q���V�����?��j+4��
5$���j�t.±Ӓ��\�p�/J/Pal�)�Ra��T4R�G��B^��a�@���2��2D��8�0�Vw�����p��������׷7����zw��6��I}��\~�S�O��=�v~�7g>���������/��x��_���~��W�)�W�ٳ���#_z+��5�����}��w��zͺ��>ޜ��\�o_�=��    IDAT���up���w�Ym^�}�'��g�����W���Ƶnf�:0:މ�jg��3w�ű��m�B�@k��:S`[v��H���	�1E�"l�����\
y!I1�zdƬ���lm�˶��K3�@!��D3�ѫM��Qr�@:M$�%��fgL�������(�*5���]��U��̛~��x٢ꕝ2d�&ȆW��I?�z��^T�
���0*�����Ě>cV�B��t0�5H���犟TQ�Ek���J��4%6�D�� g��Rȥ��'q���PT���QFx�z^j��@�8��#�����)7�	��\�pUq-�X1�
�a��U�~��vd��)00� -)��G^�J,fv�%R"�6C�z��R�E���Q�\�@������pF�&�g4d�B�f�:��ZC�\�03�c�@-�W�������d�Ra�B"��Ԝ!q�6��\��j-N�41ā�0�a���X��v'������,!\^���ACF��2
/9#2��B��R\8���� � 0�=fH��^�ą��s
쪅�b�,�d
��d�L5Cv
��z��m���$����cG�oj�φm������ʋ�Po��I�@[�����SU8�Ma���[���T >�[Y��8#�L���J
��8��6�!����5Q ��l(D�啈w�	�������!#�2#�b ��oрh�����
�Yx!�Z�g>�����J��o'b�:�}Cٰ�f!��/i��]$�d�"R����q�Ѐh��R �D@�XF�y��r���4����lF�*�P����`����8B �c�X fF1"�
[�������C�q�ͦ\�4����m�����p6�[���(m��3�@���R	>�E+�}!�ic�)�[�Y@yKG�NK�Xᒶ�&�[K��9-��	�2��pԟ���T���$��mw���
l
d�]�Q!��pLC��$Xj����ȕ�K�c�4N�"#0)��D�_[~,s\;���O�#B�{�Ɔ�t��.\�X�Z�6eDa�����.ƺk�et�H�� ���Kc�u�qc�hQ�y`�f��֠-��ƾ�vH���g/\wE� ���q]����|u{���*\=<v6�@�Emo���(n�>�o���bO��{�R��Ǔ��*���v�B��U����G��ݸ7I��W��V�����z�:?ۜ�sv�?�雉O��.�����5���w�����o�=�d��v���f8���Y�#�x_�t!H�p�}O϶&Z.F�a�,p�0 ��a:m��q��%2;!��	�<V���uf�� !������q�R��c�X��D�aX���*L���Y��ԲIu� ��7x�A.��u���7-�D�N!e�}�'��K��پ)X7e��ݟ�!�p�_v4�	��)���������S����7:�6_e�$V���J� qi����D\*qu��{QΜ;w�#w���L_HK���x::Rs�����]e�����x٢�*�Y'��hjS�5Ld����G��k�(F��ԨM�����4H6������RL��'b���%�k�7qCkQ�^��
�N��^ȸ &e��W�,��
D3�k���);��|�8�'�r1��3�!e��UF��(���&"�:�m�6:}��1 
+\?���04����\����eL�zY%@e �n%���O��j�� �ʔb��M�UHQnC6#o}u�f�J�|�)�>���J�E��D{Y���xs}��ݱ�^Đ=R��~��������ۯ^�<ڭ��7/N�?>{��޳7���S�o%ܜ�6��w�����7����xv���>��x;~:ۗ'<x�����؎[�NU�.i_�|��_����ݻ�����z�ǿ^![h���%�����qu]ۍ��8kXU'!V�6���g"�����Ղw���c5�Um��j\r��D���[RC�&W�F�������֜&���A#�P�p^�@����Wb�4�G�Be�/jP���!��l3*�L��@C:	��)p�T�~��H�X`�в�Λ�-e�q8���ClӶ�j��gm-�p �Es3@m��y�_�[�)��I��l
r�dC�,2�'x�eh��A��@Fe�(�����͎�T�T޹ hDF̪%HNMc�1�.g��)`_+#}��й"}���+�=GS)���[% �('��]�A���'�-��r� 3xI�i0Sp��R�mL�>���0��(\�=�������(��'B_Ch!ΰhb�zM,����h8	8�1��j��(����؊�F�A�^�F P�Fj�a^�46q�[Æ\6A��,�!��eU͔�o`V�?)(Us����Y� �8ퟕ�0g�(���o���B.FP9�=��C��2|��Ͼ�|�|�����;��U:o^�.��:�_\=nOw>�yquy�����ig7�|�ԛ6�Zn�.��yf�§8��z��]|��_z����?_�1��������ˋ��_�g�p��O^޿���ݏ/��yv����[_~��_}�����?���p����f�2z2��-bF������dp�/P�>숰Zy+�1$��LSk�eaD���`;����^�Ј8�`9�TI$"c�o�Z���Kg�M.�B�ђ��d�.4-c��7]�z�DrgF�HU���Y��V�����6	��^` N�(�!)�R �Z [����S���h�bء'6f�j�(\_�����W4�ԢU3�����vC�0���լ���8�4_j���쩌(*���!���;�k���C����������4�Y[}ϞDc��k���[�Ib���R��D�D*��0�L`�a�c��S%��.Qd���VG81��2�5���KԪF�G���W���,�/)CQ�h"p5,#�Ns��]y�*e6�8�6D�o,{j�зe��S�P�t�y�9�P��2x�.�D�ERи��U��0=D���aʕZȐXJ�(А���p�����^lH=f��>�>��aj�4U���]l5��svy+�M-�1�)Y���d�'?�򌪰Q��%�b���%��I���5�R��B1�JQ�s^�"x�N��'}��KQ:�&S�QTC4�Sh�1r��m:�͔�>�\�\z`8)��5L��E@��ךS/���>�K�JA��=�w��C4.`{WY�Z�h4��q���2�.��@'���д�b����B(�b��B������6ᕔ;#}����*!��Y��fh�8�&�o����?�U2��<&�&G�5�v`ʘ�Z"!\�s���hS��~u���OJ�T!�eA�5�ʈ��� Zϼ�\��a�6D����D�2˕��h@H� �:p�͋9>��r��XjZ���^!�T!�BHYG_���0K�o/b8W8��5ۼD��t s:�z�(oX�0�¥���4Km�6��MA�S#�*.�t��m�e�3kc �P�h��8�fa��	�"፡��Z]�AHGϫǜ��N���y)�5�� � ���ó儸yHͭDw7��~9�/'[:{.r�=V�N�5�W8����z����F�r�px���[oOm�ۖn.�:�HK��[�<%��{�ˏ[V�/�u��R=������wǒ���x������?�y�}3� �zy���
*ty���Bjt�ֵbwO�ƥh�|NyY��4�6����<�59�6k�=z@f���k_�tz�cŻ��D�;�]޽x�]�͜=sq�#�˓����,�&�荟��<\=܍����z
�/u����c���:����I׵K�\�d�
5e�mgY�m��H��d��ͫ�E�xIAl�h@}�ױ��N���X����{y��zHF��Rpi
Ә�d,��������7�t⳹��hy��>�H�>A�9_C���G<X����kVñ����|y�A&�	A��eG��t�8	���1
4��?'�*�"S�k�+B�^a��6�����\Q	�/c(���C8�,PIp�ڄ��.Φ(���h�KFp���e^^;o�N�Pk��B?�������;5�M�q99e�U8gǨ�f�W�h���*qbQ�:2[3��z�zH��掟+0�b��dGf���8ZR�ʀ�I\|��-\3��]mCfkb��Tf8�ȷ��@g��R[��a)� 5�8E�L�>���&�(=�f���kg5�v���ï!�ў@P`I��K!I��.L.!�\�"s��!w�ӑ�Y^Ǡ]Z/�)�Em	�I�Y�%�˅-1��AkbC�o�!;Z�%����� /!^�R�J`��=�n��K���G^W�W��n�y�p5���r�����_]�����SO؜no.�����;/ޛ������O�Wo����������͕o<޼����w�����F��n�\���V�˝>�s�w7^����0]���Z�~�fGiA0�|B.7K̦l��$�����5���TQb�yq��"���E-k5�+2��Y[��#�m3�%�LJs�s[H������@}{�2$R�p�pC��W�ahp}!�.���Q��3�m��r1ʛf.`RM�
(i�Ӱ���mKq����f:'Ǥ���&���/Qǈ�d8
��є$����� G��=Y�,��/���P�&"@"��"+�)���z�J��?���q�6yU��Y�)���1{eš��Y��
��
��a���~t����Y���~�(���\�d��M�Qs�j$�U�áS������:�|��]�1�Zv�5�5M"j�8��:��&����=��$S�s�e�\i�r )C��Ӣ������=�Id"q�����'H�� ;N��	���(x.W�6bv�Q������t \!6#^��~����3~�V��v�/�L����zh���Z�촆f��b����B�A���FJ�z"\4!ȭp�]T
@!��4M3B�Fja�7 �wي��i�nWGg�޼���w><��]�z�����K_2���p������_�}����N݌t�܎_�=�ޗ�H��c�m��W��~��Ͽt\�|����/�ݭ}���S/`�'>vs�{B����g1�\���믎���G��f{�����//������g�����7�������f׬[Cs�iX��-�����@�a�wnh��E1(Xv�ak;45����<��V��H��T�J�'0��+�9(��m>�D8z.}�y!�V�4���B�UCR�hU���8�I�բ�ΙB캆�d�L͐���~�{Rh�xE�7�Ɏ@�����b��ɛr6��3+�")�;�@����I���?h��U�L�P��YTII���eU\y��y���\�!�&�O!YeDӳ��i�v�k^�R�;vf�D�g�A/D,�ƥ��4rU��ְ"g�S��ᘲT�@��
0d@�d#2 �j8gsN���(+���jY����0{K �&��睫DD�());d��o��IN�K�lQ1��pF������әʆ@�d�MG_=����`V	c_�Ub�a�%�Ј��\��K
ȌEk�"4��h������M�)�������$��.��2 ֭]��eO�~`:Y��l.!U�����I�!3�&RT���.��jk���BT�\5�5��b�����2�����1E��H'��N�j�!�h4#�/
M_�*`�Dɨ�zJ���''HAc�"欓���<�l�p-�
K��b����
���� ��QD �-bX`�bs�7�2ơ�v���:�"�K1�//�~�$!���-Z:@͐+�T0;���`[�H���0����!$���)i�l�22����ة1�Z�i�����Q5�a皁)�X�ΨU'd؅�g���B@cK��H3�Jb�A���Ч��K�bh�J�aXaL|C6$N��!y����B-��$���?C���hh�˶�JW`4��-'��n(o�JR�S�x.5�Z�t}�x8�o`%��@���S(����q��"���z�s�)���dK�+D?�UngKP�!@�#�(U�.A^�U��ғ�Wm0���%�%�!-[`y#4�&� �\I*a��A���5��KTG����� ��o<���K���<{�D�լ�!�,��7��rY����f��C���eQ��>�1�:�Oj.|�}{}wW����w��$=�㔾&i㖫��Y�������t�;^���=lVw[_�����1��6b�39��^��*�ǘ�7�cjo�m�㦬��D��G׃Ο�*�/]c��݃0w���z�pr���捋�^���G��_���_yc�g$]��|��X�7=�q�[b�{K��q��lõ��X��*�7+�^�p6Po{1�[�L��ԐC�5K!VSa
��lٵ �m\LpM��U5*� 8[^�Fy�pj���[���M���ӞC"���y�!#�ۤ��%�&~G�W'\3�M���ѱ���TܕU�؆��%�xMtB�ly�v
���o+O,��$$�a�ָ�ү`F��v_���LSS3�AA�ƀ#KQ1��]��l��v|�7k�H�t�Z���/���E �H�����QpK�֡F
M�֟Z�kh"z��#�>L��˂f"Z�Dh:LMR��>���W_H�I3�oë6�d��MS@X��vl��N�L:Ł&�f5��!�,OH�t�{K����Ud����QWK�����Ii�|��G�Z偲��" ���G�D�e��ȼs�p4;�����3{qw�b�+E�4:�!����_�����߹�/��3������?QU
�ԭ�Va�at@.M^�\8\rP���B��u?���Ѹ��n��/R���/BX�������W?��>��������vu~|��������n���z-�-��v���������W�+}|������������A�Q���p��[־������e���߻�m�������^�ojh�M�V�֦iM�����ݕ�4b�m�Ⱥ�e�B:G�BRs^���^
=�Ŵ�A��vF �C
(�@R�|����R�15.=r{��R��ҷ���C*�Ňh��/�ڤ���H!y���7�p}j��gS��������pT��̆X1�\���X+�}����N:@+)����ڦ���ٟ�ٟ���;����l�$	ǧ#E�m����S�JbXdRz��)�¨i���v��q�S,���p �Nh�[�
��p5�z5�D(���f�H�4_Q�'�l(u''s�i�	R�ϥ I5
*i�M�6"n��hn.����?T�?��?��B.��#��UX��S�1��j*�TS�E�Ǭ�&D�tԠ��?��cY�b��������Dx'h^q ��Zdj8�R0Cx+�(VT!	N�L����GïZ�>f�" �N�d!���G��ք�Rؽ�'�K���KQ����k�A#�\���Rȴ�.��aO#[�M�P�&��{�~x}�t��=��>9}�y����/>��_\���SSx���S��ݝ�x����S�+G�Ÿ��jw����>�y���g_��??��;=[]��>\�<?ұ9���׷��_�|���?����f�t�O~������Չך����O����Y���7�]�t�z��Î_�겼W\�(32e��jh��3f��ǶOjfj��2mc9. N284�����p�m ��L�v��8C}�y��qG�'r;[L��#��� ��@yS��T?Yj�eA慷{�i/�i���c&�獏�l������zL��xHj�%��j��V�aH�~�3��d�ĵ�􆉇�B�X|}�h�)0�8
�5̕�l`=2fŔ�&DCC��6�!>���+�z������9�h����P�\i&�%pfA��<���s�Q�\��W��p^m�-'D�	���l�1p:h��~"�pe�[U�)��"İ����)�a�I�p�r�q��Kc󦖍�o�n"���řjӜ
����G!�W:Mx���eNM G_���ͨ�E��T�9�|�3��E��E!�����m
�i۩(�T>���C    IDAT���p!�1��d`���}A��}��-���\��d)uI�~�5�J�v���!R!e����'�� Z����Ǝ�f5�ф�5L�32]@^}0�g�f�@ޖ���UR��ȳ�R�Gc��&�=C�����EX4�Hv�d�M�k�`��0j��)�.}x�ePc�
�kث�����J���Ĳ���{.8��Jf�-\���Z�KR�L�P�qJW^8r
�B8��Zy!��Ό	Ȼ?#�D�����W@s*C//W��E��aϡHs���g�͍� �&�1� ��GnY��J'<�} �N�~_��zK��d!�a���3��і���RL|ٵY3~xY
o�q5j���B�m�%����oO&�m?p���iX�4R��S��n3S;�D�?�Z"�Ss ������n��9|�V��%-�,%��IM_���lp7LM_���qٚ�*�Q2��)��q!����Rv��.����9�m����JAĵ:�h� �>i�2В�����uh�vr҈siiz���!M"ygpo�"��l�P��T.�,�ʴz�*AC)Q5�+ ��)F����N�./h���17��x����|t���-�jH�|童�|G,�e*xu��P��9.߮����oO%Z��+]�$�����N���Ɵ�3��#�_v_�w��IK�G��>�]��<7@O�]=:<��y����eY2nt��6Ǘ�y.t���c�tr3'��a{0�vB�����;���NS���l��w<X�zD�ts��M�\�\\>���yv|������)�oo������n��Ҫ'b�z��{_�k=�܊�g�#�ʭiy�ƝUwC��j|&~��t���|�Z�
�g�Y�c��62�e�c�e ��'M Wd{�}@�Iěq�Wr��hcM���F��9�$���N;��S�kA��S�}F.�f��O��ɬ`CQ��\fAM�|��_8�$�!#�϶,]*��?�c�76��e��
�*G� ٱ#-�ڜ�~���`Q�+;>&ܪ�_jo��KT�J���P���]����ɥ$C��@jl^x%148~�p]/�ƙ�n@3Z�dՀc��jCP�,^8�W��&�ΐ��YpQ�hj�_v4:8�M����V��q��t�(Q��� ��%���o"��LBH���1s�y!J=mH��զ�a�Ϩ�њ ����lC|6�f{��D���*1j�k8B،�����A�d�hVBe���7U%)'8�@��QLv�J��ҧL��4��A���Z�%�lK䬮9k��_���vo�E���,;	���@5ͧ"���ob��7=�rSԛ$\O�H5�E��
��p��5��f{�<$�5>��n��������G��f��W�������������s�����gW�[�,�{���6]�^����^��\;>=?E�^��:_�7�d�f�|p���㛗>��tz���s�;�ߌ�}��i�rQN��x��>�ah..�V�� ���a���Y^ۆHL�p��R�����������*
.V�!5C�|���}���E/W8�Ģ�YcH�\���8��)J�!����d+2���.HF�E��a�K!��VϬ?���r�g:v
�76��t&��м������GN"�ө��qD����Ue�~i/���i�)Xv�-�^==Ne��,��z��{9��*�5�����y��� U�_n��GHU�єE/�W/��Jǡ-�.#�G:��ġ�)�W��e���.Q鈕����0Y^���UN�"W{��a���)��]T�=_=݋��c�=��0��'���עiVҐ>)������`�p�&�wèL�f$� 㶮�@@+��R0edj��7dH�L͐M-\�������R��O2��@��`�͛2\�G�j@V�jm&��ǎ��Ô{W�*�|p+\Irс�Ҁ�m,�MO���p4^K��GY˦�*�^x�����I@�R��4}8�L-������osvG���OO�m����won?{u������W_�7,�ʗԌwq[W���w@V��\.�lo�4�OU� A@��>�>��˳����۵1��n��zq�;7ׯ����G:�0��w�q��kv����W�|ύ��G���ﳹ}~�xq���� �k���O�Y<}H�c�@���ho��ZXM����h6���1)�q,��l�������qdOh��L�h:p����0r/;��Rnoq�/��RDH��N�)�kB�������r����̛P��h�����3�~8�|cꑛfC�E�jh�ڤ�s����4�V�@�/���ְ^�V��#P����2үr��b��BNY�ǟy�gL��h��G�W���BK�f�E�>cS(V�$���t�%"�!��(
��e���H:JY���3:l!�Ce�)�PU�#D6��(�DSdȽM��OP_%���=R-d��Z`"L=:Z8Y?]M\8B�I��d �\�!�k��Sx|C�d�ESy!�h) �s��a8f��S.�8��0;�E��M#�y5��,չ�s5l��+��9g��ygv�����R3Jd�ΝA�֬I	� )����i��8ɦ�\�>\���%��RC���r����(�t�H�Xx�,PC=W�ت�Ǭ��A�5E�a&��) X
=��2��jBR ^R�4����J��)�4�Jڢ�k��e8]D��\j�:C�WL:\-�����"��}.�t�!{CQ��!�Y�?*�DUL�Şe�5�7���U�;J�����]8�� ��4!µ�bÅ@����MA���xq�e#h��ԢUF.J%�[^�Ne��_�~�ON\�~.5�F
�p��a �+CO�p�!��.#<�l�,	f�Cp 5R�b�j���e�&$2�%��6_1bNZ�^B�֧ Z�p��W����1�*d�e3R�g�m�4qf��U�C9��P�_�Ɩ����e/�a��e��CaWU�\|�2��d#�B(k�i�a��ݐ��� ���e $��>���;	\f=S9Z�e��2e��լ��mU�Ֆ�8fjl��+��e���^O��1x�7�#٥ W3�* �_D�"�=d&�FD�l�H��0��$�Dj�U�Ԥ0kX��^��\����X����9n)���~��s��DD�.��).�fz�����.�H�.�&����_<�7$�􋕻;�7kΞ��V���������$�`��8�W_{���_��'jy�]�~�����'�[�>q�>�j��������4�5����ݍ{�~�ҧ�m,�>��N�؎gL���ؚ;ۙ���d,�X�q<v�S�-�e�R�E�ʽ��[z�o����n�n��=�������=�۷��n}��/��Y��;Ǒm�6�8s�����i�aﴏ=W���8m`��M�M���o��+2[��D� [S���pLi�1,�B"�v���\)�'GԾZL|���t�%��� K��K0�^.`;-C��j�����G��%*M�~^����AJM�Z8�y�@Ả�v�P`�?��V���\�Mo�Ȩ!�mH�A��w���f¯}��VKa(���C^F��2v/��9���>v^"ͥˡ�0�N����Q6�@�A\�t��Y�P�M!&}��@�&�_jL��CMы��QՊ^"*��є�Ng]���ug��o^�ŚZF٥�ǁ0��
!�z��p4��3d��1]����9Z���0ZӬ�tr�#����0M�p|��"���S��%���@&b�#$嘭0o��ȮHQ� �k��jy�GVC��$�"륮�\�-��B1�R0I��h�K�_������/ #���"D*7��ÀP4�>.�l}�� JL4��8z�ƀ�
�3;����u�Q�;��倞���f����8�x��������_���o���7;_�~{�;��ٳ�����x���-����/��g����鸄|t{9�5���s���Y^�׏I?��Y^i߱�������K4~�ڇx\��_��hR��
eYf9v\��us��}"fI��mjm�V��ٵ����{�q
�$�����%��Y��r�X���ж�X��iݭ7x�,:��9�O*��(��T�!MH�lF.Q1!�l}�1��&���B�q Ԭ8i�"0�K4\r>���KD�a8� ׀t��ެ-�5����_�ұ��̺54jh��Fq>��6�~���}�{�uv��:[v:*'(C����AAOJ
4���E�iH��F��ʐ�%Y��^�5�JD�+� �j^����k2f�&��N�=Z��������'����i65�@�*��GZ�2�� ��@6.gZsL�˘X�U�fFp����ȧ������؟��'���c�%�~���ۓ�K%�����(L5���Ӑ�����j� [O�V^������EφT���Bz!Ee�����,$d?6�^Ñ�,#X=;5�j�h�J���%r�ܩ���m2!�z
@�M�d�ND8ǲCx1�E� ���N�M�:c��q�b�ؗ���UO!���z�a�*�x�ڽ|��`���W>{o�/Vg���g�^2.�R_��O/��ח>%�;���z}r~4~�;�q��o�x�u����?�~pv|sw�x{}�7F,����ի�g��n���·��{����������t}���_mƏen|����չ{퇧/>������ɳ����Q�Ձ�5�'W����Ҷ��M��ڔ_)�wk�:t�X%�@�p'��ɶ���Q�@��˅&*>�&�\@����DYs�p󪐾=����m(*����}&5ޘ��H�����58A [�*FQ�VFO�!@��Υ���W@C�1f�1}6c�?�R�g�6
�
a�-���b�E�n�_v`pN�`�8.��@�agc4k-���\�����گ6p�V�B* YKA�,XR�yٓ�E�*��l4�X�z�l.�p=<�ʘQֳ��ӏ X1�S�8��y[��cy'���������g^Lv��YRn�l!iF�����5�����ɏ	�g��k�h�J-Vo�,��
��V�a�@:IY���̥��p��e�� ��0֫�\͑�����m���P��=�es	���;�r����!h���iX�l���a̪�[.v|�Zk�[��Q9��:ǡ,h�PF���f̚���\������S�BE��Ն����B�SU���s)�pap�1JאH �E�8����ޚ$9�+����Ս	މ!Hi$�� 3=볏�<��s�63F�D�	�tw]3������r�Zv�����^{�GDfeDF�>�4њu�ih[�)�G. o��G�K��1(g�)Al�L�"!��qzQٲۦͱ��zM��6�6�O6��˦?�2�TR�� ���b�uNR+��3C���������𙺂�Ԭ�u+����8z����e�k8͐-)dHQ)7�%htE5\�G��69!�	Ή`N�W:�X=���mF�P�?p%�i[ϝX���Y/is�dP@.
�]m����©I��*��m�+vVn���Q@�觎a��er
�ڢ�S�ʔ��;}v�9+)����Ԭ=�����CR�R���A6~k55��(J��1C"W�\I�b���X�q�z��ƪ� ����
C*8M"�dy�Z䩀�[^6����Zv��2�e[�ɯ��S8��k����R�,�S[�ݩ�o.)G�\=�tD4�\05^�}|)\T�E��SF�KȬ>5m!>Y����H�YQ�˕~����a���Ѿ*���6|vٝ��az>��\����}�G��,�>���_�B��;�Z�scl��!_��ɔ���_�����Uil�����9��
ǳ�'�~������Ձ3.y���[Ax���2��to�SG�R�<�cd~�PM�����+��,¥̃c�l�R��@�x��J�������3�}���D��;�\�����b{�Y.���S��4�މJ�.[.�<���ӧ>��_�P�r���p{���S�,�ş�n��S��ᛗ�{Ǘ��EiK��w�P�������/o}��)�q7�5Lol kn�m�����J���2�C���R�Fjl���+���-����hY�q�.+{^�CF����A��@ch턆!��]4�ؼz=�6��D.�al��i(��w^�&�,no��O�i�"R^��B�EK������Q�r�/5A.v��Q*����%�8P�ۚ��54'0�Q^%м^-����D�\I���#�L������
3,Z�2"�*^��P��`�y�Re�!��"��(�1O�y��E?��C'��Ф�Fh��$4�.>P:^Q�8��#�ƆL��Բ�
T0�p�,p�D���޴S��Ќ�,�K@"�z���(��fYl��쪰��3�0P�6�l�\:��	��Z`�-˦�o�Da�*{S��r���aD.�K��+	褴�M� T��������.�����'��hU+����Mή�n$�Bkx
��*H �z�"1K� ����d��#�C�����'V~�l�*���ܡެ�Ǎ��P߂9�n^���ܾz��ju�ҳw~����x:�љ_i�~�� ����ّ���#l�_=w���w?����e�^�]g�UF��
���Ǚ���ӓ���~J�S�a..�fsl:C��f�j�8Έ�a1��܉�V��Ҹ��F��%���E�-�ȕm(�B"�|˃�_y.����?u)�2�(T^=�����њl�ya���t�0��@�	O<f�D������OG��,s'�&<�R;lK=�0��Vz��t�����>s��ã�N�Ο�m@��'?�B`HA����h���fAV�jKj�i��]X�t�y��ˆ�j�@!b�P=\���r����M��v �^���@M/5Z��H�kT$�%�'%���?��T���N�^�>��#�5�bO"i|d4��D�l�5#kkv�jƄ�q���.C6Ca8��կ,Aס1�Dg#����M�|E���l�E�x��[�\U�CE��$��^ټt��f q
�U�a[
�&��"4�'L���h�qi8p�e�p��F�E�p�1!�l/flA��oQ��S[�f��aC�S����e�Q�fu�2��W�A_8}C�g^��!�7�������,���c]�ׯn��/�{zr�I�[~�����c��W���N*�^���Ҫ��\{�������'[o${������x�ξ�ln�[�^y ���o��Dv�{���W����������n�=�[]��w>�����ps��ۯ�<Xݬo������Ʌ�g˞<>L�E�����Ǳ�M�����^�:�Q�fҢ�Un5Z4�͡��!�AG֘���D��@���,BjDD9�R�OA��
C+���F�s�ġ�����2������^=ySK�@�M��L��e$� ��i�@H!s��@�|)�y�p��E�o:�������E����~�q͹$I�2��y���|�!<�YC�Pn1ٌ���!X_=�d5F���l�
�����t�l�h��t8���Z74`�
0���j��HA�"�4`S���6E"+�A��)����@k�7;þ��FO_OdS8�����gG�Hy��K�_S|��[^6��P��T�lF����fl��h�0�l=�.��.�\Rjq,Ȭ9�v����"�.���V^[mw��IG�SF�D��#X�#0�D�(2�e^���]��fFC��ƥ�Ҁ���V0�@�XF�}#�b�LMjC-5W�!�9�嚥���s��Sa�!z�Ld�&��րm����и&�φT�z��Pn��'S*2N���+�[��� �/<A[��:I���ho��m�k�mL����~^����>����Z���36/0fF[�8R�w� �ҫ�v�!.��Z�p�ɡ���[�$�����O�-�Do���Z�8�4�ZxHR*Q^�
(�G��P+V�r/M��$��-���a��RH(���(ƴ#�oH�X.FHs�|�D����4:Z�Xp�G�E��D2X�ç    IDAT��S N��]�p���c�(uӉ#��@fh4�S��f�[U��諐�q�3��z�U��gF1b�BcO�U���E!�x�a�e��W K4��2�ln��$'��Ԇ��JS��E�+��#�j��J�t�sũ'G�g2x��-0N�!��q�A�.�D�O��s9����ٍ�K���˾�)�Q9�x|�+)RoF��p�2��p�ss@������R��J�ht zR�Q8q�:
�ס!d�?6�I���f�ȉOJ�5D(]!���f%���'�W����#s� ��O���⹾�HH�Y������<��y�%��S���U/[]�T����]_�^���>���q����G]�v��|����j=�Ν%f�"���~\
tu�F���oŜ����>P���������=�=?�a5:�D�z꡷>�{x���y����}�c^
���k�M�Z<��6�D��n��z��y��ypg�G%9=���!���OΜ"[=}�d�w{v����<;�?\m�������߹�껫;��<-��k���~���]��l�T~R�o��ZCr,��9�|�CQ%c���ἶ�^k3�DmPLv�H/ʮ+��`C��O.��1^��H�!��@�u� -���^���GqKyre3���O��@6W=�4ʢ����**��)�N��a��o��5�fCx�p~�ݜj�l��;)��G.�MV��>^C!�Rw�{��x'5���V�D,�p�D�\D��h�b�1ٽ�ASZ��T�7\�t	�ϦLӹP�D���:��q���4�p|Rjj j@dFӧ�+Y`5��H4�����TkE�K�( ��wj�)�ڇ~�%��2��)[�Q�c�\%R��!�C_��95�����[�	brU�V`�ć�S�3��2�VO�c�4��Ҽ�K��z��֜О�
km���"3(W�&i���Y0f8ðA��e �B�D@)Z��/��tZd{$xL��҉&eʆ��h�,B;�|�g5	ZX�#��ӓ���
���m���Y���@2BM��!������Fӫx�,���T�m9��ie�x�_`�>9�V;ެ�Mr���ŗ�}s���\��;�xz:��-�os�����컻���/o�nݼ��\��II���~����V�W��,��2N϶W������C��_Vet-��k�@���d�s{�m��B�xZɶ�'�"��p9�]�"Ehs�A6k�\�������0ͫ��_�OS0���h!t�#/.�,�(dF���jN�5A㥠�O�Qx}8��a�#W6>;M�F9#M.-<{WG��I�"֤������ֵI��Y�ߊl�}@s�X����g��/���_������eH!��\R��5�k*i�y�;�����5���gH��?��2Dm����.zCP���4�zyqL�v��q�����p{���o���S�2�@"�T%
BYm�����e��X����D�U�Y@�&E�T�\�ٍe� 45�#��d�v=�iR���q�������������B˨W��6��>�5{��#�W�tʫ$Ql�����_��"��BԬ�J�܅h����8��2R3DFcHԬg=��%�Gfh��6s�ip�8�^pk8�Gર��¹f:�����)���w
24�p}�Iε�^/N�f�K��*�=�; N��7�~�xr|tx}��z��_n���]üq�������߹�9�Q:�` ~ey}�>�4Z�ke���3� �P������c����ف���x1�'Ǟ\�':,���8��=7�O?<�{u��+Y����w���[��O������G.j��8�?�cm�iF-]ˢ�O����1e'dۥM��> �Ek($�u�L�}��ND+�Ƚ��&����ç�c����ګ�*q��5xF��@���iRI�f��2.�׮���(�2��XÐ:eG`�3���
�^^v"L�2i��	��l�8��Ѱ��
��e"���k��@.*}|m-+C�P���)�W���!2$N���u��U�8]�� 饉m��Kq�y���UUI�\2�$|�f���)�WƤ��t��	*�Ds�֐���&[�[`�PKS��K�2fj�*��K'A��aę��������OCT�^�ckNBI�6q�6Ax"��8\�l���?\oCS3CFQ����8J��Ԁ����K%�\�H�R��H�	�����qUI��������Έ�~Õ7��T�nI� ��F�l��Hގ )=��̾")�"р�D�,oI=���H�GzR�]^C.����j��³�)�W;<}�h�3����#�
�U��^x.vs)���ŔE^U���h�15CL��m�\3�4
Rٲؚ��P����Q��A�hz:!�iF�;�-����xG���ɜo]S�)/}�7/���Ka�ڬ���Ð�W/�7�>o��\��ϕ7�M��Q�^l��%/oʓ�@�d�`�W�FF0DP�G0\_�L��Ɇ�kU�3g6&�6�p�@��j@�3$�8B⨖�\��|#5"��ټ��P�~��������`
q$e/A+d��VF���0eA�kµ�\�I���\���\���5�D�����~1,/&��J���Y#�F��%*#/�R�2�q������,�D�!=�\��L�\yْ��_lH;�f8Cf�ԟ�����dd��~���8^�s�g ���/yݳ��ŻKdF�޼�%ρ;�Q@l��'q.]��ͮb&(K��FCU�\D���\�eT<C.=)d�����Z�[[xH��UOj���Vڥ�V����ݭ�6۸�����s�e�?_A\)��; �R/�����q�.m��Iۍ\1%���|����'gN0oԅ���Ԕ���,=��\�7���;F]�\~��v���9}���������^�߯�ܢ@ϷN��ߍ˔��c�W,u�p�L�i���4�Y�*<J�%Ȯ���<��N�t�����֝;��s��M�d����G���?\s~�MW{ۛw��n���'�����_m�/o�[����陓 .���z����2�-ⴶJ^���bh�+3�� a"p�mݾd���id.����Go� ({4}�I�٫��&�m����F�"�JQo�9����F:R&��րC=��z�?cw��W�G���7�����L��p�5Qj�E/���J�q�@�c%�Bʮ�����w^Y��@���������xYÉ3�22�h���,e�L5.C^F'0EI:ur� �xM�!���K+P��28�XHF��5C=�p���esU�ag�,�t��\f��d?���U���g��,l��By1!lm��8p"�,��B�W㍜��)j��m�)X��4.���!6'�+��)��m��I��ij�c(��Ŏ�ˋ�X.��%;!W�������!;MZӌ<STP
�A�]��W��W8�e�WR�] ��k4��S��Ssב�w����Y��Nz���9`P[���;>��*�"(^5�*ӫ5���b���ؙ<�x5F'7.�m�O/\�<wv�n�s��x�߾zq��������O��o.������'{���v?�l�o���o��zR�����ݫi�4���q�������C�z]=P�'�z����0C����t����֛�ٙ�^CЄ���-T4�\^h�h�-8Ͷ�'�=����	'"|^Xrz�F�h�92)MR�lMQ^,\�!�6j�����:!D$�g���A��@��T^:§� Po5�'�>�K�*	"���3�C��P��b�{)��h�A��3׺>��S��-����X���h���˙���/�J`���R��[�Ä�@G��<q�.�Q�!ʫ^G�Jؒ�\碵�!m8%! �!�t�	�lAH�h٬!m �l�� &�,
�<볰�кar���C�Y"��Ϋ	��z"."J�`�t�To���S 2M���Q�x�q�Հ���o&��:�e�w�-b�8^xl��V�eCSp���
���3r,)���PO�2��¥$�&Ȧ���m��C"okg�M!����.��{o�z��@)�)�2w�)ćZj�@C��,�@`���?9\UX_8�Τ�Mh=�P��i3q �X��O\9��ɓ3�/|s���[�^ޯ��_����7�/�x�ſ�?������W_y\�o��_��|�'�7w�����ܴ�r�����!��'���#p���b��o|�Yo7g��GG���~w��������s������{�sv������z�><��yy����k�������ܜ�޼�����@��?��l�_��L۬��m���c�-K�l/��j��%�e����\����wY˱��ʢ0��@8.jl50���t�2q�0���]bX��=Kޱ3��I$��UI�4L�"6��*.!��,5�b��i�v�	��U��]�y��7��&ˆ�P�e��#��5�4�i\b�y'eC��h)�� �T���hj��(�0r^6�\e�@��*LvR�S3f:m6>�Va����)kԊ�Em�Z�^�p�e�/N��
�ѥ' �I1��٢��[$�V�I���ۑ�S���=�W8ä^<�A�,�\��3��͆�]�c8P�V
6�V���q�f��%�Zqٙq�4��8Ճ	Ѹfv�S8SvF
!U^TL!����5�}�-�l�!�T�&JK��6[�p������M0��!�BG���h.@�I��I-����d!���y�A(;#��C�2p�ĳ�&�&��p�
��7�S0}}v"\Z�z`C���S n
��,/D+�L'�!C��,��`���#��В�H�w���� ї��~��In��L�Q5`QS�Ȕ� ꧩEf�ٝfYҜSFfW�TX�_�]I�z]��z��7\:�iR1����Ɲ�
g��C&��b������*A�dlX
��.����#��s�Y��`�Bؼ�\OQ@}�µ'����YaD�\�@���.�PI�K��9g-2�Mi^e7�kNX���\�j+)�b|+��Qy�j� m�5�B��g���5����3������*	�6�9���!��\v�Zޔ�~%�2��S�'���͋g"Ub(���")jzd4�2KơƘ='�$ �x�z�=}����,u`Ql�d�E��ճ��}��4�ZT�^7��,�DB��$�%����C�g:��^Gs֖�׬!}�S:�\M�H�V�OgSDx��y�5�"m�2���%��S�y���������K��yC4$]f��
�B�� *0�+��1����2���`��G�b6�Ñjy��σ�=�}��"�[C��g�qWح�yP��9���뫥��(oT�s��8�s����@�5���y��+-�`������:�;��L�c��gґ�Ll,�dc+7�>x���>�m�L�V��N��Wۋ�����;g�h<�X�uy�)Fn��w��(�>=����{n^=�<{v������́_����s6y��_�{V���x#C0)u��N?/:v�Q��b2Vui�6b�
N��z:l��0Ⴇ`��$��ޡ���c-wn�7��lw[�D�H��1�(R�hh��eA��m��%��ʆ���ah����w� ěH�8t��()C46~��N!l`4`|k�	y~�ϩHgt{�[�Z('.ؘ���6���b���r���<) ���,���C�`'g�SdM�E��p�́��A��p��P%	���Eu��H����edP��2hK���e�Z��8�KB� b���Vۉq�ϕ!o�3��h��̹��8O�A�FMR2� �^H���Pޢ��Ȇ�29#���0e�@��g�)���e�2Ф�dkE�
A� �ϰ�l�b&>S0&N��ȏnnqj��߶��8�Wp�x� ���;vZvC�yE(J����P����������D;I\c+X��hv'���I��k��7-�����ЀQ���XY8�&�P7�f��Y}Z��F3T��F"wg./%�'gJ�ՠ��s�p댇ÎD��<�������{����}�������_�#gL��gepx|�т7w����ţ���ﶾ�������G�ǏQ�A��������N�����{~�+�vu�M��l��Y���x�jFS�[���j/D�'e3�i#ѱ����Þ�&D��,/}�Zp�y�N"!�.��N��^,��*���J �TP'�p�拯���k��*�4�"j��__2D���]W����b��֗�P[
WS,�f?b�����t��'�|bgn����b�{"b���?��wAOU5tg�cD�k�]��u�*@#�T�z.�+@+����i��?���w/�I��5Y5�'��t}6}�4�\B�Է�Ku�M�:
�" �h�^w��1��W�&�n��ڸf��+{�o�f�v�ѵ[L�8N��nIGl�w2)� �ҋ)�@��&�k3!�:��b���cG1�\�l�@�A���hC+�W��)���3�ؾ�!/q�} �n6L5+OU-5����)H�kǙ�!�7�3��hNfj�L'��pD>���H6Q����M0A�G�BkR��	�,pn8B�\�īy�$b�Ak��]���
K�A����=��� �_\�~����/����������?�q{w��������w���?r���������ݭ��B�.��xM��~u��{5�&s��������.�.�O����yt��omo��w�G�=����'�/|ufs��w�y���G��o�z��'���z���z��'w��䋛��ۇKWL}��Ah9��[�<'8�GIv9���@�]l���(ʖuP̭h�,�=��w8h��M/&5x�2�SODis8�(����n��l���%%��M� g˨�6�ޮ'%v*��H3Wx
!)O<0�<��Pc�J'o!���a�Y���WP��[+�V8���SD��X�Y�e�ÅN5�&V�BC�(H.��.0|��Bkl���مH'��˥��e�@,B5,fd���@�C������		���	G��y�{�7L_�B�8����ra2g dWR�q��Z�B�Z|L�u0�q�o抜W
��6媂��x3 B�1��"�5�e�ӄ���d�W@�^j0+;�4�'�f��e�P:^D�3�%ոp�I����;~��"�jPI�ؒ��ؘZ{#��d����k�h�B�YF ���7�Z��l �P\8�&��K!D񢖄�K�!V?��O^:�ȴ�j.���.����q�hR[�Fȩ遼=/PÉ߂7٩�ɞ�$n�Z˞C$>�1�e�!2�t�C� ��"zQ��  ��wfuå���	�_jöu!y��Fl�Bp�!�̹��"D�*:\��bD`4���F�Mߔ��f�� ή/��T���q���,!�flF��g�V4g1M�t\��o"���*���䚸�/|��^�d�4�邤������;;^CM`!�h���s,8}��1J�ak8����R'�m&��k�����d$�୪lyB���m�����e�rC.4|��r��s���hE��+�8!zdHu�'��p1xcB��˗+$��J���:�����Q2f3��Rvj�8��A0k�s�Xxd�?�ح�4�ħ���U,�(8o�� H�t�L��Sl��fY�z��鴼�1�����3��_�v9��uR§�%hL�8��"4�*��I�@'s�D�pJ'�P�lF+�0d�i�)Wmg0&D��Da���dy1S��țK�0�����Q?��5q��F.N׽�5׸wcY�qn�kQ���/�J�޻w� 2w����U���]KbuVW7w{#��x���/⮈���������o�?��ObJ�H_.^Y����+��vcA�v�u�Yi7��=�v{�:+1�b���?N�B�	���]��t��W�}�ٯ�!ȼ���{���ӷ=5��~�u�ăg��7�g��t�vu�U�����P?��	�G>���N�����    IDATl�\�xx����nuyu�⬋���֞wt�J��G�.kk#��o{����熶Mۈ8c����z.�f�1�>��Y��X8��91������ސ`{~���a4����Z[Q�3[�h��e��s��^��bTp�"J7'��6�f ��O���1�Ub5�ku��9F'R<��)�`R-/B'�[.�p^.��z�1��𳀶�����h�8�ͅ�G�~��eKW
QϦG2�cQ?b�f(�z�pF/�z��dt�BM�*���K�8����F����0�"�i) f�x�USP��N՚��O��Ze�G_^󭰙��FVC88�p=r����
�1b�2�B�~"�f'��и"�*�,Ðў4�ч3�3r�!��� �I^,YI˵p��U|[��� ����8t4��d�\���ш�	WO8q�p`���E_ô����j.�K���Dｌ{E��n��; E������ǝR�������Nl�TI�b������ZY��A)��A���R������d�Fʁm��7N�չG�{h�_e����c��:��7w�W/���|���j���o��� ��=�l��ӭ�y��Ȟ��Ks�ۇ�gO=~�������s��M����;yut��ո��{LH뗳�N���C�p�2��X%�c�`:M>g4A7�fʫ��I.6r.|
d]챀�j+�9�#3�/03��UB��!�RS��ʨN�ul/
��3ή�D ���ji�+�/$���e��k͗Q <�Vl�!@�&K:���K�7��͕>C�Z^h��M����M������g�y������Q�w��?�{4!�Te�]�tht���WƒB�T�%�bK�s�M"[Е	�]R�M�Ԑ-����1E��V&���p�QkX.��eMj����W}�ڐ��f ���8��@�y��!��UQ��� e$NG�y%X٤Ѐ�n���@4
�^XI���OMm�����JM��^
�y�8�������C�
[3u�k"�m��>��@RR7A�kMZ8>�!���"k�7�4�Pk��5�a^òL$|���(�P�E:) �ϼ�K��aF���3-��2/��V^�a��*�N��~��Bf���o�3�!]!8���H0�@��p��=~:c�Pw�������W/?���7W/�����߼|qw{���;������ݭ4�6w�������}������9�����o��'�����0o|;8{��?z��?��sW����<:������ߜ<�=ܾ���:�H��[2_}����_��W�_o���So1G��v���v0���Z�6��may[�u|���ж�g��x��m5Y\�WQ^�d�ZR�V5��E��%�P�*`���4�z=&[�f #�[�dc1����mQz�G��d�q�ڼ�S��[s��So��8[ňBc��(/~��4�D��s�"bKě,�t8S���ŘE
���\�"�5�Zvx�������R�*I�g#�4M����8iΨɄ�Q%��jt�g��	�k6P�����O���Fï����-��p�)��X��<[-D��,J_�@!�fdϤņāĤ�I$��b�ֳB��4H �����8��,հ��~�T_l�3u�������R�
��w�^pb"3�͢(��%�����f
TaQe#8�08�$Xm8��(J���iG���<�1�#jw
I�W�~��j�M��1ZƐꏓ8D��v���5a��~(��8cSַp!���L3<��p:����Z�7�T?�~��dw�M��&��&`�&*o`
�@؅H2��P�#h�tR�KG_8���s(�лd�إ����y8�fG �%I�H�g��D8$/�Po��Vxx4}�7pr��XM%B�
!I��
G�Ҧ�BI�t
��(٢��)D(�X��O�=3��;qF��3Ԭ�)%PsR���lѷ�hv�ʲ�YvC`������!�(I�IC�.�8�Vr(>fd�����@������j��[�y5RljVOvHL=r�E�X�W�,�-���)�L3|��/2�ƫq���u���@��'�հ>& U@��c����kG��N�B*�a��<���!{n�V��5�!l��ZC!�z�p
�J��ir,d*0jJ�ތ]f
���h
�R2���@CL��nˆ ���:�C}
^����Pƶoje�BPv�%�=@Xmz
�dٌ�l=[������t��9
{�2�����"!��v���'�#G`;Ga�%ѡ[}
p*�s`ݔ��F�=��,|g�eD���w(�`���x�������85`��ިȸ@����<T�L� �O��)K�w`:�jG8؜,�m��u֣�ƥN?�9�&�a��om�����Ə��=?�m��ٶ{�k�=ʈ��K��n.���q?�r�%P��M;Vrk.E0����������k�={i�t�]K�����mO��~��/�]��?�?8r�� 8e�}}N�����]��wg'�g.��7��;m��4~TG��窭�Z��A��FI˟����>06ق�!��w^$m��x�&C�%K����1daD�{��B�sR�vK��[)K]�&*�F�d腠I�����Ɯ��f`��?+�Q���Rj�6���\��#��YEpv����5w�ϥs�W
RD�^�dڂ
�",�5D���5�+K�b����4��k�9F^M.!z��[�����@�����i��,�Rip�y���<�N�+�˖E�`�.ٖ׍�
%��@Mc��ڼ3��\z�D��
fx�&��wq�3��ʫrRl��h�(grA�C��x��3��{j�b�f�		�-ov/�
�F����Z��(L�A?<0|ޤؚ�f�7���B�����l),>��"H�,��:���j�G6�؁4�>�yA���5.H=����UUG���n��k&�W�t�׮��2��v �=�Q<��O���|yڃ H�(�IƔF��o28D�p
�KR�:ZK`nvwQ+�}rr�`R�j풲�����:s}s{������?��o^v��o�}�2�������W㺅G��l������с���ѭ��.�z������������_y^�^{�[o���=����p�?w�5��Ԭo.�e
1��f'�m�����&�ԣ̞��"�fIM��j�ta�bÑ8�Bl��{ъW �&�a�;7\C=��(D_��eЧlز��!�MD���gK�pQz�P,��Y�g���A��D깦#)F;��ys=�E����w���'�൒��|�������bC;�]Cv{�զ�]�&����;�f�ۂ�(������.�j�\s�9�I��f���g���=s��t��H�]g�AV3͹ h��T�X�p0W9"D�D
�yU��^a@��7/�?����t���yy�S"[�^��X�J&n��܅�"�/�YF���wy��"������pڏ>���'V1�m�C=��=A�C�dCLК`��f�h�� �\7jt�J 2o+FJ��	��hZFoL6�3��@!��G��jg���q�.|}y+l��Ӭ�hl��]����e�*EB��Eh�+u��4jS:�����J��Y���W��&C�Ic��������|ݪ{����|�\������뗗w��ݍK�q����r�z�[��{���3^���=;wW�'���f�p����<&g���}of}�s��ӓ�'?�ُ�������ϼ?C���'��C������?���_^�����WϿ��������.?���;ܾ�v���iӛ����Ƭ�\k�h�b���l�lMUB�z���[D�%Ё@?)LC=/�a��q��#�����A0LDώ�K<�hq��̋���,6�*�A�W#~C����cٟ!�Ɛ^=����Z^r�ԦN�s��p���GAK���iB�����)5��-��@F��j�J8�zv�o�"����R�\����R���D�k��E�B,D�Ѧ�(�	Bp�gāN���ȥk���2��U��\��!j�f>W��J�!p�����!p�
�񽨦�T�p�| �,@6M`�2Ԓ-*;)L!�B.M�iT���@f7��ǯ'KSF���FB��/X�8�Z�%dw^^�A�a34��Y�*W }�Y�@�m��?u*�\C}ɥǬ�9�\U�&�yV@u楬U��}�e6��PaE&.�:!���1s-c�C�!�AT�GX�-W��h�5W���y���E'�����R�\���׮l�R�:�0�!�ljr)B��`�h�&����ΐE
�1B�8�-�}FP+]R�R#��BH��>�3�~����Ѿ�t�CHiŊjXF}�D�1p�F�+��2&��(�@H�KI�*<Ng��,\��"k	2v��F�ӰՎ?��M���EUC�$*�!C������!>������D�'(R���kI�C߮%]jD�4�ҵ�x��R��������)�����ό�M�J"��3d7�Of�@��b�l�,#f��!pC��2#N^��OJ�ŌPI3�(=�嵧��c?Y"��)B�-$|��v�dqf���͝�6�\��j���:���ZC��>�RУi�������4wE��Bp4jzH
ɖhvt�q2x��ц�㦟���=�E�!K��#W�ZQzd�݃U��+�7���zታM�v��>}�ᇽ��"ќ1�A�i�Ī'�ʠ��n+����u�"�"����{�r��@"leQ�z�D|�:g9��/��+�2M|y����>:Y.����a�E#!���~�r���t\��U�+���s 
p�:Ju���$�.���B�޺�n����[&��k�r����ᮨ��IŻ<8�bS.�B�����͓�{�Y�׎����c����o�����Ry��+�n�v�W�NE�C���47+�2�����n"7�^�������/n��7+_m�=|�c�sz��닓�'���<�i���5.�޻a����eK�.V�m���PZ:H.s����g�q���������r9�h���:9�����Z��:_g����,II*6�^��gW��R�}��>o|}j)�/)�L����8l���X��s���Y^�3���ڜZ�Ν�����Ȋd�h�ƦÖB�@3M��!۬)T��B�+�w�RFS���E�k� ��k�2�U���#��CJ�B$rf�� �5L�t���vNH��8��
�RYY6� ���U!嘐�Z�� ��ѱ]4dgt��D�ٰCxYB
��e���7���N�dg
"�8�)��@T�e��ɛK�A�Ε���y-25�1�E�Nak�8�*)���2�g����
!��R�W\T��k�.$W�R�2�b3�@f�*/�,0���ց�`�uZR�(v�c�= �UCt$�\Ppy�[��
�������v����0�ɗ^�6�(8N�=�Se�A(��� �W�]�i�7ӱ ��r�ݭn}�`�p�{1��n��}�ŧ���������lO��������l���Ͼxqxp�λOO���
�G���x����c�]۸�O?�8?�C7�wG+����{�ǟ�N/�^�n���n���o��b����֔�l�vEX��,�YC�x�Mkz}��zی�ю�Ip[���##؎��4Km{����p!D�^�{l��*	W 80״�4�U��N\�rU��s!�)0Aé�A�fȅ\�%��J�4K���M��q}�%��>��풐R(FTo��կ<q�o��o\ݔ����eH�����k�PF�l+H4��|v��2Y�Mr�vzѼ�*VRd́��d��f����NlF��K���Kl��o�"f15L�0�'VF8�����r!kh��82BA`6�D \�^d�gd�j3}F����%r���FK�%ɵLW5:dcq���_Jg��r�ge��,�B������mg������1e�#Uh�MG Т5��Wy���y����G^UI�����K���Z���e�Ԭf|���[`����L!&P`7<>6>��!��U�E!x�8����(����_/\1�d�U�pMl��c����0�j��,9~�r\}|r��嫛k�#�ȗ�ݮo/=+g��|/o=�|������n���~y{��=^����*�m������>��==mώO��>'��eGg�o��_�l����fߣ��׫�W��_���_����oo����ܼ��������o~���~sy�����zx泜G��k�.g�)�Ekjl���XF�v+c��h���a�s�ۓ���\��b��-�2Bp��Um\@�eeeJ
aӰ��J�8lF��T8C�l�pCx�j�g�ԘM�R��[1�Ϙ��6�7�@�V1ͮ83/�P��hzކp��jx�*2��Rh�"L&[8<M!�EU PH��@��9��v��l�Y�js��Չ�¶J������JńP�����Ea�G?��6��#�"��UK
��DR�Me�a�tI��"«ń�y!\��Y|7{�B�@3�P|���#<Y}�Ԉ��s�vhWF��E+��F�%��L�0��T�ڌGx􌽺
��oC0���ת.D����E�Q���aό�F��f����� *>[�p�=P�o��T�^�����S��ZX݅d���� 8ɖE?����!�v`Y�R3Ԛf5W0��dK]�	N?�1�	� �H�1ŭ!N!}tU�6]������<���hl����j#������7���&�@`�e4�i������W���]�Qd�l���l��W|�Τ�v%��i
�S���G0L<\o�L�\*)QU�b�s	���feDӧ�[me�3f�Gϥ�=���H��dٻ����,�7��g7ԋm�`'%�fvq�1�y��!Z=f!����B"d̗&�Q�bs�[�2ƤS��F\T)˂�!�WO��/�=�"H�L���!����F❕�09�zR6��I�}k�P	&U���)���P3C���&��^
^�p:殧_=\�����)u�a��%��)��6=�W�N%^�fv�Y�L:A�ͫ
WSH���7J5�8���
g�ak���CPT��2�(=�H���y�~���]ev�e�#�)Dv���1��
fL{��Z:�ҥ������[[�;�'�<�O�@kg�3�1�)em�~�f�[I���>e�"Rm�F��:7��,5���i�,�����'���}c�~�j'+X�jjb�kO��o"����6V�uD�+]��-�����W�5L��@�Z汓��_���e�r�혚����}�c
��=���Z��:����Z�|���� >WK�g'݃�c�߳|{9��[�(<�	����m�G�ݙ��������������{{�-A�r�؇��G���ͽõO�na��Ԭ����Ʊ����n\ u��ם0�7{N����'�g��|�:���u��x���N����ϧ��Z�^_=��S�՝J�w�f=�ϳ �.No���wq���w��n����]fl[WTi�F-&�ZYCU�H6��g��I�*��8�(�nɦ�Ԣ��q,8�c�}&�(�t9pd� �pC��������Z.��'�]�K�_�ȭ�t�첋*K�s�Z.`-N���2R�2�9��߰�w���Z+놓Bj@��h�0pح�jmehm�p+ܤ��2�s�L
��$�A��Wd"4+;!�3ձ��j�T�U�D ����LM��*�f�8N��թ�5L�M�MT����,{u�*�m.d���[y�_y��SS!��K��W6A �F-/\Ac��&^oC-�^lRՠ7DH�P�K�a)�����2�R�L�@K��9.�#ӄ�ij�W��+���P�z4��b#�)h��0
A�*R��,d�S+P�Th
�{^�8��&���D.#W�L��	Mkg��Y�N��m�p���({ЭJ�k.p͚���*��g�P��ˡ�!*=���"����A���ƞk9�l�@���(���b    IDAT��sz�7_�z�t�zMh���f�������ϕ}�?^}�����|��g�����^�>���w��T�w�~����q�t3>Ҹ�쌤�<?���Ξ�����������'O���y��q^^��&�q��r��O�*o^\lSV<�0#�5��[M���X[w�2\t� -��^0�M�:�m�j�"�4�7�]�h�͖��%-�5i���
oR����j�KU��v9\�&��Ť�O�Y��	)dW��l� k��r�,l�Ѯt�����<)u��z�������W���<~"�ߵ.F��Ű�[m)Z"���tl[Ͱ���v��ׂ�u�Y8>��c*��-�(�wYC4�4MJ:���K�
M��a-fk���Շ�!;Wۻ)5CY�^S@R�!�KoF@�8�S����e4�z1��Z;����B�����ճ6��s����4&�>�Ҭ��T��ۀb���a�jr	�N�}���>��S�L���E��U/z������;>�KGyb)�N� �^!W��2Blh��4_.�3ڠ�	)PO�8;����244=W�\OC6�5��I�j#L��撈]�q��*�^�u���A�B;��l`�2V�^��1b
�Z�$̨DR�僛E���(z;.G�������ju����w�~?s�����S_&�=����MV�x�}�'7�H�K�k?�����/�{e�����������s�ʼ�ߐY�����ŷ��������������ϼ��߾������������������/>��եo�ݸ ����G��}_�+`"�fm=����Ԗ֚d�[ ۂ೭����k֡�c�!�v`Q�D�q�ǂ�9D_"=&�Q�.\�ʧ����%���1u�y��L��@��%�A,f%Q��h��˅�a6��E#+ooUq�,@C�6�R��p����&�2�+ �����e�I��W[R!�����^3�O�j�6��dӟ��@�ؤ�!S�8���P�o���^��&��YH.k�<�ǆ�Y����@=<�!D��/�)3�f�L��aj^�,jk� ����3�#�gxI�R�ܣ�R�n��i:6�g"������*Q����>0�f5rч���0JԐ2���I5��Y$f�`S.;D������悀/�EcC(��	ID��PaeɆk�L�H�+A�B�]��5aG@��G��Q�Ԅh�M�@^���(��Eo�9M�~�?�q�[ǯN}
��Pk�F!hm��e��f��ؕ�y&��B«�lۅ1C�R��� �-��� KQ��c�ʛaFEЋ�)�8�p�,�:@��y3bNYxU����-z�C�l8�%��m_���и�$C���d��`3��a�]8BWF�,?L�b�/c"�
�c&2��g��+`�=h�jXl)�s�r�5٤�2�/o��8t�e30��t�I;���3M6>&���-F��O�
��K�֪�8��Ks�<���[��M�W,r�Y�c�t&��Wĩ�R@*IOJҊ1����	�S�\�/P_x�fQ�4��^�=i�p4�\s��i���M<B���fDH"{��t�-5���I�0��n���b(;�ϩ��R0&R`��)�N0q��KlC����b٘왋B����� �Vf��m+�z��fR�7WS��ND�E24�J�[�K�� Vd}.�I�h�@��3\s4��%gLS��,v���(�(��V�
~��_�+p6���X�O�J���P� ��i���Gv �&��)x͟!RT�G�`���Qv8L�y���l������ߡt5ѕBc!�tc�xJ������e���z�,�+�����9]u53� v�o���<�n{���`�k��ki��c��n}��$-YN=������o<mϖg]����e������'�{��nq�w����������p\k]�{�;|X�<==9<{q}{~����ə�9�ݚrOx�"�h5�#2�ãqrw�/��]��w��ڤ)^��{����={�t������%�S?=���틗_}����jN�_��x���O�{��j<�w�����c�F����8<�<��ߞ:w�T���z��Ă��z��@��6Z�|6�׮¶�f���e/�'�� U;�6�ݩ=���u�8Ț@v����!8�儕^�հx�ɺ�&Ɏ���W���!DiD 4J&jyыL�z��L�#3m&J 4�8�议}�_��3
k��8~��Gܸ���撡ߍ�=}���됁�Vay��0���t* �7Y�$J�?6��Y%���D\vyܥ�ak�s��,0�Z`�FGF������ QZ�R�;�o�z����D"dj���(��\;�2�ֶG
�8^�]��8��,����<�hl�jC�s\��2��t�t������V���da�k��L8#M���]�%h�L�L����WvR5CM�jwW.E:۴�t-,��Dz�*�p�P�hpy�%1"*@�y�UT�e���js�}����i�S6�`I&�눷������ y-��f(M%�*DO����3���4���U?N4L
R0:(�!��E"C.�'���XUI��Ņ��r��B��X���7��8�G>�����Eya����:V*�K�Yz.�����6��)=)4M�d8�������%�o�x]Cmϳ�K��}��ӓ�g��y��/_��W�����������q������'�E<{�����ə�N������ޖ��+�N�N{s���'$G�w.�&��_��>�|���nM��Р�f�f��T�_��}<E04�ť�2@�G�c��2W��,���`��k�3m��Kߍ1�-���*�<�1���U�ְ���g�*n�e�G�Ł�yI�q��J�[N���-c8DS�����q�fvN�#�'�>��s�ݝ3��/�7�����G?rSʉ�eU=ںM�\N���-C��#�p�j=Q	tc��3Y�t�\�d�*���2�.�A�i���@��4U!pɥ6Y���,=�54��Tϖ�������Z+D�J��#P.v5�y��i;yqH��	2������a^֪J�OA3��e[|D=�9��վWVo���f��E�fx�#4n�;_���ʽm[��@s/SR
�:�Pٚ����ӱ�h�AM1��,��iX
[7j�ȭ��谉(�A`������[F�	�U�kȈ�m��T
�5Hڌ���Q��L5Hސ)R=���|1�ch���H鿕88&͖� h�z��)l�d�!��'�z�����oon�o�̏��bvu���iڔ>�o��½�e^o��%ޛ�km<�z��u�!Λ�󓋣S?�q���;��;;=���|y���/�����w�����y��������ƻ��oo��\�^���z�Ϊ��Z�E[s�ҷg�Y�߼V��y��w���ov�4�^H+OVka=juZ=N�&)"��D@뱈�:��k+J���a����M�u��J5$���j�*�0��M_?��%J6�.���4SKP�!���a|H5$k�)襈)\�!~�bӏ?LFv%��ޒfG`3�)D� Mͼ�@j���f���ͥl�z:�)C�Ė4A=�\�&~�U�By�rl.���Z+"\���Ȳ!�f�,�Ah�dӟ@���(g�o�WB C��*,�-6�p�(�V��av=�y�>e�Y.��o�2�8�:���se��y��	z�N
�G�h��#*�C0E��_>M�R��<k��R�ׄ7G�v�'���VF^�
CH�pCm�i�or�ݮ����ɖ}Rp�ER�D粩�8��U�U9�즳�o*���x����d!���?M��#�(˫/��pvˈ����Ja�ժB:X@�P�qC��c���1O6d������ͷ��tR�޲�s1���W'0 �!q�ʀ�+��ۈTo�$;���+�����њ�:Z�9�3Ñ��c���@�a5�a�3o!z.���Q-r��5Y��4EQc���·���V��MT��r��>��q�(���qu,��7�����5Q��c���Ӭ�JB�0�q
M|�k�U!i��xC��P����1#P�%��%*0�P�>��z��#[�,���xc��k�MF\l�t���
��4��գ��5rCC��ȻY ��	����n:!���:1k)�K�PHsW������*d���h\q��p�����l�`�W�v8�Z���Bf�R�VҼ�L��R����C�F,$M.�2�ò�sb����{6�K_3���������~�����-��̐�H�J�ټ^�{�� 0e�N�"��HP?u����ԧPU|x���r�yV�*�J�,+�H��Ґ�^.�>>&�C���5�Vs�ӭ>�ܲ ��5�d���ٵ�>��^��Pu�������ڮ��X���ӟ}����̿��+w7�hޞO��w�{���;{r����큫0���o�|�����w�Yك�YLWY��S��<=t�p����5����N�(?rO�K7�A4�~������?���Õ�^߻���M게�������>�	^�ؽT{�aƮ;~��w־�������yzs���"�W��|�������o~�����S��t�jOM>�������9{�xn�O�}�Oٸ�R�����|k����WK�.Ws�v�b�Qf/¶9m9e�˛y6$�ޡ� �r�!y����
�C�l{I_j"hZU�[�SFcl�@*)5ò�T MvF��g��ReA捣���jRT���&n�N�b��k�������*�]Nt��t�W���E�T}Y���~�4)����"ȅ��%�Y��qў�=���Չ�n".��@*Y^���hU��7b�&ʅV�e�>�%Pmj���hmHŪM�W �fH�H��j�q��e�hxm�@CLSpѕT��]g�@�����=ʥU<���P��j���E<&�Km��.]��E�0�JahIU��r����dA.6d���zћ2�&�n4�RW3g��Rp�4dW�gF�����P�����#�x5^=DOS`��S�M�j�����[
�x'Kk%�&Rl�h�Y�ns"cZ��b�@[N,���El��?v!�k��	���>��9#��<$fÉ�:lA�-��\r�AJ��(%C�� 3�\z!��8���VMb�	oL7]~^��7�߽�|�;OO�]]������_���룓��>{�������׿<�p��w��{<�>>xc��r���s���e�����_���|e�]��x�����}�����'o'��YIU�T�e4�@�7�CͽI5MQq٦��3Ď�v֢ќ3���ȁ�h�Cl�B���ԗ�Q�%eF��Hǫw4�5�jV$W"M^a��@��yټ!8b�D����ȮMlC�j����Ȧ�>�s�R|��'�h��g?k����͍�?��O��O[:+���Ä�ݣ��@:��ThsJM�������%��_��[�������$3bZv[S��\(� ����Z�=�@R�hj��5�x�hj�8f�S,ov!�hl4��\�v�iS����l`Q)�5���P�`8&�khR=@[b=�� ��NS�\�yfd���C��`m¥C����^���z�s�������Ú#N���z����ڬ}�ᕴcT4op�J�E^k���t!zMV@��2d���oX��է�0�!�&�m��">��h!�TH�\yc����b�o
�S	/W�¹�d�[%�z��ywS�pi�d;p���o�8��wׇ���w2����w�l}����z���:{�룽��NO真Y>b{x���+������S?���y���e���]P/����}�_(�
�w�^���Ȟ��H|��ȷ����ٱe_or����5O����� ��漘�!-c��h�8�� ��5��m}L��35�p/jqew�ږ����"g$��7��t�)�a��x�I�P`����4L9�&"���Z�*/*M�$PSF��2�w���ɫ$�YPh��t��)��2�H5wm@L��@}
��vVF,�(�����Q�WYR��������9�4L����	W[����e�,j�U�� q��V�bhOVX�ʘ�Y��#��0��B��se'�0�ͨ�F'C�'q�
K�z�Փ����@��34L��D�f�[ERf3��(�5}.��n"ri��(�:$�~"bSXB��Eŋ�Q�"NCj��Q��A0�/�WI�a����h��e)�F3�"�$R�v�0S��&Ux���|�ld���#TO Cc�jl!8�(}�)��(��F����F��N��.�א�>�����͋�VT.K׆���24�X���bA�QF��� S(�%*dp.`K�no�A�Py�f�B���1ڟ1���j��(ȥQ`�vn�4ğ/v�R6�:��5}uµ�gg��ń�mR�O�WKq��BH!�M��4��Eգ�S.p�_�jN��]����]��sѷ�� g@�V�!od��Q�K¢�5��o}Z:8/��IA��+��JZvGV�2P��AJ��Z���14��W3�<�y�I�r�/m̋Ia˶�K��ꄤ �7G��b!������q�h�Z�=r=�"d3�2
�D���!��R��0C���^1�p�ه���iF�S���1��EG�f�Է�S��a�4�"v\ͨ�d�UFfR+�ۃ����3 U.<>�a�͐-cx�X�$>�Hq���h��F/��f���ׄ�q�+ 2�����o}::�F�+�������CE�kȘe�6ف2N�B�|�"ks��UمjS��l2��k.���F�@.v�c��Q�_�&E�\���ݸ�(��/�l�������룄>���Q�AY��;>|rz�s�>�y}㍺N�Óc/�ף���x��N�������	�}�3�Ύ�y�ݧϟ��7��+I��7���y��f�t�l>8r�ӧB�������;>�yp�x���/yO���S��o���㡭�5������ݥ�G~��힥�w7隅E���m\�קK��ΫuZ]?&��ۋk*�<�{��d�U����ݛ��������=��~�i}��~��՞O9��ǧ���p���W�߼t\���Oώ�}*���r���;��t��n_7}׃�m���ߝq�`K�Km�
��h�\�MA��y�ؽ~w��#��P����}���7� �c��b�hZ�,=���%
�t6�"k�9Ô�?.�m�9�����B�	QL�l��YϨy$/W�,�s�m�(���zK���8W������2��ye�q,
o�Ѩ�t�* �M��P)|�([,����o)"��pg��W��t8.Z*Cl|���k�FS���j���Ij�x�b�b!z�k����ޞ*��Y�̅�����Rw��dY!r��iIKAG��g�bh�(��6��Ū������T'>��g`2��'Qv���0S��7/��W�b�֐,&!A.�٥fk�U��"�$M�j��,/q5 Dc 1�	0)�
#eH4>:%�Eb:��\�ų�9r�3�l�uZA\�o��d����Zj2���f?��o��Vu69ۈ���ū�v@
lP�!׸��Ph\l�z6C�6�U�u˞��\��Ù7��O���\=ܿ>����9ٻ{����-���ǣ���}�=������{�����a�oأ�@��\���Ɲۇ˓��{��Q���x�>Ƴ�ә���<�n5��$�<�Mo:�׷>zm�V�����q&���[l���jy���D�I9X������~���������J�JA^}�ԯ�m+cf�ǧЂP�w�AC|H����.v����� D��k���	A�Ɛ�#,�^a����~��������A!�3��>��?�#�:�ӟ���j�BN�)�7��,B�%��P�V�(��ɢ���3�!���z�g���� 	��)$�j͋Wj���kTk�$
���*�K�r1r	�[�ϒ�HBT� C��D���)�jښ���G��W��l.����&�d�!��    IDATSҫߊيbe�DH�>oq<4!#h�<�y��Y���GDR�M�oFBܭ��?�c7&�0t�ۮ��Q]6��	�ZZF�����yuDЀ&bct��,MR٤Z:Sc'o�Ѵf��D��s2x�J2���m�͗K+'��/52[k[�ŋA�D���=}���o���W/p��Z`8��#�7�->M�y���m�x����a�~}��~�ɋ��	���7+<^���������v��7��y��;i�{4=�a�/M��D�t�sߋ�'�=�������Ù�9����<>��p|�3����^�A�u;���ܧC������sb�j����������i����[��m?�8����� |z��`G1fc0��B���0dl�ڃ�S	�Ô�J�lk}����a�R�$�0E���U.��aC4��z��B�G��2Z��J�����E�7����d�����,F?/B�hzI�h��K��'�I�ĩ���OSKa�� =5L�^��
����*�)���6K�OMl=ڪcӟ@�֌�;�!��T'~��Ȉ+ b�Z"�ͥ�*˖�F3�2ā�΅����������${�DE�2��"��/D��hI�Sh^�"@�I����hDZ ;~��@���c���W�hB��E�I$d%q�W|ᆁ��+�-�-*Z���(T�a�fX�h�pY���q�J�Θ����8�i��Xͤ �SӇ�\��J�Na�8Փ>��0o�l�zF���\�&Ѹ�D`y�5<[��8��$&|���	��[�"�Gl6\=o�>�L�ß�I$>)���A���IR���Yd�bz������KY`yG�����D�2����2* �8@��S5��N^:�z!���'�j���"h@���v�s��0��r%^!�y�ǰ���c1I��
lX�fH�Q�a�Ϳ�2�eh�ru��=0�&��+�H	�CǐK+�h"h�Ù�
�Ų{8� �>�!�8�R�I�h���X�����!#�y��=FL4`��)�u:p`��e�"ZS��h!M���a�-}��["��rŬ���q�R"��"�p���X+��+L��pLF�p��`3��88b�SIH�EI��%�[%AR) C*`£5lm�<=M���8�8�^�vuS����f�qg.�hzmc�ä��k�ᕴ�fDm*��bvˣ&V���,�w�L3S!�h�$n��Uv�&�и��dP �͈N!^��:�����y�M3��R�k��bfPK_�-T����GgwG���=ز���Q�K�G�h!-��\b
��)NL�X���X�Є৩�Rt��T��M��'1��/�z��C���;��x���3_�us�՗_�v���֊��F��/+Q��5��'��M�'7����4��ǽ󗯯�.}�����Ţ����Q���,���K?��N���,������ON���f���+)��f��ɱK�ެ��ۻ||���W�\�^�3�>�47(�uk�؜֗0y�4�������T~��mO��ծ��~����~���0a��Q1��>�;}z����įo��������������������nn��ܛ=���c�; ��5]v\?n�-�:�nd�\��R��e[��P0��]��Q^�=pT�G,&�#��%2���㵝qiƗq�����`��厦��.p�0qw:	�I0�4�ٓt"HQk��H��ىoO'/�ݐ������7�S��e�){4jV�[�]�pIе; =��pg����=ؖ�&�b!j6$¶����6�B�]�+�㡉B:����-�$���i��%��i�Ԗl�JG�K"88��J�*.��N_1*� �(���s��n(�f�-�S@`��]mRR��p�)�򚂥�H��<y]������g�g]lW*�tʂ��p�ՠ	�$��KXo�Z�*�8�5�m��`�a׋�X�4�[���wǅS^g�O�8@�Vov1��Y�b�*[uo�����_oHD�oX��_��A���XH��ySMc7dw�!I3����f�hvM��Hj{$b��S��7b*ފ)��p���c�)��#����:�̮�֮��D�\�[qB�l!l�fb9��(
q���n]�.����q��Vo	<%�+�g'�W�~�_���;�� <@ÿ���\ܽ��]�GO����ޥ�컸��������M�r�F�W���OON�Լ;xܶ�Ņ��w0���楧勫o�_���Xf��pw�F[�sl*�՟���y�پ=䐆h�L�7MK�X|Y��2�=�@:lD��Z"�Ŧ�����\p�ZF˰���ɵ�7Qh�v�bM�RK�*8'��ag��/*eL;V�i��������Q�I���O���%ެdFN!Or�i	!k�̨H�l��9nXp������9�<-a�Z��D�储���Ёh�j����3�lI)�T���\�!�^�Z�	*L�@5gh�2�3���^�^CPs��DHR�S�,=�W0���4�Z6�1�AL����4�r`U�
th<�Y�O>��Q��6���٬��;b��h҇���c
$B��P"��(e��+�a7G�z��pI��HA��Q�!�H�f!�w���H�QxV�H%Ia�[6�p�l|���A�q��3k�a�D��jY��ç�z*�A����LƸ�蘻p�F�~ds��תN
?Y`^8����m�et�K$
�
��닫��/.�֍DQ_��r�r�΋���b��I��_
ٞ�W�������ǣgбOVޞ�~��Ko)��z�����j�_}�ҍ�[b��믿�ç�և��Ot�=�?y����w}���o��� Η���󫫵!��7���Bm�5��F��pL��&�+D���&0���T���y�OP,Cߙ�/�a�t��!�j�ah�D�,���¹����q�T��h�!�ʛ/0�8pC8Z��DG?![ਕE��ZUI�a�'B���zd`#�bՆ���-
!5H^â�<�N|@�VaUU:�=�w!j�&8Q��t�L?f���8���J��2F��@�@��$[�g8�ƖBIՠZKDg*D�jUF4.Q8����) h���i/RT����-���4-e��(g�@xEF(W�j �8;��";js�<�pi��`L���K������h:=l��8��r��I�ٛ��aZ"���T-��+�+M^�,�+U���j)��!#kȆd��Dї�@��Z�l��4�@�p˲��?cZ����[%�r1B0K
�i��%��-����
�-$X"��hz�8�q�G�(˖�j0����cS��``�V�2��1"�E�o1�*�:C(s\R'ت�f��#�Ճ�����85��p�l3�H��N�[�BH�G�A�[��(��ū�*��䂗(�Bd�L����p��+��_o��	�5�H_ϋÐ�!$�b�!N"���
L������!hY4�~�{�eԗ�	"4�VU��'����'N�Q���v����+�q���Ck�!�mؙR��#@�������L:L��3Y��3R�W@��`�4%�0���	�O��B��SfQ���1��/<^1�Q#Ő1�^.!@����4�)����z!�h��WF���fFzH��� ';c
����h�D&�a�2�9A�`VR^=)��K��Ûk7��+`����X٧f�2FR�3��ҬC!�b�$%)e�8�ǥ��ۿu���Ԕ�e��a�eɅIʹ�2��	&�P8e.H�����0}"�I��5�p��
���SH䤊��k�O�6K� r��c�ن��:9]W�|��6T^�������U�k�B�[s��ڳ�O����������:u}j��o�xYlv~is����͝����zy쓑k��~��_+����w(}]�����ZR�{�6���܈/::;�����k/��������������rԹ�>��Y?��#&�솩SťZ��z�a|'�ոU�����9��w}gҪs�*�j�N<�q��M*�0+���e`��]N�����ɳCW���|�������;��<�9v7��Ow���%��8~�˞������퟾�>޻{z|�'D�v�ԑ��i~Zԧjl�oe^kT����ѳ;�h\V�f�Ů��G!�h���=ks��h���+�zW�\�r��\���_F}v[��Rke�&�1��h����L����b����m�\��c�-�>fى'(���-z���dN.�]��%G��kB��rY���8����q]E^���2rQpa��u ���RU�k�Cy&:ф Ч�W$g7���lS���ӱ�Ԥ#(�!B��(��2Q��
YlQl����)�Rx|ū	���6|^�B̚ժM.We]˵2�7�]�&�IJxF����Ȟ1}�-0Z=<������,�u ����2������k9o������璵,���mo/�lC
���m)��Sk�q�f ���ع�!L��!�t��E"#��Ʈ��2$�8<[,qF`Y��r��c��p�s��t�=ܞ�m�h��8�D48�w-X:�ܝ���?y^�[p;�]CT�$�ZzMDˇ��1�G(V>v�
B�f'7$5|ЄM����I��������G�����+?z�⫗/}wދ�w|�����w���wYχ��	/��-���༸?��-�O����阇ۛ��U�O���>|<���X5���y�4_5��ͥ�-��<��µ��)�ѳ��P�t`���#X�BDY�j!q ��Z�2�]�A!�²��A��p�&^lN���?�
I'G�6k�&�,5vS(���D��*ŗ���b��m����a(;��Y}x�����?��C��js��y��>�(�@\� eMIRB�����4?��S�����Tk��d�憛�&r�$Y�&�g =�;��"4kjN�j�TG�A�l��2��!;�G�-�@^�쇎T�zC=�&��(Y�G��5����5��kX%�
�`"IYp+������4��ӯ<ˎ��!��	:�4"\�D�-TŨ�)��6��?���H����xm����({�q\��*y������nS#h�qY��k)"�JDZ
���ڦɅL��pBsd��nR���q����fq2� ov��<>�D^NJ�$����"#0B�w�р�,T3�/*2��l�W�F��ЄK��~��7�N��b^ܬNN���+����3Vm{~��ʋ��/_�z}zt��o�Y�l^�?yv{wuw{��	��pO�={��]���կ/^����[���ƣ�����;�<�~>�Mͣ�ӳgg����o~����Ǜ_���׿}�wI�i"S��(��tM��`�i�ہ:�&�I���5a���i%yS(!�����#X:�K����!M^�^I8j�)P/���pM��7.%A*l�А̫� ��OS����åc�(\�\��O��d���*/D,��f�pd��@��2�#��kVY�|��Vجy����2M�o��h�S�(�w�Ub����Ѵ&�%��$���(��¶G���g��5lv��\�r��B��'�d�y�5C� k�=��P/��8yK���Iߌ�ȥ��J8/&$M4Cx�#�(�V�A�V����3�B:!�p���fT��)��aX��Wye�q	TU!�����8����F�-iL%yJ*^l�������g��B���DzCMH���B4.��̋�A*Rl�Y�ۑB�Ϡ�?k5:�P�7�O`�^B���>z�V�pQ8�y�C��	I����1x�\tp�w��y#��H� 1� �W��F�y��gh8��e�i�����g�z�'W)�5 B)�)�+ͼz"d͝���f�+*�@})�����$2�����b�**[/�� �ky�@�d2j-��"���4���7�!�2"x̜!�%���!\�I7����Ӈ�j�����d �)<0�n����R4$��5L��ƖŐkh�l^x��&BG 0/|�~s�	�G�<6�4�Z�x�X���\� ��𿧋�,yGy��V��B8���p��a���#��)���]<;5}�5|��D*������+#�M���8�Vy5R�^�C_���p@��7�!0=��q�׫� �H���Ȑ&�-��\vER�4�7$���Ր��
� ө�4�\8�D!F+j�/�-֤J��lތ])�@Q���3M�S�|��K��)'�r��j^����lk��V�@L�SSq�ʹ4��@�he7dh�k^m��NAr|"*����~f��*K}L�8D(�hn
��;/|�g�Y�ܣ�*j����.Z�_���������/�}G�O����or����4�+�!�]N�e��#�]��{�{r�2��le�zۺ�~����c�3�
uAw��~<x�����>^����ǧ�0��K��<ݻ�|p�rA��G�֎۝�'�z�;�l�;�7}��7պ����Hj��R?�Z"�\�=kRj0߁˶m���*Һ�8~�������������g�����^�S��ކ�z�]=ٿ�8<�ԇW�߼�����ۻ�^�?ٻ��Iw8�nd�38{w�>�y�>l�~t{D�MNoOm���7�C��a+X[�����i�t8�xG|My��Ob�tL�+��5��@V�+W. ;klΟ��'R��fX�ِRl��s�^���#���@=f��D �����PԸ��y�6#C�qeU%�8VC.�m�h.2���=�_�Clu�ܹ�E��c�ʭ�^Id5!��\��:�T!�0����i�z9�8	W3W��YU��8p�����e��e�;�y�j��(�~�	�Kj^��J��.��q ����Ǌ咋-�2�&KH��kj�I�#�q��N=���h�0Lgĳ1y��#|�0����>�0d� l��m�zeL,5� &Ka�Z�Q��bhŚ�K�8����ʛ���C9�z!6�f[@6CE�q�R-���� A �Ym�jX�57��� K-BUms}sD�yi��Y����yK�a'NQz�v��"�i��`R\�'RI�Nd'��Qٶn�য��) [z��c�U��Ԫ�WS����z��j�Z DA�
��
A�,���J�Э���+PƢ���c�ު�K��������?����?���������w�}���/�O|��7�x���!��@#�C�����޻߽��^��|���d_��<�\�|}�D>��m?�*P��:��ێ�zj�5�Ԭ�
�kM�}p. �%me�.}��>`���4,){�B�!&��C,�m���JR%��h&�G�x'u:&�(#�!��^��@��%M�`d�h8�Y`k�B��Rm�(����	�X�A����/�c�#D��h���G������N�����OVO�>�´�ٞrd�Ǯ�^B|��?��?J�D¤F�٥0�Wj)�!N�jM�&o"N�fWID��ڄ$h��UXe`���2���1�)���DB�ah����WSa"��3�eK��+d:=�!kRh���ܰ��48Pm��4�B�P�4�˫�����nk�/��/z_�m����o�=����!�h����!�V7ow.��9��Í�UvU��M��?�'���!�j5YZ[ǂ�|��z<K�qT%�Z��J����|���ͅ���b�ꥃk�"oC6�����Za���B�FA/�+2;}4M�eLdz8Z�A��F-N�����`3�e�ö���jH��AҤ#��dR��7��k��}�Q^����mH;z����x���������jrc���f�����'OOΞ?�# �&N�{﻾f�گqy���E7G{g^������O��N�<{�m�^�Ő[�7���9�}���,H7�jʲ+E��fdvznv���hq(��R[�N�E�ŀ�Q�)� �2&k�#�S ��"ǩ'i
h��$�RզW���2�DA��@?N����pj��˒��zmk�:v^ $>�\4�a#dH$�/{L^��"�tS�@=W��'Z4���.J��hsu�F s^    IDATp�E���kb�F�m.����j[Л�V^^!U�7Ԫ���@�t"�)��a��Z:��D��U^T���<���)\�;�ô�����(����B������(�aX�jC����n���Z^C�DiS�p��z�)�^ �y!1(s�/{��V9/C����'ŀ�8����:}^��Y^
b�e�V6{w5�Ka�
����7~�BS��bB��r�aC2���/;W��]G�P��(^�@=�J:����(�~�q�¯j�a%5�����MG�OԊ��7�^8�Umʛƛ
���y��zQ��4�7����].)x��d�e�4CL��U�ɫف�*��u�-��0����Rl���Z!�|F�2����%�moT��\�V����kUذ��UC�@:��p������n�z
�V�z�Sa��l�N^�p�^l�z�qf)x;��K���(
ASO:i��� �y�b��hB��zټ�����0�Ì�4�a\)�e��-\�\+P�Ǆp)�-�f�E	I'}I�h�#��7��+}�f��j�V�I|rA��诬[�P�K� cG���ǯ���[Л�C� �R`d:=�a5�"G�׀f=E�&�q�'IgW�k��i�R(�ͫ�hJ-W�!$caSV��0�&�~��*����ZV���Mmt�([:�iNI`{,)�(�n������)��H�C�B�vfC=���*I�%��'dזKT!�j�Ol��!4d�K�2
D`4���1�W��G��0y�Ȫ����"]�ɲ��7!��S�ٹ� T�f@0�X�^kW�x� 8�B�;ݷ?-�:�>{����5��nP���\Q�Ĳ�mL�ng>|���_|��g�ݢ;Z���Z)�\cp+WjGz}�D��͝����/Y�(�g&?`y�Z��7땸��ٶ������!�}��������IJ���6�,���\� ��X_��S*�XɯɸӸ��Z^�#�Fٵ]����Lx�3�
z<>:6M3_�F�W�.�����~s��8e`�=��05�_\]��3��{wt������O������zuw�������Ǿ��}Qr�σ"�2@�s}��n����i֚;.�m�o�CGsE�<Ȩ���{.F�����A�ܩd�p�E���E��W��I�=���.Zz�oø��)\��Wm$Y �}��/��	�F �-$[_T3���+ӖE8c�5�e�C��i�g:��#U͢, ��@�i��O�d�Lh���ߚ~�p�%�e'Bm*��Α�6%5e��,V�,�u&R.F�c'U"�Yj��K���!��)��ID��5a��@�3�Q(������kL+J���a�h�R�iUI���IJ���ސ��&��X�hv��R��c��A3��!#P_vL͐���Ӳ�.��Ä?j��f(Wj�����&D+)�u�U=e,)Zmj0��>cY�
G�A�+��e!�o��:��Kj�x5��hl�͢�"���{ Bn@����)����n	�����0��F�*/DO*M���,�XK��-�|dp9�h�5wFws|��E{�>"��W,�s+�'麬�f*�v^���(YS2U���oE���*�1k�����`K��n^G�ӡ�e�\\�[�~.�v�������½+O���������;۽f] �6�k_${��۵|�����|�f=��zft���WoO��t����o����Ӡ�IO��ެϏ�6ڭ��ū��U�`�D�X [,~4��\@d�X��pl��m�kk�j�RZ�Y��d#ސ�\	V-�����B�B"[��FA/���qآ�*NxCx
3M|�Ijp��]Qt��Fk��mGq�Z����n����r�uw�)x|�������?���}�]�3�����.5k6M��lC���x
���������7�"�w�WW�!�ڨo/L8Gؤ/W[�����*��8�`S�&���P�,Pc gw�! �Z�m�:l�\�C�A�W�a�!�!��J� �V�\p�D��Ն�8;�2���F�:X��[�!�xԳ��,���DdqD����-;�W1�\&���p'���������{G�c%��Գ��4�Gjj=Щ�MS޲P�88��F^ۆ�����t�
Q�^�V��-#C��-��;^������AoM&J
�Zv�j6�Y�[.Cs���chR��H��R��$on����e`���M�Nur	ߵ	
��%�6ɺ���T�6�7�^���^߮;��+:�������b��u<�ە�>�i;�]{5twqwu|pzyq����9^��?��u����_��{;���Յm�i�7}��g�/~��/�ۗ�w�'�'���a�Qa�B�*lY2ୡ��e5�V��=���M�fȋi(�J��9y������G?����O>�Ē�i鈲υ�TC���B4.��o����A��l!�M~���9�!j�Jyi�B�2UEK�����å����fe
�x����X.Q!�L��M����lv�ݪ&��\bEi:��Εr����Ǩ �"�/o���C�'�Re�z� ��I��jtx�2��'��`F�>j��b8��(�9�[��(g��0�h�]O�W�����\ }�#�$j�a�������7��4�dG�i+/Pje�I��q��E��cq+R0.�"�#�f��G�8DxC��\Djp`x��	���!��H��g'����S�>���B���>o:B(�1���V��̂�P���a.zR��a�I�ϕr`� �=�V�F��p=A�����xkl>�^
}�	F��H����=>q�R˕���ު�g!D��T��\)WjS>8�'2H˘����oؼ�6s�)��y���/��y��2��b�I!VjL�l�&$�!�(pɂ�6�R��A��h�SҤ�hbR.����y�pd�X�*5�!����V���P�㎣�C��zd.��2�V�+cp���e�Ό���G6��#�ҁ�E�!�ֲ�1���K�ߐl�$6{Vɐ�>5�j�@�Z^"�dD�k�O8�l���:U!p4���?A�![�������ar�=�b�q����W�6��@4S�˒�L��^���)�*E��M6$�I�,B���!2��d�4/LvCH�4̪BI�v���W���Bz�"��)��P�&��8ç/
���1Ħ�5�Ȇhp=�T6�J�8b'
	Gne��\E�i8��H*32�}؂�N�V�NS�楜w6���VLG�fjRӦr����a)$�ARS'�RS�/I~!bSơ6!�b���B:S�"�����J��e�vKm}�q����zk�}��z�+`o�^_���؈�f�9��~_���#�3x�a�Rv��{����Bׇ���=��i+�G�	�ʹ�|�c�����a���W�{��룖�G�O�.���nj�z����Z�2;><;޻�~�j��<Y_B�>
�&ޝA5�N�c��m�n�n�j��fe;���o���&�E���=�R���N�;������sS��W7ڽ����g�e�����GE���^<;�8?zy����;x8���)�;_�6��J��O?]c������}֩{���w{��{�M��ء_���2L �kh����$�i�0����p��A�u'L�0���J��JW;Ӌ�.����N�a2r�5j�l�q���ՠ�8z|-Z�-hM_X��V�&�`X�'���@�a20!��� >��j�+up'N7��V���'%��mh"��r(�.�u"��geHg��C� 4��G��#�+�tx�R�����/�d(�ݤ$�1�P�b������W�D�T<>q:�Px��4�h�-zul�K!�Xd�l;�d1q+_�C}Ey\ՠG(E���6W}LvU�bN��DR��g�g=ټ�ě�M�BRh��)�$(�ƕtd]jƤ�d��Z+^�&�:�j��Mk8������-iC�1�,��e#��,�g�	V[L�"�\�ؓ�N6)p:R��(��ЙEAv!MC��t8��L�++�5v�]=�I�&>��In�P�b����|��+A�*�R݄�Z����Z3i¼| #�E1�;��큛��l<�i�)��������j���������/~����J�����V�{ ��s���۷\l'����˛���sw���Ƭ�Z6��e�K�rW�6S�z��&��c���{e�|��J��	124�sh�Dx�5v"�mV%%�5�j�M��� ��,�m�Ŧ6�++X�Q��'HͰi�6$�5�����ˎS ;5C��M�͙&Xm�B0)�۫��\�w�mn!�Eq�����v��a�bj����ќ<�l��I��Ŗ���'�j롄�e«�׻� �A'K0M�VmS�#۞�*��7q=���bGP��j�h�5f^�(��L5 $�4�l=1Ճl��Y�&�0qx� \��zL�@�"0�(æ#а&Ys���A����ټ��{зt����4&�(�9�-�OaZ�?�P�j!hH�IA�[U�g��o?p��OUC<>z߇�-��g����q'՛����V[�ح&)eHJA8/�Ts�裏
�7#6����a�T�(H��\�da+���<���p�aF|C�F�]����Za
-fQ�V`)�ՉG���a�_�U`��M�
��ɀ��mq�F�U��A�7�����>����M6�^h!�[G^�Y~�ӳ^����B��L�9��q{���g}�?�D�\���<;z8{r���/�>��7��_������<�x�}~�~�UI�
����Z�to���Ҵ?y���V�45!��J���0���oH�m�R���b?�v�a���H�証,UeXAdI���(��\�z:R���ɋV"�!��l}��آƩ/<�p�:U�[��92R(*e�����&Ȇk�z�i!����pQZ��V	~C4��z�6�Wʭ���$*�!Q�a�b �JM8����N�S<Z��Fӧ�!���OGTv���gH-(Ml�0�7f`xC��Q��\ۂ~W�F.��k����!�R���6����E*W����a�:�9��D�7�y���]|��G}-�p)*CxO�J��6b�/W+/��L�ώL32sd�R�Ԙ8�0�R3�5�@�� A�ʅ�T�G�.ܐ-���4j�Z���M����
�� 6�-�U�Ξ�N�k|QSy���eDkj���79�>tpE��d��F�rF���ג�Z|}ü�%�߁�e�xs��2���^R���7Y��s��>���dWC���e#h�_υ��̐Q8MFd��88��fTOjB���	̈<1�_l����1Z=�)xȘ�Rk˱S�A��NQ��Sƙ��j
�8lm������ѯ$ò�ِZ�u��bv~aαc#�N�����ڊz�t3:��i�.���'��
�5���Y�[L�F�m�%�`846����,��©!h�DK�+Av� 8)$>=qm�K3��4,�!C���в�Sg��D����L`�/ō�75��$�,8�B�̠lU�U�6�Uy�C'�8�Z�E2���h���VL�Ē�%�����aʫ�b���ݛ��m0"�D�@�0D��b�V�o��W���(���U�,�����0����7k�x�pLF� #Ul�]2���JS����;�8z��X��XC!�3�b[.�kA.uU�u�dg8
�j�o��QI��q�����_Ϧ/��X4�ɦ�!��4�I��7�������u�E`��I�t�: ���$��@�,�����R��:�󝫾[�������mB��Oxn��ޤ�z��|�pY���k7�V��}������z}��vSt�o"�+����������3����޳gO^���>�����S_�*ˉ�?z�k�>�is��?��9׊��O�:-���Y�Ǐ�����>}��U��Ϫ�Qo��ܿ<;�^��K��;���/��\n{�y�:�?ݿr{�}���ç�_�sruqy|q�xw�����{�;=��q�y�,�Yu�p�n�MЃ����WNo|:�~�f�~i)�C��_3���u��k.��	�vK����\yw.���y���?zH���.C�&W)xql�k����j�F�oHS!Y��v�6�suh8�J�0V�֐C2*�]k�h8.�d�M�H+��z3�l�_�&P�l�I�8㊟}��D#���@�8D+LDyN�t���i��8B)\�A��UB�NR\h��,~5+Cv�
��5Q�s(��q֋u4U��Q�x��Aa��o.���!���؊44��³��Ua�a�TU�(��Ԉ�xe^VO�>��G���%��S��,K�S ���p}"(,)������)D��&��0ጊa[�&���"���AK��Q?A=CC���j�:����l��n� ��g�UFvyK���7�l4ז��֜,��HU<��r"V���(�^��@�fs��D���R�ӯ�AxÒ�������.�a\�w-��b<���p�s[YT/1�5}��gJ���jU�Z+�"���[ޚ�"�iA���Jc�%�l�.R�4sS���}�������j芭�� ����?���m!p�@�aR�IӬ����pg��P )���[Ma�$�ۚ̐af��5�r��(}"z
\�µ2B��z�@=<�J2d�0#~�Q`�Y.�c�l�SL~�Vm�C_K8��($���!��u����9N3���ve�������駟����n+&�]%�����ɟxC�p^ǷO[
4/}|��8A�c�W��Q���~&��+�Ie�)P֔�M���i:lC;BDI���k33 ����*�T�^Bz2+����˥ɨ�NIe/�MU8\&D�H�ӄ�Ue��f
/�!����5�#��X����,2��x��#Td!h����);���#�.GJ�)x����#��`ҫ�Ԏ>}5Xv�|���t�4CӦ�)P~���4���i�?��[y5��/���SH�@��YS`$�c�)��#EY��s	1;�~c���p�&�@p �sA2I�YFk� ��ަ-W���M�������Y���u�y�l6ə�%g��I6�I'@`8A��?ȫ 	$�ۉ<cٲw�Xl֖F3������%+�q�8���SO�9��&�w�,D��9�|�ֈ�`ʄ��jFT��@N�Nc�ߝm��n��k�E�Z�=��cS�����v�O��� ������� �S{��S�������8-D^���H���7�<��϶��1ֿ�)�v���f�ZZW�PH�d�+*4�|8�n������3W%���3>Y-��S��m��)H���H�uBM9�L�L�I��[�ĤN9|#>�"�FM-�!��+��PLS���ɯ��|Lc�B)���@6��J�T��������89moLH����(K������������V�H
�M
����n�I��k��/1�Ӗ L�N4SF�Be6R��ʑB�д����b�$�g8�FQ4~����)��\�-0)���Q��G:��U��8U�D����示�������"�tN~�*�x�z���&5˩C#�h�iE�(�`�J��D{):L8C��j�����Mm�"�t`���D�9|U�s"鈖kZ�Q�^m�|�̦�M�iQ�Uķ��/�,L>�\f���x�D�D0݈��4먨?�lf�@x̺J-�Hj)�����`ĉ�xkI�-�Ĵ�A���V�L8㧟�)��SK���7���i/��1<���ɉ�.g*�B����72Q�m��3B>}�齉<E�T?��
�S!�m�t����	�ЩnHӉ*Q�6n��[]�����Ԙ����1�ҙ��CjL�,��F�e�e��ѩbjS(�TVw+����YE�RN���Tj5VWJN"��|j�bl-�iJ���'�D<>+ͅ�@�(΄8+�g])%�bQ�?`;��	�X��|&�䷙������]:\E�r͘r��f�U�Ҙ\`%�OEL%���J|�~�|R�@� �!_�B�|��«5j�̔�eDn�6\24�	�#X�h����?�t>Ñ8�    IDAT�"�������4�&%B�1YNY�US��m];��岢�rb�c��$�^^�j������
����ҟ.���i?p��1Ncu�a0�i������t�8��L9�Ɋⴐr19.%�0�A�l�Y�B���t�;2j�NR9����m'r�jA[���l�����������#���4}�����Z�D��(�t�����s�:<��oz}����^���f^�����Ww7o�����햨�R��!��؏�_�=<\?ܞ��m�v�X����mg�灎��bۆ�r[��룮�%����x�ٿM��3/.��1��gϽm���n��K���߫o?��TQOx�%$�u(������7׻�.v�8��ϟ�=|}�?;�s~������S��y���*�w�ޯ��G����e��Sg�v�ש�[�MoV�[�\A'�k-�du5%r�LAH�ڷ�7��Y����>w�{�B���0/�~���߯C0�z���!BL-��)�So�s�����p���o]B(%�!�?��\�ĲB����!����}��xF �~�w<���V�t�$��]>��Ff���~�Y#�u�IS4�)�e� Ϗ3J��p���zڗ���ײ�Fʦ�4�B@WX]���A*��\V��N gn
�n�p�Vo@���� u�$�R%�Lq�b]��6�{L���K)wq���R.ZE�ݣ�k,}���P&
ls ��!m�� �r����p�('�n��B9�����LP��y�N8�ē��B��W�H�)���F�w����l
6jv _��8.���"dW��[:��@�p4�/��G
��Ȅ\b#}dƇ�bzVK֦���){|�=����B�x�W|G��D7��5�`�S&����Ͻz(h���9s�˔3-v@���Մ(�+��j|S��i7�}ɏr�k��Qc|F�r�~|PO����g�z����j{��ɖ�|��YZ�k��B4:m7M�ê-��O�i�kY�X�`�dLNE�4��!0H����9tLS�`�D0��(?Z�D=���1�(p�fѦ!J�i��K11�� �4+gB6G�6�B��blRB�P{h�ZC.]�6����_|�
:{)�9þ\�ٟ��g�}�x���]V�+
��*M����׀/��ap$^�zE��-���.�k����rƚ�@:ݐd�
1���7*�*��ZHQ �Q�MHS.5F��PSk��*aE��UD��P�b�ᦘ�"ޢ ��	�YU(�L��R+�楰��*j��o���p7����Gn߄�	|)�_QR��ԡK�V���f�[�D�?ֿN�M���᫦�Z�kɽ��Hͨ�[ї_~٥�橤�ltb��� s���%xU�$xr�0H�%*E>q�i�sJ�p�j��Y�~Z]Rm�}���*�b��/�Xu)@�)�9Y��9҅��	4
A�4-�+$��TI�慖�YoM�C��C�V�A��B@SY�&���i\e�Z�v�a�d⮔%`��J�0Qx�G��6�OW��Y����"~�-���?�Ͽ��3�u+�_�����Wg�e`ך X'�]��t4c�4D�'Ӌ��ʍ߆�9@F<M�&
Lͱ����(T��*�с+�#N��B��i��8�YL�_ϭ�Z��.%���IG�S����/ί+SQ4!05cm�Y���@��/]t
��L�f�,���*��iz�8E�Ҕk��������e�1�RM!B	�4��R�C$�>�+E���9����DS4#��	�IGK�0�,�Dp� 8YF
����K��d�UL�\#�Q�gmQją�5Som�Q]֭!�2�G.?A�h>Ǣ"�����'ȯ��ri*�z݊�^���BˉIMH?�
1�)�1����!�~%D!���rj��jU-�V=4N���I9�Z)o�W�h���)U�}WL~=�wAH���Ⱥ��F ��F!]EH8
N�A v� ��o���l6M�T�B�������6����h�(ߘ?͠�KԳ6B�ŏPc�ȪJ:��j��J�;-�z�PzU�ATiK�kD:5�B��io���U��YV���4M�hE���P�J�@��ш#�����)�moߺ�]�%��,�L
�S-c�z�c�/ez�G0�I~F�'%�>���F�i�$��	�}W`8�ߨ֔�K7n���O��� �)�.}x�F�1F���D�&�;�/j��JG?�75����J-�'�S�4��;���ۢB+�Qb�Z-�ňUJ���h�Yj��MĦ�GQ[��������|�������:�u?#��O܌K�	|s��0�P�������@�9o�ݼM��0Wkq��(疺ѿ�J�����$J�N�$L��O�:2�a�%>��k���m��5JH��
C���[�B׫/(��5|0��p�1��\rE�h��~M���v9��B4M�(@H�͜7�ԟ��ߨs�sT��p C᠍a^u�6���S�z#`u"B�H�吻4���|�՞qϖq�e��u�E	��
c�ٔ�����T�'L�AZ~��R��6k��[�y�#'9!85�/Zzҭ��@��TPQs����W���X�o}r��N=�ﶦ�6�<1������ak-+u3��4�=Oik�zqv����<$�߼�r�]��=T�����㲾H���-�45y\����Q^��$���P�9���7����0h �^��c;��D�������[���?s���,N/^N��Qi>>Z1��v��Ϝ>�%��l��`�4A�DozcP���5��6��Qur ��l��d]�̐y������S��؈��|x�,f=rs�5��T~�Tb|�r��\�現l�_C���M�g��n9GOcS�IK�l�j�D�?��0��:���8s=R���i2��T�kN-\J*\�W��/��O
�H�0�=K�]Jg��͔��i�} ]ixӚ����+�̩�h<߸���m�@�Ђ}᝝|��,6�|D9��m���~F��I�:�pOh���?ɦ��~Dq�V�EK�?��	򻈘����vk�Q5�''&�̝��X{�{U�o{k*:��i@F�K\ilS3L�
��ixbʈX�Q�� ����	J���(�#�Mx%r�ff��If]ҫ�����gɼ��#4��QV�}�c?�yo����)$W Ʊ<Q�5?ʚ�ɔ�z_�����I��W]|�����]��=���.��\hrQ��������Y�Y����V-�@2�k�������Q��}u�3M<��g�R@[�«�Xl��>��TҤU%@�@�h�X-�}n^5k�*%���\;7%�58z��X�q�UH�YT�M;�O?{�\��T������NR�σ�$�"�o�vE��}� _���%ߣ�]�mxX�D�o��)3�6#��d�DN�u&�Q/<qbbn����s�xX�6��=��8�����"�s=Z���p�5���]��f6VS*�)Z��2�֖�C�� \4O��k�(���%>�X��ϐ3�	#�"1�~4)左,��e�_����(�e3]Kд���Y�{Ӣ������?5ʚ�_n�8�yku�n$j,�Iw�)5c���h?W�E\Y���qa�U����e���Owi,a�T�N���B?Jp`QRZ{��y���" ��'���}���L��'jھ?ũ��U�Ƙr��f��^� �95�rp���隋�xa�u�R8���gFC��8��V�gv���~^eq�!��Qi���d�(�qXݸd{�������L��H�*�d"v�g�ko�mv�f]����sA���ſ�t��f� ��a=E���u<O{�%�A3�ki��1C�����VI���ga�~�ǁ%t;/"�� �I�6k�EP��R G/����}�HQ挟Iuj�[J�a���n鑈hD��ׂލ�i����$Iխ�7fz4SXې���֕<��
��������v��'�
Nȋ�2����Ͼi�T6@\�����u@pfL{�������8���"����rYw��L`cR�X�;RM$N�Q��3��4�\$�@<�d�(�|�����b���΋* #��:&��@e��RԪ�n���T�%��A�>E*�z�����|��]_��]�ifMk�N�hW�na�NN����X������ ��h
��/٣�Z
 �ߨY� 5�P�F�sxXGQnZa�p!�����M�<)E;vU��� G�.�@������	$h#y,)�ְ��m���8w�6�5�$|���i2exk��`��w�c&�V�b�	�#m #Kֈ�gc�~���U	nUQ�*a26�ZË
F@��S>�g*Է��"+x,p`� �(G�x1g��[8���n�B	����ϸ���K"�j�W]CR���@kx"[���T���n��tցJ����)l��*_�r���;?7!�"ɱ:"�{#;Ha�~�A�҃V�X-P����>���es��:�a��^���S�:[=[������X�*5��s�D��`�WTI���yj�|19�U?�>'X�	�u�[6V�rd�_����&lyߌ������i�S%�	����ą'啵7�:���d\�]���C����h%�`��S�5
��;�4M����R~8�M�H#B8�Z��x&=Ȧ�/�q�۔�x&mO��U��뛌�]��o���r�cb���&}C�o=�*��eu�'���D�4p�j.Í$�G1<:{�CB.ê�I	���@``��31�y��딓P/q]���o�t=D�H�������ȼ��2p|�<�q �!�ɷ�d���}2GkR�v+k��P0�J����ݠ���oW�y���]Ԕ�pj�i���X"���*2��n��Y�J��`.��
��kx���^_����|N�\��[���C�E	 �������qȉh��	Ԑ4��#R.�Mlz�˦��x4��G`+£�% >m��?Un�j���y�F��jIԻ�%��ԏ<U�QRm6S�PÓ�3���O�4䲋�N_{E�
6�|���ngo�;��}�����]u��7����/};喾�3�bRT�Ks󳪢I����������+�&�uGc�i�?T�lͪ������.��ӗ/Md2}�vQi��"��f��1w�sU뗊�#/[��?�//��وܼMstǌa�����_~�yy�l�{�ۢ����e�u�7q �������b\�9q@��_J��'׻�nm�jfﴚ]J�q������ׯόF�^{���L�I��`����&G����w7%>�]l����8o&=9�����h	�mg|1��B���BQ�ek<4,I�[����]G۸
�ۊZ�"�κ�OE��/����x��0)6�r�B���?'�0�Hj�%��?�72���O��!�\�+@��-��K="0���X����׃��ܝg	��U��"Py���!�C}�>�R�R�L����OQ�n��4������O�������#�<7p�J;���Y�������,e��8�s��#ɚ��S�&S�p18���0�(75	�?��o���Cp6;9��WW ؃p��J�� ��FR=+����26s~T��~��`�j�xv���CI�,ݜ(��-�pW�*J|E��<�8���C�;3��%�4��Wq,��z�cKJ�����I$�.}��;�L������"�A3�ɿ\s�p��̛��c;R��rӺ�*ƩH~ܳH�>Ló�K�#��ޖ��-@"�yVׇ݌|P~vHp���;����k�bt�3'�{���g}l���Dދ����R�ٍU48����z��we��꼇0�z]�|��9�x#�����]�	��d�N�!��y�+���'{Қ�!/S˰{"Y�ȱ��C��g ҂�%a�4���Z�վPJh��^h\�ˊ�ދ�yeB��ũ�9�v����Q��]SF��F`���{ﵟv���$<��ȅ�K-S9q���n�9R�"Ls߼��ş���B�i}�x�:[����m���`\��SդZ�<���]�WN�R-]V�S-&���\Q,gzq��/����X��
M)�I&M(^A�N`�Q���<�Y��Y���h��b!�\�d��0�}FQj��$G���PN(�zt�~\���7�m�Yy�s1���Y��aar�v���C�W�P��*��Ob���ʐ���H��"��� 3mۜ�>���켐�`޳�E�������B0sm�G+	LOo���(V������Ћ-��Vs���u�����;�O/ݧ��ia���nA�/�v��j��v��B�������f >u�ɝYz�ө��d"�1������G���U��k���[��#Y�@MX��$+��S�4�%���\0G85��6]�(
 ����&?j+�J=�Z�9�ؤt�X��t5kR-�OD�����r�zfT<sD^�vJ(��m�����\�p�G��'��˰�Qm��^��!�$@��)D�?!U��Vyɱ�T#
��r��
u���
�o�ch�n�r��u(�Km�d���;��B��.�rE�Z2��˙#<�q�^�����b��'8�6��:�`���fu�o��>��]P�-2�`l%��%4��ɝ۬�b�irք(��iά2��-d��d9Y��gށ���S����N����v�Ϡ<=��ʡ�x/��ҷ�.
�/��:Y���]�R��z�{��D���7�4C�0���$P1��R����[*�rG�jV��I�(7;6}�^���C�8�1�˲q],᪎j�G��X���P�u��`�W�Q��[>��~��){��~F�{���Q�q�r�v�rh�J�1t�MlS�҆w���;��_��bcO�ʞ����/md'��ԑi�Y��x^	���z2y�T(<i 2�V���
�E�(*k.��ֿ���;F������<0c)�(�>ȏ�
�@���Os������A+�q2���~�z&#!٧VCu��9�~�ĤO��*ځ��h;&�֗�"I���vt��8���<����L�o`��]y6���M�C�]��p:�րMU7 | �~?81�u�"ȌOKR��U�.q�x_0�6��LE�cYf
&x��\]�&bB'+6m%��5Q�B&�Q:z�D)��0`�����ah���0��11�,��g*u���},tݜ��t��(n�4QF��#�%�
[��n65-�)^��5�Ѡ���s�.c���2B� 附�`��95���d�'�pxY�zXEԋ^3��2�$A�ѹ��J��"|]��C����h��ĺ�X�A��B��=����h<�/���e\'��P5�8�\R�xS�o]�����Eyy���L����)���u����L�Cڑ�?��u��A�^��]�� ڣ͟��w������D�y��K�_�c�G�#�����W���7G�rZ��o�5d{�ܳ;�ZB�׎�>j�?�T��4��#�����~9��w�*�.����! P���I�TO.�d6���_a܏��ĭ�����]w\���e�
om�]E�~jI<��Z���F�mr�������N��춯�;�5�Vc�6F}7��fs4��o�Y*O�nƅ�5Ħ����7��4�&x4�B�:�~\�*�g�h�����)�\h����D֖�=�O��L<Y&�'���C���Lg�l�Q�ğB��5�%kƶ˲<V$zT�2��	-2f�]��Z�ϫ�o[��(\+~����us��cʣE,L|�i�g�j�,�OU�c �	�*z�v�-��r)��ę���LHg�)S��	Q�j-��,aҙ���}��c�p|j���^��1��u
�u�n�l��c.<�LWc�a��t��&��KŀEʱ�~�Z�y�@R��j��d������Þ��~�˦��+���'��f�{5���������S��`�a��RBF��Q����3������/�����A�[�R�K�&Ŀ�Aгj/�_���F�?�`&I�`�B���q�mI .�}�z�61.�j�΃ۣ5�
�ݒ����.��>U��'HBU+��wuO�Jc���'���t��E}�e�5��䛤���m4�4�"c;�KGB˭� ��rl�^z.i]�L�iɽ�z+�jT�gi����i���y!�<]��!&�6��~����0ω���a%3����,��3/RQfn��ʲ�/�#��ȷ�*2a5sI_�U����ȇ��	M�� I��g�`x���$V�����e�^{���%zPǌY�Zb�c�yx�)�T8����z���0^�,��I4�8AN���ڛ��4 <M��!��o���Y�?q��Q`WL��(���M�~6��W��8O��s�D�����e���.�8�gy�ĮI�d�n���߮M��c4ж�
g���5q�]�~6��)T!�a~��SpOY�)R.穼 ���W�G�Hz�5+%���}�!�YQ����̭4��-a0�Âl�3k�b_����ߏz�t�)�L�V���E����&������9;���'�3]0'��
�LZs��$P�Q�wG��>���;��LHT4�
�8L�(!H�}5�6��:�[Uӛ��UOxUa�����*���jg�u?w���=�~T��	���(q��\�͞cY ��R&�m�� ��I��!A�_#�p�L�ѷ�?x;��(�?�2&��]^�M�{�7��3���8��vй����ՐP����^%߿&fDMx�c �E�;��
�(�݄����ϧ�@^�'�׉Pl�<�GX��M��	̥E/�X�b[V��3ۊ�bh�~�]����F�C�={��{e�6�y�XK?퀇ɩ7��̽;�Çgٯyj��!���-N�1SC�q��t�����
�b�O�Q�0�i�g�,�}^�������+��(�$6�����|�6#i�[���30`�ap���S;D~.G��:}�G�o�v�ǓC��S�W�*�P�Q�6����(�y��*6�J;��Wq���z��#l��"�R|�Sz�jܖ����9��b`����/�8l.��S�I�dݝbe
�%?VgLeP,��?��.�cm�P0��R���ߘ
P	��50�����	k����o޳�V%~&�0�1�5e�a�t)e�)8� $�Ӽ��jHT=F3�<5T�C|�kĦ�X�#,�zxr�q�[��i�$l�q&l�rj��b��vM��;]8���.�|���E.[qYAI$�����ިK��\�V�F2~�v��,(p�ꄃÐ��1p����Bk�q�S��@��>�*1�+�������!N�����d��|*ܛn��_�P��ʣ6A��ꓰl��A�܏Y6��~2K4bQ�=�j��L�7����u�b�/�T��}��h���c��OX�Ͻ�aUF�N�r>�,�׼%-��Xj��
��h}�����p�k�^�ƒ���ػ4� @^b�bQ�y�A"��#��� "����b��|�k��c�"��%�ĳ`>�G@x���gU���7�ŋq��A4�������&y�FC�k�e�sEN��q�)I�Wڕ�@�y�����[����dSk� �S�9臊��;�~�����9�r��L9�;b�r�<]�]St��;Y�4���U�ꛈ����lZ��p���I�-k\6b ��eC�3ԧ����E�k/�j�ֿ����)#�;ܣ��������ɑF��o&�r���,�F�!������i�	R�n���^�,����%v˂�
T�6M���wOe��J�K�\���$/}��7�eH����ݻ!�	�f�p0L�/���ϵ��y��m�ɻ��ݵ��?���g$o4�?�e�/I�,u,�הp��fG=:�8X-J�^�:���n��uz�jql�����N|�Y��R���K�����qK
d�u�0��V\��$�����՟�f��&�w���N���F�K~]V�w7�FU8��|��\�^[lh>��c>X�=m����;�@���<p����[�;���`���lR�l�ޡI�L�����y"�T��ǿt�3��UN�8��{��� Q@Y/�Q�	�Cߑ�K�����љ�x?�(˫b�f�3FU��4Ą��E��r��q$]#q���n��,�"
k=ٺ@�(��b�k#�h�tD]b%�v��_���j�	����u�$m-�P�ۅ��u�&R�)�4ւ�ȑ#KڀX����X$��[���o�(���<�Qx�f��)Y.�s��ea��j싦6�h-�;�ه���m�M�UM�������::=�5�/�/�93Ү�u�l1MM��+��*�%t�Kha���^G+k�6Ymhڸb��t�����@���*j�W'T�V��+H�	���	V��3���c��S�[<�k���D~S�o�7�ނ�{9vy�$�-ء�HADGŞ�B�T��ǟ ���t)�%!EOե(Ѝ ��C&��V��E�'�|��|O��"�Z������8�R9��c��/��j �2�Ɩ�?�C���w@x����fsm�ߧ�j��M�]R��%�� ����{�7T�����1p;�q�C�W^�'}�9�]v%�� �����ZD8�spZa�F�����Y4�.��`۪��Ed����>��R[��ݘ9W���m�!J�Ҡ�vh}^�\��G���dgP=I����5K*♷y�g����՛�>�1�c[�����e:˖\ԏkD��������>啯�gE|1�Y��⯙�;їq"/6�.od��k��ŉ��g��k��)����l�T�L�	I.>U1��G� �:=��Km�U�sE�^��P?���*���?�'ܹp�NR�}����җna���s�j��?n�4�!/x����V��d�Q�l�9,f�i��Re�g�E�鏅?f��ފ���K}r��}ӕ������������܋�Υ��š}�7L��V^��ۿ&4
�&:��(<�p��Dw����sRP��+,|�HtQ�_�����s�E���b�Ѫ�{�Vĩ�[�)�2\mN���M�2���	{A��hu	?p�7��ǃ��	4f��*����cW_Bz���\�[���~ʼ�8m���վ:�t�/X$М��B?�t.V%�q4�p��J�唙����Qa"]=���#N��R�岹�������'�D,D�m����ru�IT�}X��D.���U�ĉ==C���/l�)*����)��jjH����v��)�`�>�n� nS�'��c	�.n��L�!Ŭo_�RJTbz�h��Jxr�I0hU�Fe�K/!H4}z�����x4�P��e����������<Y���� oHr���k��*��RH��]"����0Tah��d�'�Ӑ�0�D�K ����D���zA���ay��
O�h�&���K-�)$�t���;�ﮣ�YG�Aq@$7��@���`����v�m$�у��L~���e:N�J��� �V��P!@ɭmt�X���_p��y�k�x�~��A�n��(0��<]V�%X/9A#��d��	+�=k���ЀJ��Hj�k�u�0я��ӷBr�t�ZV�_�a�9@yn,q%:��d���(4 �2R�2ͫ���xp�I�����M#��Z��¿ ��V:T����J��y���L#?K[�}����c���_�Q����lB�c+��i%Zr��Ÿ%H��_.��E	#�I�78��z+2��WPQ�	��+�ZL� z�C5�٢J��F~�iҿ7��a	]����-��"�TҬBV�w ��OMci�V�����5hj9s%2��Xe���;[W�B��z]�EwP\�\�Z2w�s��ʮ��#�(o��4Oj�SRO~h]���	"l,~�P� A��N[\u���0����#?��9>�C1�I`p2�E�}W6���bӖЁ������	V#*��Eu$W�T2�{��Y��G�c`�lowyv�z*���ھ���É�|��=��AU*#t���������l������̆�t�T�����?�
�`�+mvؕ�;�T~/�&^�t�� I�6�p�w���F�~���8S������Sv�!��ȇ���6t��w��G[�Rřȱqt�=�DO�v��84�;h���?XP��fC�c0����Zu�Nתq�ts�]��M~W]Βm@m����J�s���+�������gy��[����x)#ҭ3�!�5��,�Ճ_T��d������9Og��o�ߎ%�e>�m}�N7�Դf���<��ɟ���՟�W�;o����-����w���k��Kً��b�魶��"�]�X�4Lѿ��;M8��?s���� #�?�.u\�r{�cq\H�����z�t44�?U��oY|��_dfv�zq�Q���ZV]ʲ�� _�������-��6�ƙ-s~��~m��f���D_����	����~n�#|]�ۖ�d(x=\�oH�m�O�E`>Th�$�ix����>px��i�Z]����p0v��rv<]�6&��T��:��l;���0���;O���o�����/�P�+F�{"����4t�R��8�I��c��xU�@]��*�y���/����y�m�n7��_m�:D��&�Ʀ�yx:��(#���P�fL�e�[�ŋ�SHE(��Kc��Yِ�
]��9M�I�/�ghLLcN���t��d�l+5LR�@I�eK-�L��Az����Bo���S�q�7L�o]�`�������<'W�:8e���rdsew���<�Y�rfȬ�/�9��e��O�R����I�=B� bN���W#~
4ϛ#˓�DM}��;\�uYyRI�{���+QxG4�����)+�)�
o=�ۨHQM�[���}�Җ4�$Ʈ NA��&�2��`K]�F)g����&Q�����&0��X�Zt��m���tF\�,����Ꮕ)/�ޕH�}���џ���$;��J�ھ��s��t��T�Jp�nO�а���u,��%�Z��>�����<Z;�TX�1p�4�(��8������@�����Za�qѪ��q��ZC:���E���-$W����+� �ǡe٫�� �����m�T� ��KO݇ۓIQl���
j/z,���x�Q��I���nS�n
z�Յ��v�"�{����ҟ8�I�����Ǌ^R{>ƎƅŶ�x5f1�����C�����[�9�����r���^��w��K|������8%zخ5Y�0LRӆ���k�]����je��6~J�(�`�w��[�0N���e�)ݏa��#����ܭNF��h`�-C��jU:��Ɋ��L�fF5��ҷu9��R������wm�k��z�n��'���N���o ���4y뭵#���#��g�o����R�[��֋k�u�ɆOb�Sa�������K��ޢ؂����%���"��� �"�)��%����t´���N��H�
�6�cV$�;����`W�yHv��I�������8�V���=��e�.��ϧ!&��N�2�n���
w>�9�	�bmw$*��L ��e��9zۜg��Z�ޫ���!`	����\`�B��C�����K��͵�UIFiP}R�&�r)4��NW'4��Z��c�1�7]���:�U�v��/�H@	"u ������!
7"�H����l�r1��1tz���E'��.�>�4<�'I��g/�M��'(�wغIr�h�1�P��������fXi���h�/jҵ���Ā�1�Y�-�kA�б�yJ�qP�H+O[Sf�Zi�	�Г���Qʒm>	/����`�U`*%����P;a�����z#YC��\�ho�VYt���p���/��n�F�H&��"�[0;����0�i��ʠ�>� Z�y,�St�C�{�?0T�k��h������Y��I@�|!�vor�!kU:/)Z�<�S�d��Q�N	��jP�qɽ��|E|��'��i?87ͬ��[�H��
F��b��6Œ�u�m$~�`�&����'���dC�1 ��`C^#Jn�%�n��z���x"sN�hS���p�]�=ǣ!��@)s�ն�(C� ��	{��&�a*�}t� C��*�q�F�O�~�Ս�F��T����$G��V�Y���Č�z���4VU�v�Aiwq2hb�)Q�]��Z'!Ư�M&c Q�"TL��]H՝Ļ�0�S2���v�PR �9��!��bW��1�����ro+ɯ��ە�pڱϞ)j�+ٸ
�H�:CR�%M!Pz�b�5[<-�3��QWE��y��t^KO�n�7�oS!~��B\WhǙ�~%�F��{?HYJq�fW4�#{:�Ճ-?;��	.ءg���(	�����!}��T�7�qt?��P\o��0�+!���۩�����5�t5O3'�O�;��ο/�<���`5>6T��I�{�l2듍��ΰ��5����v�O~�5xL���!G�TJGiZ��c�k$z�x�,g8A�4�/F�����k�u�ܪ͒����5��=g�e�k��=墙��v��]G����d�'��B�����)ϓ���#�h#M��a=����Lwg���"��P6�n���s뽯������6�OƟk\ϐ��-U�%w�Ȟ~N:^�M3a�}W?Yy+���w��L�+��{I�ݤ�*z�Ge���S~�շ��ѷJlc�̗͆S��t�����ӡ?�� ���f��[�s� ����6�����6�\.7���knl��3�����<C�����\��|g����e�R�\��7�����pGS��9�o����Qy�~G;�=�)��7A��F3���j*�Yt����o�o=s��v
�(��\N��^fZ��S����Z �^���>?�Օ9u���1���V'w�lj:��o��DyA��<u@���4wp�ժ����yH����:x����	�/V�Ui�v��9�f�LutX(�!2�9�܃�-��ǔd�{+��x*Y|j 	��)=w��#b�O]���zc+kL�f!��a�zqo�	�+�P���a2	P�h0�zϿ�@M
�8�^��~��,-j��o��R� ��p��6=[1H�b�<�I/�>TE$�O��U]�XN�N��/�,=�/dV'����^��%,�&�;�F��zR�H
J�xڸ��;��t4e�/�a�6���fdC�b�g'V��:$� ��Y:��s����KIX�%̖��ylV�h>�
E��U��cm��v$xiU���(���$_����+�nJV藮	�<�k���P�`����Z�+�e۞xqi�ju*�XԱ��X[���g/P�|��I���A�'�,K��O5�hv��`�������X�w ��}yq����7��V�ތ���:���L�</q}����!}j���|���N£KF��5��gg��p;R��қ�@(���=�r�O�~��..#Z*6�
���it8�1��n��K��Y$��4�%{5!;~(%jǊj�� Zǿac6�A��}���t޺M�tnZl2�#/S�s��2�Q&�4�k��=����Ep�Id�v{�+}��da5-���"��8Ƴ�rGn�.�J[1w(A5~���64���� j5�)W#�"�D+��Q|���(橵�8��8���E
��"���$;�N�R!����N�~��?��M��Ow2܊��γ�:���tR)*��B�/�f�9/�X���N�%�"���p\�W0�ށ^�O���Oy��&�`�B%�|��1�(�;��[n�_;��lh5L��q�*�`F�Ԛ��0}��-:�/��թ�_�d��̺GM�*�iH��2�1aH��7H#�_]蹐�JG-m�%��0?�15+�<�X�w\�m?]�o��"Jp#�)O��<�c�^)>K\;��}b��ab�ǳ��q�9�ֻK˴�B�}|~��.���y2��F\�N�����L]E�H7�.ǳxN����]��˃Ӈ��TB\jY�k�$��ƅQAx~�澸�ʴ�.��00���Ί�s�W�0����y�@�d�Բ$u��e����PD�����u:���ڎ�
� hUt���΅����K8��"3�����2��]T�xeh��R�e�%��&)��
{�L�Sax�aԙ�#�Ґ�Pm=�#y�Ad�NY�PR��c�Z&*�ݸC�����Q-rӵGV�4@"�jd#����BX ��i@b>�Gh���&��G�>�D}�s#���z�
Z���!)ҙ�Ի�V0���t�Ԇ"��B�'^�r�a!�gZd�nv�b�F����'�
����[�K[I�FS�J�<֌d�,1MO%�L]��+��[I�j�TW���uY8<1����9�2�)@Ta>�3��d�M����)	����}u48a.{fPG��-5�*Y$�ЦC��uIR�Gg4��	��a��Ԛ��Q�pҴ��#V�ZdK��iz �ގ��OĞ��Ek�T���F�ߏ��O�r,���.����W����&�����*iO�H�µ`�A��ǳwبN,�XW�v���0�A-ze}F,�"����,�$3�C�fe8Ƒ�ɿ���@o�	�Y�ԛ�&��=�d�%pX�Ums���8�B��ڮ�ҿ��2s
Uڤ�^�[�1��.5�2U�o���\��{T��\@��6`Ȼ�ʄà`-O%�F�&�� ����-��'��2�������VÄ��izE6�B�ڥ��c��J�UH�d�s�(mw/�`�T���3�*l�JD�65��bۣFj�q���ݬ�60����M��TR��!ʀ���s�GT*h	r��B~���2j�b��F����C$��ϩ^���z� ��,�~��7��XRY��9x^` 9�Wi�����F{�)��P�s��N~v��ͻ�?,?��:�q�+���׽�������˻�wSC�Dn�Υ���ؓ?#7�jً��U�Y0��V7����n��n3�o����1C�N�%���t�{�}}��������?w�e��ϗ�O��T.�9;ۏ��B��{�����қj���Z�w�٠Z��'�����WB�j���hμY�{��p�r����������>��o����J�3�o>�m�e��v�ۿD����{�ׇE�{_�:y���@Gg�\�,v�������\��{�x�~9�J���-m������}��˫gJ�;vD�n~�|g�n����]��-f�L�s�W�!)�����}!+.���g3��֊����as���*�	���+�{K:a��؃W�2��Y��1(�	]S�u���mlv?%?����i��7<+K4�|s�#2����,�1R;��C��8%�c�Z��Z��Q͕�+G7��Ww����lџ�F�����}�\�%���@�ii D��D�*x�8 T�͒���_�D{��!&܀��uX����)�����_iQKџ�}�lD[<-�?�2��ӊ��!s�Q tlNf�|�~�ixhj���(�x�D2j&�O����T��Pq(s����Ä́�iv�%���1���J�b�4�z��e��9�,h�Z��I�����<�c�f�4�c�	}�!�&/�@3�2�(�@�T��~����(FCy,j��wU�����\���FKT�y��l�B���36�Y/��zj��{
��)`2=�}Q����n����l8�Y?��~�1��	�/�J�%�k~7}��r7���y�A�:�Y����-B���·��v�s�l8��	-	-{[y<����BM��a��!�3�0��16���L:>�,(�فj�
<�m���uKD|Qc��cH3� y�tȈ�R������C����$p�]N����oюO#n��{�������v��I���Gá�,ei2��ۯaB�k��p�p���ܝ+� Ӡi�Tl�? ��
i�Z8��Pe�������B�]���7)̹��:��m?B�"eÂ�U�1Ft�(��$Wwψ� ��b~�,�9D�r�W�#��?�o���\Va{j
(��8_e��л���gS���b��yɂ����T���
�{!�4V��������(��MTAqP~�)�5΄*�tv�C���"��ৢ[2����`v�&�Sb'���(�
&�6;�a=0��^ᬄ,ö$ �l�#�A!��%�>�Df�^�&��!xp���*��C���B��(ru3TV3Y�����Žh�?y6.v#f�C�c0�������ӭ�Æ�]Jj� !I���"��"���Ryac)���7f�T�Eɚ˂���v�%�h	٘mc;?���7,N�幝!��)t$�0�@�0S8�C�[��c�z��>C:E���ңm�]�}h�����b51�O+�#X�B_f�Po��,�ԓ	��ż�L|6M�eD�C��l3� �����L|�@�6����D��'u��t���p5g �M瀨��&�^�x���34э���e9���_aЊX����O5�E��^��!hw#���I���=�:ެS�Ow����x�U%�	�~y�� :@ſ���T��^V��a�����-0���J����8�j)��)d�D�cjE'dr[]��e��&E3���!�PQ�\�@U�ebh98r�D��C:Ç�B��Tn��Ѧ�h�pv�3ʑ����r�D�b��P�\H�W�YT⦌2�%�SW
@�p~-!@���,�-=?�(Pn�h�/4)��%jj�*Q�p�Ӭ�`V%��\�MCZ�t�JP�I��T~�RF�6 ��~�,~S&+�@>�2��0��H,jL�)>9��ZD'�s�b���ѩ+Qю�A� p��T��U��Yb)S�P����SM>��H�Q Ι\���(+$>��qR�P�)� �ҫ7�r�D�j�ɒ�)�)��Q���nd����JK���R@�T�$~�҉<!��,fx��}/��h��銓Ռ&9�K2���H�)-�Ȣ%Rc�8B�#  �*�xj�i��N�N&�H������Aǵ���9��(�#崊i-�F�U�R���F�,8�~:	��n���Ǘ�j�"��M!͊&U3���ᴺ���ꦟ2��-�b�Y�@���P�|&��
oG.�(7Pz�t���1���)TzFY��HDc�FN墝�q�M�a������d�f�\?q��ȏu�&��:LVV-є��ȲoB��k~r�������㽦�"��t���U@���XWȕ�)�A�kR"����R��V�|�F�0�>�����}lR	�����V�?���S��zny�������h}|���ZW���s����Q��7�����U\߬����N����P_����f}F�3���.=�����J��z�x{�?�O���펇����o���p{x����OY����n�)���_����@���Vy��FQk���+�#�j���Eӗ��?���.�r�݅�������;K���o���.>�?���ߏw�=x냥~����߽���y8z���>?zNu�[��x6��on������\�t��O��n��k0�n�[�<;���t�q�vm7xW�S��;��R����:�ҙf(#�:ؽ��R��{��� ��<���1m��Ԥ�]F:pm$�9�	ȈG�K�72�D��h��|!S�%t�`Yƥ��ȢFV]#_V)ьԘ(~��d8��fb�|�����;�ҽ�[.���Pf�9�v����8О��Tˮ�!�^�p>Y
�-Њ��3x��@HS��a�́�R�VUj]�iOB�2��ZG�V3�v�B(�U�����sސ�4��#�Y���@z���##Q7S����|ƗR�|�jCc����)3q���������9��RFf��]�O��tK+%N�m�.d���G����xޫ�5����2�# .GH����FH��A���e�ʆ�>�\�̌�8�����q����\c�9�\�ؑ�wE�)X7�+��r�4C4�ű����Z������	BSv�zT�I�{\:�p���	o�U^!zL��M�-5�si��8M� �ɖW���1Ķ�������T��E�� x�WF�v�4���}���&\=�9���V����'��'1����4���e34���D�R
����MJ�9d�q��������lz@{,D����-�J� �yRC�:4�By}��.���j�_a�9��ֈ�����#�֪��b�ѷ8h�S��֪@^Qz!qDa��yq�dR���VZ�zLüb�JH�!����Z��3�Rl}YD�G��XJ�+�J��ot�y�|ʕ�Ӵ�4�>�i�5�i#�������G�={��:	��+��8C@/lQ>'���w�cK
tΝ�'O�x��+���K*#[Cָzp� E6�JŴ]��"kR08Y.C_yz�lF�c�%^"C�
#x����@K���0Å�fW��Vꌤؚ@��Z"�b1!��('����z![���k��B4xف��ҏl���]#<s�&��굏�x��g�wf�� �iχ���86^���"�f�$Q��~��0�����fj����Lo�r�ֵ�KFᦀ��pU9B��^.�2$UX�?$
Z��o��HT�+Cǩ�$hH�a��<ÉJ���`(�P�0C-���N�a�C;B�
0}k���񲷜w]^4�t���dam�sb=?����vh�����K��&�ŷN��Y|L��2:Z\ly�Q��±�R@?���s�##<��5g���8M�;oyq���Qp˥B^MmB�v>!�1M2j2B�\�5���g��,�L��,�5.��0) ����Ƅkw����2��P -�א�!�W���P� 1�;
��D�M%*r��x��3�a���Vg+v-���xqdԋEӀl�fXa*d��f8:�l|��)���+�gDp̔`��K�f.HC}�3 ���Ly��"k��7>�fd.M^"�St𑫟ZʆE�K�('5�M�W+cF!!�M���!e�c6d��5!¥���c��b#�����d��o(P����@��P+R�)6�w�;Tl8P��v?N=|�����7�U2�?뜸>��bC�	.�V^��M�
-��q`Rl�b��q�$!�Y1C0E�jUI.#;cV�t�j*1̮������<���qJ�6ۡr�z��tM92$��+Ӷ&p�9l�b3�P�<���tH�0x��eg'���c�k�t��ʹp��Ӌ(2���\��b'D�DV��\�����3�!��zQ��N�&)8��0�iH�L��ʀ���b�V-��fh�AЈ����QV $plYJ�>AF��[
��z:���&"
����,)D�'Q��l
�;e�	�#�-�`��M��4!y�����	/ضZ�X��@C\
dm8l^�^�C���pI�Ӥ�j�Q�����(�ț�o�C+��Z�]*�\�dI���֪���-�M<�!��D�ij\��5xj!��Ei���3xS3��5@����|[X=Wj����adC��D�)�=.���VC�*,;�7CC��Z=B!��T�>��b6���P��	� �I�=�@4�Qt:����kl4�}أi��N����`��W��� �Rx[���f��{���@�^���A"V����Jr��/����e��-���9"�I�!��)��"�%""�T|�7c�������@�=������6�Ȩ6��~]�l����Mb+{���^��Q��]eC�W����� ���$�]���?�AD����D�*��T�D�SR_��i�ڊ�[_ܪ�۽�^�_]<�g+-�wD����~�>�賑,g����O��釮���/�n?�ڽf��.v{?!�n�iN�\����VL�;!{��ã�G>1�wG�LI������Oc��������_]K=9�8�9���������o���ˇ���/����7�P�s�����ߣ{�����{�Kո��h)��C�'��\{��з�>�AX3�Y�#_w{��彿������{�Nt�l+m���Vo�5d=�5���5CwƐ����e/Yu�τ8���q��D�a�:@Rl}�]3,�a������4Ul=���Rg�SS�!�|E�\�'�#k�j���9������7�,������N�R�rSEjd=�^+]EV�/��j\%�ŋ���kv�}��P�B�Tm�B�6N$2�f���* A4���!Sp�_��FR�!�:ź�0���u��{�-��a�e糛r���,#}dC��z�ƫ1�*߰��RF���&�Q�hD��0�ٌ�W�I$���(\S1���۲ Ʀ��f=jp��#�W�����,�r���6$�!�f���F��z�%�%e�q���<�cɋ�ˀ��N��6`!�t��CT8�c�c"l� ���(h�V�"t���454^Y�(/I��}�Ӑ�u�Z
��c=�)%Ga��b�fףe�߈k��¹�'M�r�U� D2��2��bK� 685 ͼ�ф��g1�v��r�H��V�9z]a�Ԏ��'X�Y&^?Ӑ�s��7����p��T��f��pYh٤Tb
�U��k�p��R`7�@=��_$���!�Ŭ�aVm��U����	#��D��*H��Φ��2�f�y�Ζ�C�¡ ��8�j���g�y���?�飏>��ҥ���������7}-�}w���d)���a��p?�>}��M�Б�zp�q<ަɖ�z�c���QN�޳egFv�Ri��Xk�-��q����@�k8�0zUv2Հ��	AƱ&*���p�^�.�zhR�k!D �h��GO|��v� ��C���������N'�z���̂x�B�6Ӗ��j34NK'�Q,P���!��d^�he���-��&���K�+ r�咔}C��&ı�@�?��pOI;���G�S� �����w��v��z~�k_��L��,hr��ˮi�H^���Z���
䒈��nS�Zʉ�}��d�g���S���م G�ǴP^#s�����@�l�H�Xj����x��e)�xx����Yg���j(	H�N��r9��8Z�ëY��}L)�ehզL�-u=��C������Y�Y��Ī""�z0�#�N�\�q�TB�d��(2�W�X}�'���A���5e�ƫaVv���I��W�9B�3I�	����!Ґ�!9�������4l^���,y'E��
�Oܰ�x:lY�n�2�BL<����!��ԪA��S_�!��HDM�aU���	,�!��_)���u�պ1D��=�Rr5�t6��%�,z�&��n#�e���Ȣ�	v�TؤR(�@
EeW0�,v8U��@`EsM�W�d����o.�d7L�aj^���@���h�zxk�'�w?�D���\�Z�v& e����e�DcWIe�������y5CIC��iC���r���@�&�6�!cf$����z�0�0j�h���U�����U���R���p���B��2�f�HU�鸌��:`��aΊm�+�0�R �JZs�fAaZ8�ް�WI"��LA�&C+Dy���+�X:�hѐ���p�F���� G��Zj�������J-/���pC!E�-��2p����F�5�siBJ
g�Al|m�2��5��t��#|�R�el���U���啝r��n"4�VZ�D2�a6�h�bc�/��gĄ;o�A��0��z"�����5:t��8�ؘ� �P�S�&�>�
(�r�j��� ��3��)��ꁣ�lw65���8�՜=�R;}�N�0C
��6�+�t*�t��VR���=N�JH�Dq�o�@���!@4vSNDy%Qj��2�V��%-Jx�0���G�DiRG�;EzmD2�4"���/k��	C�=��%ZY�}L��P����e�����Hц"�V�ʴ�2�,�]����"�1��;�&��C~+�'�s�b���
�T?%��+q^�&d��p���^��!��F�f�P��WƽQ�j���\�IDJ�u�Ug=>f5c���	�5��0 6W�%�^�۶r1�t��ͨS��R'���$���ܹ4Qՠv0�����o���ң>�b��)�[�k�Q�����Kj{�g��u}��'�!n��۪���/r�V�E����T��'0�)�ʇD}���WN�w7'�Ďv��w�뽎��;�q=3���H/3uz�sE�c^��;P��k����=�����[�
}x��r���C��xh��O<g}pqs�#�O=�����9>���/�����5۝ǒ�&p��O��5�/��_�{����V�D�L�/o�w�n����Pӫ��dU��"颺����l�C�z������1�#�9����-�:��(�QqD�.�    IDAT	�[n=Y��XgIjQp�=�0g���*�V%�5��=�FӐmp�ƕ ��~En/
��nqw�������:vC.�����j-���p�p�;�a�쾍u�l
����	�f��n�{)>@e� �f�S�e���-pR3��6AU�Ճ��/B��j�t8b�!΃tꇤ ���b��UR�8&�)��zXҐ꤯�ՄW�)�$ve��i�R;�����պU��T%!@��,
Բ��A�akl��ِagĿg��BH�\��3hys�Չ��9��4[/�=.���n>[7oCd[Yx�,��fЁ�+ �^����~�����)��`s5_Y�&����&��>���&DI�������4�	v3U N�ET�����`
L�����1L�����2�z�Z��t���o}�[b�f�<�cE�w��ɓ'*�R�N�Ī���`P71�Ɩ	^>Ci�q�Ϋ�M��V���w
�4�
��[��q��y)Q��A<p�gj6��4{����A�ei�;��#6����꺻g$G�����B �z`�V��%&[m-���5����ԋ2|�Ԧ�lM��r�-�2�1$X��i�aT;�R�?\� Ff34���!�9��v�{�6��G.O�=z�����	O��={��6�|�q0�N�=����~H��?��%cҷ�\8��v��,�Դ���]��h|�K�W�4|T�(dm���j� k}̔��FC}+�S���a�3�¥`kRSA
�@=�KC����2���(�\ta�%�x���V<�b�ڇ����h���:�#d�e���F��V�î�jpᲨM [��p�z�Jv/��jr)��+
��)�B��ѵR��S��� xPM��J���ҡ"�4)��.�>HP"
���.!���g&�J�5�j��2�*q K"�(D.C^|5`�*�`Yx�Uhp5�]ןh�d�B���)�3D�5<�L�NR���G(4^}�l
���8�3L�Pk�`8��p���E�p��Y`�Іr�-�5� �
�h_r�}�C��� �E�����(�{�X��ƐR�S�\\�z:��Dk.�@eT	�~} 2W�th�p�4�B�L�G�O0Ry)�EB�jU>�2d�p��S�N��X4L-f+��!�a�PɈ�����N�pf� ��<���%�)�K+��y�g�F�1"������+P�V3B^C8[+*~j��cH|��F�R�Sh�eX�΅ֵ�\�����dC�0Z�y	�J�$��o%U��HL��,ȕ-c㮎�+o��K�� .��P(u/6q�t�
� 6���RT��9
����TO:e<�®�@=�V�씉L܋=�YdY�eAC�H`F��1+U���q� �����%����q����E��t߇���a�~2�����P����ᜨ #2f��N��\d���KaXj5CMx=|�[�ְ(�~�j��1!�H^=۫U�!04x�v$䪤
ǁk�';4C6/�������1��q8�b3/��MY�[��u�ū���b�.cl�
Nd�5�aHR�2�&�Z��Z�B�*.H&"�@6�O3�R����R�N���a%7�:` �l�5�V�����->�p��MB�Z�qTh.��-&�^tBFYH�h@��	~��/u���B�"֐W,[CȮ��t*7M�VC��in>��a�tbVOv=f�cY��@���f ���L�!8�)��R�b7���DJ��0 >$|Ø"���d�(����E��n�tK�^����� elmZ�Z"�i���M�+��I���%|����fH���ǯT�3�eEF�eȆ\�W,������yM�ֳKa��P�!3��3����,�^HC�b�k�첬��&���
����b4��z�!�ahRhB�Uo�%"$�,!R0&݈Tm}�"d������Rf�˨��Ūv��j��^�Dq	/�D�k8~�*!(ba���-;B���ϰ,�
�5dC�jݧ�0�����4�I��� 4q�*a�"�Y��<T��E���v�aT�<�R����|��D?��s�K��<���ٻ�]�+�L��Vj��u�|��V�N�o](�|��ğ�4] ��/{�����B��s�>�ة;~x&x���|������vq�f���7����g�~�=v><T�y*�i��U��z�9⮓Y���l������t�}K6����W�7o|�>�������������O(wG�=�<������+�����?�)�Ս����g;=Aݟ?<�z���+��<rВ��UZS�D'���3�m��!�v�3��'����/���n?�)�]Jw��m��ݑ��M*7��o�zR��~Dt`�+��	��c�l!��h��)��H���#��4�ogm4���ݪv�ٯ�!(LF^�zj1 o}��Iċ�ctBxSKj�
Y��D^!+�����W"�ZUF/�����՝^����o�(��O�t�=�OM.`�w��m�*�I���"a���Y���Z��h�$Hm��.W�πȒ�~��߉B`W	�_:"��J��U�����fi����^aD��&e�E+Q6B���1dgOj���93?Z<~��I�0�^�T��(���~ސ[F-�n�W��e�i�k�Z+i�-c�v�aى�t�O(�;�dՆ	t�1�C�JO\%z����6��ҹ�
�<��dh�є�)	�&oC8�cc��&X8��'+ě�R5kR��bz�z\�1�=����gϞY��6�Jҽ�!TJ�� �T��qj��>�$W�j���pL3&\�9�×�J�Lޘ\��\�\��z����65CQ\DZP���~�x$�`qiz'`�j��zٰ2B�8Z�R����l�U9���X���cn��E�?�kb%�WX�4�[-w�����D,ZL��uN5�d��+ ����Yse�}�YX�:Ƨi���H��h�]�z�-�_O+_�֥<
N��Ǐ����{��4�y�?"H�x{I{y�_��P�ˁD^�2vZTޫ����Ge���lÅ�QA35I5:@
h5^� ���Z�B��p��&[,�%А/6PO!2C��!�U4�*	�+\,oC����1כ�a�\rM^�PT��#8���j��<5=ZsW	qMl\,\B�Sk�@L)�e �V��N�0 �Dq�m�]��:�M�V�!��P|��q�&��+'ʐ�����s����XI�\�y��!�K�J��Є����-��\�`�}��Af���aC(2zmb��UU� pe'2j�D3B�R.ʞ�T�e4��b��	&nsZ�������_<�z���[�g}��E1D)��!Dx�-
���dm�=���Z-��0�R@:�j�S�O��V���i�ȭ�Z��_.���Gn�J�OJ/�*q{�wƤPI�2�a�S��6�h��H'�V..C5��Fh:eas�F0LMx����C�b����QKʬ�%�(΀�/#���y��kpFMl�
B��Rc[���`��?��)��e��dq&�@`�Y�h���\�:�dH���j';GOG_�-o�5)):���b�SD�nbK-C1�&ŀ'����4����N�1��A�4�4v���.EY*�M���i}�R�Һi�E�4��+C �����޽��L?oQbף�[C"�J���r \��Uҍxw-
R^�j+c�e$D#R_��hq
���W��DȢJ1G�>o!	�5:]�����b��/
mj ��2��
gs%[m���P8�(CF}�}�i�R��h�	ɛ~�м���Syzj\��ljh���-������t\s��z��1�#R=J�ˈ@��1p�e�b`*/$f}�p:�S�\1���Dp��ݐ�Q�\l��
!�T�N\M_�l�k�C�'��Pc��IGh�Y.L|`��Ke���0 켃��l:��,�	�(`%�5�Ώ,��x�@��S÷h`'�5�88Ă���SéN�p���z��HC|H:��a��!8�∅�5L-�ɞ��E0^�Cj�Z�&2�rO��od��g��_�#2�5=\�iF��gр-�F_��9\_�^QDc�ҧ�1$�[X�!�h��3)��\�S�dI'��WT2�\��H
�G�$5d�#���#
g$Ryz��G�ihs�X��rx����O�fGY����a�z+�����@^*op�����Rن��eGc��f�E�Z�"c���O�";/>C�����І�hx(嗩.D@�~���5���m��G��_�B=�eK���&>d� )��8cr!ׄ/����8/�U�b��s�i&>�T�S����x�B�Խ+K��ܵ8��g�zศ>~�Af/�S�F�Tr�/`��;���*�Ϛ�:f�_i3H��׾R�%S�Ϳ����Sa>�)�C��"�t�or��끟�2�JZ��x�T���r���U��޿m��8���������Xw:�`��m�ũP{��Y~��$��h��C�'�v�������[_�ߟ��>������0���]^�nO>{����|N����~A5�m�i���c�2{�[k�����_�t/K���f��?�y|����^������iN��W;A�N�Z�'�_��W�"�<��yl��[o��f����5`6��[s�����u��$k�Y9	\N��\�ڽ,[�w���E �m۵�e�֖Ί����կ3�:h�h\z��h�/{�..�>����w����p��rF�D��'pz���������*K��^��dcv_�〟��'����ݔv��z�/Ql��p��V��k4Mm5��tlL.%����%q�S�!Y[f��K�-�����ɲ���;
�c�h�8ͽ�b��B�d3Tb��R��r��7tJ��Ds_�������PS�j��)P�(�Ų1����5.��\�l=&N�8M'�|�U%	�@�a6${X�ax
�E���\�M��l.v�ʎ��F�|����롆m2�klQ��(�E�P,\�@.����e�e>g�� UR[�Uة&KM#k�;�k�x{-0&)��뷸u3?C�\!�8�^,�*G�xz6Y6����4D34A�Q�[�_�җ�( z�ML��_���a��WF�vWO�|&�Q�ld��i��5��y-�Fs�5g���Z�	�$E�\B,�j��(v���1��B4�"�x��E�L����-u�g34!��VU\@�)88��0��akF����V �!�>P��"tؕ�f���T�$�b#�����l���֐M-���+ ����Uyp��;w�h��y����S����MǕ����>�ߟ��g�t4y�ꑝxWR�n=��#�/~�ސ�poH^��ԕ��o�+Y����cF@V*�
��7��x�ق@�6�N�
�le�,�&2Y8L���g� �n��jʕl��ő�P /2PUi�58��O�	,6M�U�p�S ��)������ڴ��uRT�	����eǁVǕ�Te2�@��f9��cÆ�H��B�5�yQ�X���?�Q���.�~"��w��k���ő�U��i��(F�>h�~U	��b">5(�	�y��N�@���U�`�,�(�mȞ�b�_k�5x+���Z6o�F;�9&bF����C_W�i���и��}v��l�<�Ć$"o�2v��	����2�)X|xR^�{�~/|�f+}��ciK-Qϧ횥Hʾ�eK�P�Dz�Y��������x�7"j ����v�C�šɅ�o����G)�l�\����UΥ���]�!�F����X���D��
�6^�bWXk�8D�����+�����(�h�(da��]Ck�O����X�v�\�hŲ5��*`j�Ol)&>�zͺi�D�Sv:���Z��k����9�yS�步���-N9\cB�S^��+�&�Q�d3���lQ��k�pj%�e��K�G��K$���8�t�j�\�D0G(��e(#Y����/���S�p�!�� "�᳁iB"j�z��h�<CFk�b�[�ᠵ����I�1��&�FS *X��fW��설	gx��g5( 'G�J�RF4CL^�[�N�0šr奖��f/W�� Z���Qy�qؐ.��j;,H
�ʓҀ0���y�:h��4�r�l=BQ��Z�z�Yg��Z4!�eat���	ݿ�Tf:�5:����t��ńj�|��p����"Z�)��)h����X�@�E0�����)�^#���2��
[٪%�hG(bj����H�(��&J?ޤ�Χ�t�[�G�����f�T*��,�KOְ�y���U��	���8�b�j����P�r��`̉��rŏ9� ��2;�T3ex=d�ijQ}��7�s;R��N���w�0T$��r��?�� Zʉ$d(�/d�v��as�h�P,�� X�P�L2egO�L!�dSVC���$fj��Z�@����\�^�Z��처��,z�z��(���ʢ��b#���HA?�y��*V_�ݝ�D��8z�����_��k�!UX?AN�~���l:!�Q_�z�U�aF4�*n[L�!��1����Z�${�K����`�X��h[�u6h���{ͺUUe�U C`I�0,�߃�
f�5�_!�JG�f�J1(���;E~5���2��bU���V,����\�ұ�P`�j�t����d)���Ԥ�n��D�HV�r��a�5ͅl���v}��\�nO��M�5|�Z��=��~w���xf��
�W��폮O�5�x��s�S�7��\j����zF�>�x�Zo��-E��]�۔�'q�VZ_6���w�ެ�ݟ����=/]�y�x��~�S�Jyw�<5o��ۢ��|�%�v~���Wn!�����O>�p�X�6WZ<���3>�yv|���?�r�������=�T���t��3�O�|,�o���5�gR}E�/��ݻ7���ЪY[��������D�D������W���3����:;�n��T0�$7��-\���hG�:�
Z)�1;�z��ru���_�vgk8�r1z	tb9[aF��'{ۊu�������:���&/f�]�R@��#�,l��0L�>W5@2D1�M�+h�Dꥰv�ָ���_�ҝ�nå�%�&)M��k���E.�MQ1%��
p�	asєB��&����~�����T�(���ɂм؝jl^���nā�ǌш�l��" 鰕ae4�z_k��s+i"�ާg,0)������,*2P��ͷp8#;�l�F>)��JY��4����	�#������@-$;���*)����(i/���3���e���/^���r��e���OF�(^�._��W�m�Sa�nS#����(>A��$�ӥ$j�Z��VX)谫��/��	��4
�-,~���ϥ�QR5k�zk�>�gY�q�L�-de������'>V�R[��sM$BxI�eH�KWzU�,ܰW���
�1�[�D(@\��U9����E6Ԫ������{}��8��*�W����aL�|M�d1�˥?f5��VT%UI�y�p��$���d�"����8pC=\�k��9{I
�Y���a#��MDA�A��:�����r�a���,\�����j�z�f�+ò�8�{�'�ϟ?���f�G�ɯ�뮒N�M��J,[#��Rp��cH{��O䷿���]���`SrQp�P��^j�Y���`"p
�Y!�U�Id֓Qxew�]��En����� J� �&��[O6;�lC*C��1�|k���%���r��5��S3�c�ŪGO_c �q�ʶ�+l�e=�\��聆-�^���)�W+'���`�Ԙ�&�Y��zB,�͵�B��Sk����+�-��l�tM/����9D�_�RIv΃�Rx�I\"��U�Q$�?���dq�]E1L�ےp��q��\���F+^�U�X�(�0�ը5)^��P��Yc��BF�� �_�[�i������PR^q���Zy�@�R�xR@�qa��R`��7~_    IDAT7d3J��ڐHY�w��A�[�RV�my��_lC���Z����S�[^rg��e����q��0p��JM����N
���V�KD�L�Ő�4��zǧ�*�p��SH�Vx)c�-�:�Eqi��qu�t�y!M��4�oĻ�n���j���!o"J*�a�d�q�M��ʫ�媱_�����殤�S �w��+$���كC�(�hj�Û��LX�뻆TF��Yl+c��#�@^Q5.Ɣq��C�\��bX��+��\���y�>�*	�I6��d�#��K?F�8�����������"b�WI+����&�P!�H��� z:�G��S���.u�%��;&�6���s�fP!]T�+/�6_W[/V: �q�P!8��_�N�\�^Mم�H�zC}:��S�}���(�T(*�!l:Z�-;�谵WtB��'Š�&�����u���Ż�,|g�%S�ƀt>q v���X��#t ��i�z�,\��h����\�l�D�!}�Q�҄tH
��\�i� ѿҀ��
��Њ1+#M)�#T�~�q5��%�����+ܰU
4T0W��h�˼T��B���eac��J�a�1��&$�\*!ޔ[�z�%b��B9&B�t���둛{:4K��G�ٰdxH����q4�N�b
�$yCR���֧�r���V\.ً�߰�����j��g�1�Y�~�5�C`�i�h:�t�T��D`��-u!���3��
nY���Bf�p4=eN�b��Q���Ϡ��`��ᆕZ�[Ī��4�6L-H�@6�CC,�>Y!4!MRΘ�{ʦfM�N�-�D�fW��74MHC��eL�	�י4� ��
�q�H\U�6d W�a��#UO�2
aK����&ޔ'��pz�T	��5���ڀ�s�Å0��j����K
�HZ`v:��l=I2#�EO��]��:eW�Xu��[ȔW:�-A��`���M�/�&^F���h�!��b����۾qaZU5���2*@�*��MY�F���e��U뷶E�J"����z�߭3f��w�n���Y���7?��=���>�Iߣ7�1Y/�=��ڲv�#�ǚ'G~8������j<�n�:��*C���鉦M�����g�����z�ݥg�'���������/��R�'�������L�'���?�dw峝�]�p����^����ȗ�zعN��l��<���#����g|�Խ�3_v{�xz�������=�݅�O�n/-���N/Ώ��'美������,��o�gW���k��Knw��i�7"����?
zz�Y�>�y�p���c����'Po}v��<۽����������/��]p��7�����}p�}�@'ʼ�g��#[3;jy����h\&��!\�2������v�x�n���;lw�Z�A!;Cv�~c���%�D��!\j}e������/DCȨ�+�R`�IJ����C�A�������ʂ��'��B����'�����e�����v�.�l�2�t��b�2x�7l!��R#Ȣ�ո���È��8	��*R�"�B��zu��© �M��G��4d4����R������G��m�J���6�D��}��B��*�7;C�,�euٓ+�,GY߂#L�}��^v���yX �遑�X����Y"�S+l��#��NЫ����a떦��ޛl��hy�\
n���]g@��Txs�,�~{��N��8�c3�Y�+��&�Pyͽ>/�����A�5��@H�˘�)���ɚ�yiN�,����h�ԉ٭r'ۣ"�+�z�����L�T�d@F��BG�y*K��6Z"�]/����`!l:*n�@HΎ�0����2��(.`aJ��A�Y��*��e��F��R�)�nY+6Y��A2�I�]�hU(
�?!���A���9��Y6�H1̢�*o3-�@+�0�M�w��jSy����0�Gf�(�V�*��}�g���}��� {��?�zI;�^����5"�q��8�Qsu��0}����ld׈Ǐ��:3�	l��x�Bȼ�p�=U���=�RO!�fg.:
hY�tj`4��/J�,[��Ro(D,�ٔj��p8��T6Y�Bh&Bǲ�-P����l�	��@
���R�m(����k!ꉆ� }�K�p|C���K�Ydx�fLg���s�gAR����h8�*���U��pZؼ.�r��k���i���Q)6�f(V�"�pJ� C@�����������}�H���Bm�.w+5�;��4��L�t���h����^CF����P�k�jg!;e�I����s���hl�
��z��4ш��N�0�d�R�����ܻ��2;G�Zu�L��"��@�	���04I�\!ͱ�B��á%Ҿi�E�,5�����fuΪ
�҄��A"��@�K���;�b��0��7���d�V�i�pd�N8o��K=�zQB��eX�#��%¨�4GA�Ė+r���֭D����(Џ֚�KM������C�A�� fk��*2�G��D�%2d�5���W)�k�g����w����e�����I"{GN�J�IDC.ov�85���uZ��z�[���t'��m�&c!��HT.�)��0�0r8��pv��CB�Q@`Wa.6��Mm�85uj�����r1�|���`�d�Jǀ��Fh̛KC6/�NK�� �f���=}LC��!��p�Ap=��[\S�@-=�"��J��m�\mMC��T���'Eְ^I��0�C�D���P�aAl�#F`�`���S{eXj!�hS��(/�%b�4����Hv�p.�V/�������BDU@!�U��+POG��,Qޘ�hr��,5���B��#!B BM�b7�nO#'�\zm�*^�X8~"G����l۔���S�M�KDH��8���ҪS/NK��!���J'<&#&C˕,[�oȐB�!�!.�)���P��)t���	&Δ!oY!�k�;��f!#P�Xaq&/�A��p�hDxS�l�s�@��Y�
�,��fId���H�Z+���W��	O�\3#^L�!��� J5C��@4ކ��������0��>��s�[�RLl$�2�&�U������u��\�e)�!o���i6�!�AH-ev�"��aj�\�f5����~�Kfx�������T � �-WR\��%/����b�ǅ�x[��Dke�P DU�Sލr��/rˋ�U�d��7L� ���DZ"!��7���F-�G��s0~y� ��ѥ�0�B=���~Q~[���<�X���%%c|%	��v���ЏU��pʘUK0\"�[�G���tp����tC�R��u�S�Jꨯ\~E������������^����p�̇���k���߉�=7�*�M��>��p�G��ۛK"�_Փ9C�lM��v�x���ȅ�I���v�a}�S���v]:=�P�̞�����멨߅���[�*���Έ����>�遢_mv���?{i�_�`��އ&WA�p|��z}�Ǘ��i-�Ԏ�>2i1<==rfo�׳�k��<~y��7^�����d����������s����/^���=O��o�_ܼv�3��z~v����'�����7�/N/wgd��|��/v����zz�{����WAU�٨�!�����~-��b��={fO}�H9w{|��M��ϟ�:Ez��9.# �6ߵۖ�#��i�\���*mw��ې;T�=,q��?���7�!��>��r�Ð2�V!ٌ�!p�E��-{�We��pm��hB8���8\F�l����� N�8P)E
�3�U��dZ�c�n?��O��s��uâE�/V+E8�^��o��4d�Y�
@����`O�j	6G�&��O�q�>z�����H�y���)	�0�X4!��qwT��T6�X͹�ܘb��;�q�t�K�eg�k!�g�љ���5:@��z�o��K�3�����h���SЬ@��b����&��E,˫ ��B��sI*���V����h����/o�h"�aZ[WJ��_�X7��r�}�ͻ�k��� ��h�=�=m{�A��H���(��U�w=�I=5#�)ΐ��ޱ�<�( �a�h#������&Bb(T���H�k����w�}��M��� P`+O=�4�nM���zf���ZAZ�O�$�$���U��Roª�S7�&V��l�,.3}�ͳX�VT��iD�[YU)��<K� ��!D�j�khE��`�ѴD,�m���o4���jZ�Q�M�Q�E�j���\%eS����r�Jǎ����l��2�>0{�r���!8��fQF�JB�!��#DF���f�(�����{�ݛ���z���F����I��Ξ��P	)�\N����<��J��,�"���>��&>���	Q����d�m:�\�,���D�Όr�Y��Ig�
�t�2y��+KH�-#/C-TC��u�3MS�q��x�\�U+�a/"�S�u���,
Gļ��%W� ��cz��h�
z�
��\ulol8�&\
M^��`"��D"@o�Ȇ��2�l�)@�p�0�:;����Y?_Bl�!>Z��P���?R���H!H��Xo~0J��(@%��lCӄJ���SGׁT'e�5a�l�22�[5��l�l��B �U{(�Z;���04�b�rQFkI�����!��z����'2�0Ld��xq,qj��w=�f1C0��c�E5�!����T���@����G��)j�Зt�)T�(��h\y�Zʥ���'([�ޤZd���adL��
!%�������~��Nj����[�j^��\8�y�*0~�E�gX����W0ZC����!fZ�z��Xa@.v�l�R0j�$���O���M�Ҽ,/MC�%M65 ���!�.-�t`�1(�����@.Ȁ�/�Kz[�z�p����&�M%�@"���e@�!l1T��@��������) �^d�$5��ٵ���K7)v�
�0WH"z-�䂴�t���ճ�!M�t�O�c�Z��K�;\�\�7N���P�?e
2��a�!y��tA��ҁ�;�h�	7Ԧ��CF�
L%Ma�!�)_��y� O:��!�Mنt ]�Ny����"3G�-�ƽ;�l�R�[=dI���@,Z��Y��r�P���D�����SfT*C��UIR@�]!�M�],~��t�DM�S��lL:8�q ���9?�Z��3��^T��V�^ [��x��s�__��dd�Q۰���z >o��cF�.<�Sy.2S$�V^�� �\�%e�\[p���'o����
�D��=��1:��F*MQ���0����
�Z��Q+*$��_�U`��a�n�z��\g�d��Г�E�`��\�U�����1D�!�@������)u�M��m�w���y���J9��[�O3���P!���E!ᐘ����82j�S��V�)L%��@��0
�O1�\����dX"vW�J�k52�hlFY��J36Cc��La��ڄc*�W��Q����q���X1��
4�$d���*dC4�C[��^1����$��p������l+�G��0j1�h8C��#8�� ���l+�Kxk�?�Jpt�F6�(������J"�U��߾��p��/<82��wm���ˎ��RIA� �yf��Gf����C)�
y5��`B������"�A��![:^-Q�\ruGk�%��ӣ뗗������^R���K���������?)��N����O#��n�������pizۺ��m׷�����s��ח�j��ߚ�r����>L�"a[���}%��c�>Q��uc�׵�v�`=���C��g=I���O!��__]{���r]_Q�1�����Ԟ��\��.N�H��5;�l��[�=���_�֧D�G�}�����_�|��/oO?yy�SQo�Ɵ�|x~�����������?�ݟ�	壡��_'�Ǿ���
��p�V����}ϭO�ʹ���Li'��^�bn}�U���on�������~��u�h{�`ݲ��As������K����تX=���/�^���2�*��
w�<�z�M�����6^p���^��O�<q�jۯ�ZPL��&.�:ۅ����	l�� C [c;CH�EG2Q��%*W!#ŀ���T4�1룭��]�xM����p^F�8�e�
�������l���S���n��f��� �8Vb�>��_�v\��5��4��N3����]�:u�8�M��mH8q����C㕂���ꇔε���s��S�>��^���t�@��0��H���C��0La	m����M-T=f���*C���)c �����y�Q��r�r�(dѬ�^ �6�8���n[�O`�Q7�9i_���<��/J���t�q�������׽)W6����8з7��>�; �K��쑧Ǣdݎ�Tvd{'&e"�H���^3T�T3�7��Ks��k�B�y�j��a��y�s��:ZD�ǩH_���35Ż������{�%��z���-�v	HT����Z)��)E����U��$H�2�ʵ"��(>
�r)�m�˫�\�@@.��r��L�UP1z�%�����ZI���`
zjR����7,W���V,�f�B�)�Kĕ��-0������h���r1�h�Z?�79�V��B�4G$fՒ����,]Rp�J�5�!&["�W^G�?~a@,��מ�ᡦ��@���C��p�Jrt?~���&���o���O�>�u��8&.�&����`� `��^^E�#mPGB����ͅ 8C�@��Q+/BebF�g�b��%�(��J/
8�Vp6\S0��� �"O�K<P��t]�0� 41�]UA��jl�Ȁ�����\_�	ΊI�a*��f/�HA���&bO%��Em
��A�k�+�X�&��
a���E4N�R�3��~�s�y������P�X%iBdQp��!�z�-?�z�p��Xo*���bv�p����a�;���:�Ph"mB̷ʑ�4��p�~ޘby�B�C���Q ��Pن8���B��2Fn�`��hh�x�ˠ��K02�PY�n�j�B
v�u� 6���~�>@�`���Z3j�*���*'}�0��r����V��6.54�DF��CզQ����*V�z2x��΀L��ABJT�'d�+�ˤBͥb(P���F�+�ˁw�HA�Fǰ@�0�&$�zCRU�m-��)�ak��7��S��	gdWO|=�_��0��?�L��r	D�i��GH9D���Ԁ�T��C��2p��S�z5i^�	���D�ð��"೹Z`���*I�
�ed�-����I��>o��!��Ȍ`!�T)(fj+D_1�O^k_�ԘeiA��4Iq��,٢���!�kZ�d����W�����P�>��l.�VII�᥃IDR B5�E�U<#~CQ��,�K��"$�[��$y��g������� #N��&�xiB���������&�[+0�&8G���p��D� {�4w=|�8M�N�b
���a�N��4�Fn�r!4C�p���Zl���S�3^��s%孟2�JMaZ�`��b*aX�-i�0����?�A�i2 ڄ�5G�W¦�N���D Zk�P�C�锴��-J�i+��4�j@�0j��Lm��~��2䢃�,��,Q�f�J�M�\�@���2DU3����UR��j�0�����IsB��>Z��`��!;K�\�z�1�8��"g�#�
3��C�(4mR��5
��!|e��r�ďmz���5�z�D����(�z��y�B�	�`6B"���'^j���VZE2������۲����G����L��3r5�C�ʐ����Z�ҟ	RS`�Ig1��@�ې���6��p
��bkl5�ǐ)�Y���֝�ؖu�#�"2    IDAT9��[uk� ,�t�o��/��x�O�	�c�,��54.��5�9������6�X��E����'��w�r��첤�Qm�
��$0�0�h�l��}.���,U�fG[:3�N�'�fD����o'T��.���>�'�>���L�`�!�t6CM�;�D��<��S��>!��Z�D<����PH��|D��S�~����R��R���!Ӓ<O%�aCݭ-0ZR��ue��-�BBl�N%�������>֚��'=ky�Mi���k�hr-����v2��'�l[f}:@�	&�
������8����x<?�&赧$�l���8��y����&��v����������o9?���z{%xtp��2
(�s~�NwK1�oU�a��a5_�d=�ϣ�wXߏ{�I������iO���?���[�V�~<~��������<>y�Hy����S�x
���מ�M�X��������홵;�~��G�Ã�CO�������.��t�Ԛ�Z����S�=�u�^�{on|��~����˹�kP?���N����6)�5��o���(�K����w��]k257n/��[�+�0���Օ�,ƥ-ה\kR�%[��]}�h�5ہ�{���p[���»Cv����f�a�ux���N���-�J��:� <���y`�b �y�dAʲ�h�6sKJ�$rk��(�u�R���.�uP�uS�t㗲���\�qк�ڢ��	NNXϴܲ�jU�W=��)6*xm8�8���l�1 $Ő��	r�ubCDi�D�C���N~E��r��n1�0���9'f��3�C��! -7�Rꓟ�i�	3O��Z�Ӱ����D!���;!f�A��'cL'$B�����w��}��J6Nb��gW7��笙���y��\���26+�駟�~����]M{��ù��|�"���,�,��]}����Z��h�=G�yI�--��l5��� �to�E��$���tC�L$���8�2S�� &�t[��ڏ?��KI���]a	��T�a>Z�7�u���`��Z���*��ĠCH6�PI���E�	dNC0��B�VQt��[2�q��'6��Լ���'�|�{�kU?`*"���=R��f1�D�j���c�0L��~6-e&+<?��=��$<�]�wf�)�A����a0��J��4䯜a�%��Y���Q�cT?�$�]unE�V�w���v����~�#���(�0N޹�.�ߍz?��o��o�i��#���8�w4P����(bhU�`��J���a��a�lA8U�1k!Ea��p`�b�������"0��E�1t��H����_ N�U3:�����4��J�*�����\0FY�B�3x�d+��h )�������`����h��jv1 t�i��h�ׯ�l0iUA�}�-�t���i`g��vZ�,�,�!0�[������ӖV��5�YH��B��կ"Q?���}+�,�H٭�r�"�*R,fsɦ	�̮el���Rd��� �;@B l�Tz� 3��	r���l�n�	��C��Oo��e�'c��#��	�I�[�hr��0ю�B�`�5�*B3%<�R�%��ٌh� �ӛ�*�S�,`�,j�E#)j(��P{��Q�L0H�yTDK7������JQ �]���_u��e��I`���=�Ŷ��޵�pm���ձ���&��0�'�*4�0�?�aS� �n)0 ��7d��iR��9y��IUP5����Gb�x�"��-d(D�0'� [�p����Jl����yT�N���sz�FH����	3U���R(Zv���n�1��_
s���X���Hu��"�t(��؞��&���w���#�C9����ARE��,E�����oj�h9�2@�9i�`P�ܜ4�H]aka���ګ���mV�~�xb�h�~����P�R�\"C4���0��P�ax؄��nxR����8@��B�\���	�^`I�@�Pu(���6�B��$�(�IP?�9�pm��S���0'B0N��:6!;NbXW!�f���F� �P�8���#��l�5\n0ڰ��r��r9��|���U$�9'Đ�G��,cB���0�9��8%�j�܆<�+4Q�B��ΐ���U�$�+��4g˛�F˳{�6��t4[!����B��g09[|��.+�J�e�I'����Y�� "�B`���	��JK�29@�S.�a��D~)B<9[���z0�z��a�-W��&U���hl��FTu� 0�ӕF;U�'%;]J�E�n�y��Ӂ�l݂��4�G.c*�c��0���D9�Q#6��t��[]��3��Æ�\�H�6gCj2�aE[X�<��'��d�������x EcN�	��xxOz�'������F^�5�s��OW�f�W��&plE��ah�I׃��#jHzvTn����2`KT�%���F���G��B�����|]��a)�E+��f���D.ǿ��{ls����9�G�>���غ��ӽO��WA]�zv�&f�l�}x�C h�Z��a+#���S�D�����r���w�������ދ+�������'�7����v�H店y�`��n7�t��r�����w_bm�Z=�C�+e=K��y���?͘��x�����qp|���ý~������uY':+q��+n���x���۫��ǧʾs�F��N���C��0r�ԭBrj��Z<��^���m��<G{ޓ��~z��O?��O��z�ԏ}�2��۳G��G׏�x��;�}��a̓���ャ��}�r��X�վ9zu}�gE�����%�}��^��)Q��9������m��n��UDmZ7�z���,�k�.����}Gkb؊���F�#�+Ev ?�;����Յx\�]��0��o}��w}0�ك)�&G�j�����<��yz�{i��+n��I�f�����	0�o��℉�$�?<#X��U�!<$$Z�ȃ5��q�\T^&�����f/�'O�0���=���%�P�ag��𣭐I ؎�t$�����,�OQ l�&�F�[Î)������8Đ��c�l���5,׮Ә#���4���_��_����]�D�ط��^����	�GmӨ ��/=<���Hd�nU1�o�M��z	虓`� C�����545:< �6�]�Ig�䄇�Mb�!f6�}:�q�T��{�Zvl�3��Vܙ�`=��D�d ���}筯}��6���c����ɕ��o�E!��M0s���=����Ԓӈ��th�fR���qd���M_�&�Li �  Cc[rj�]�*Nh?@<���m�5�m/I�Ϸ��m gE7�x��3�s';���o��J`+��JuO7�2�w0H��KH�5J�-0?�UP�ejlQ=�î6"@�QEY��!]:m%
����C�=�[뫴5i���
;)[꯷���b���t��B� Κ��Qی*��h�hx*����x�O�s�V�Ƭj�!#rZt�R�*a ,/3�7+�9ڡ�����!8%��@�3�4S�������ߝ��}�{����;���i�:#x�:�յV��r<�tv浍�\:���j.�+��ۤ��4Y��1`%�u���h����aQ���x�·n�8���L�+EK B갣�D�1 �yv�	,�A ZC�� y�Ճa3�dӐz��~`D9�[��:�*��A/�Ҷ-����ɀ��N�ِB�����J�
�uD"�=��;���wsJ�~n����H��[����u��c��o�mll��ַ>��v��N���:�2�њ>*�,C�38;@`�Jxi���)ô�����Y4�6��\���u�di8$���vt����i���0B6~���0�h�)��K��&U��)
F7e�D�&B�"������?<�VX0IC C�RlMݽSԞ(cվ�f`�:t��5�$?�Y�o5
�1�� `K����%ɽRjll��C`YH��l �< iw�B��4?�m�PHJ0$���Y=6�y-A"W�!��9IEg�Ɖ���"i�K #C"԰Z5S��9[������`�ŠJ�� �����=lEk&�\u���\�ꆲ�"#��t����	5`d�;"���[ȆCҰr9kX�9�d��L®��9���E��r����
X!�J�N�����8J�ι���B�����9�*�=<!+ĩ��ҳ#e���Ĩ����+qz6��p���`�`8Q���N�1�!�1:�.;�P{/��y��m�9٤��`:0y��gJ���!*$���y�)8x�^�aW�!��q�O���Ut�:Rц��B��c����Be��0LtHj@:���CC���yJ����P�!+����&�ih?g7Zt�?g�6�r@��KA�@6���T,7���v��"���U�6�����m�Vq�HK<9���c�V�C����\)�s�	$�CN�:�W���B<�b�/Dg�V��a�l�ṭ�h������쟖Q�,2��R�#J�`c�K��*�7�QJ<R�`j)BCQ�M�CK8Y�luck�D���fxr�	rE�T�!� 5�����/��y��0�Bc2�UFlE�5�_9C~�В,���0��0ʹ68��Z���=��v1^�ܓdC:^�Q?-�4CG ��;)�խ�3X��#���1F E�YG�l ����Y� i!H�<Ѳ����)!?)��B3�R��!��%���ԃPUiI���M��W}�>+W�ِ���1LK��C��a�k)=���0jX9bL
lî}V��D����<�Ps2E�^e6�!�(����}<���G-�s����Z>W�Ą��� ��Hk&έΚ�n�8y��x���(��Y�yn;��l�a��?x�N����[}��:�������~Fs�=�S�u�p=��
����D����Nw='$���nM�9�o>�ۗ����;�&�Fq��
�]Ze�����/�?}f���V�������w�j��ˣ�__�J�Jz��f������ԙ�����j�C@��t��yf'�m����啖�nN|���{yu{v�����}w&ݿ\�z{xr{|���У�G�����ó���_~���x}i�{���<r�У��.�ZOh����ჽ��~b��#w�\�����T��%�~�{6��<:׭�c��'}�z�1�S��?>��L䪦+��<7,��+�C���rz�x�����D�kP/^=��n�|��_��O���:6G��f�����zX��B��5�m�	;��m�M��0����Nz]�!g{>N��r�l�a�9�<� �,�4�<09%Z^��-���b�Ӆ��n��Լ\H�4,����0�<D-CN�J�e�a �p2��*`�D��YH�d'z�c��`3��a*�p�g�k��Ðw�����\��	Ϟ��I�і�\��p��l�����'�a:?M6l�<�Ζ��2<E�d�e��x┢slea����R)��dT]4���:�¶ڮB:Rx��8	�Jt� �9���_?8{�_^�h��=��˴�~��͎w��ʟ��_x����?��<�V�&�.��h���X>��C'N�#d(�ᛥk^�"MV��yZ�����l� W���9!u�Cf�V���R��e���j�w�=���7�DV��Uz_϶�%�Ό�1����X	<�����N(�<D��khn���&�Ղn�@"ڴ��Jl搳�:<<5V���\�����#T��G�[�-�s���i$R"��\�B� &lHv)� ��`2D���I+)��a�*Z�6�:��'�G��V(��6#�R&1� ���a��P0�x�������##2B�۸����G�-%���:;���ƀ���,ѣ�}���lhs;�Hz;�8�u@%�R��^	^��׌\��n���6В��!� TB�3eF(��P3�B� '�����&
y��L���"A�O� �!�.���L�[љH��	'CT��l�65NH�t���J������d(�F��Gc�I� d�A"T<��H�f��W���d� g@�LNZ�B���`���[���[��R�]�cО��a�*��xr9���f&�zx����8}������	�~6)0bֶ�=�=��ںlr�W:�����*�y<�֢o�k^-��DLW���Cӂ�C���u��ժcZ!��DƦe��̐ːyG6|l �ťf��?d�K�i���Z�� +f��8�nZ���d!�a��$��E`�6#$5@;X1�+Z��7�y��o8���~��梷k��D�0�*�Rz
ժ�c��NOT���r&�C�B��m� �QN��I��r�I-�BB�<�!=#BQ��y̝����mĿ&gm�!X-6��e�4P����yI�G"��5�I��WQ�e�6g�y�<��B<R��$�Pg�Z<��Q��`����`ȠI`H$Ro�0�C�tF���φɃ�Uj��8�V)?M�ζș5�t���1Ì<
�c8� �����W��IK	�ΌJ�Q��v*��7d4���?!N 9U��L"q�| !�z��(r+��*s��H� ~xF�!;�	e��"��2�z��hrͅ�=$l�H�18�R��.@9����?Cu�B��^�ˎ-�t(�yM?�z��+�`�r����o�:ֵZ�g:����q�i��@~C��kF�Td��-��ن	c��*�,;�`9��Sh���@���r�\$G�,}�N)4O��o���
��*�xx�ƺS�ͷ���iȀ�3r`�EB7������-���p����SB����+W��m��� ������E�&�O��pVBJ�!?O���-7�aH�М04���|�?��lX��q����#�Jp�^�i��h��rk)�Rx�Q�#���(p���eW��#���,�`�� 0S�ݐ����[�O�u�+WT!H����gc��4?����<!v��<��C2E{U�!c��3dQz��*�8�4�ڎ���<�0x�P���!��B�IKTW����,���Ȱ���Ȝ��H�gm�P	�i;�y� �@���ĐF�_�M�0��ch��0���d�g���U��F�ږ;~)c�%�H�i�g�.@o4[b+']��0��s�)�O�^���4ǀA����?S��r �jј��O轂��� C�:��Cp�6���S�M�r�M\
�A���*�����[Y׍7��룾v��:�?l붛�U9ps�r����Z%���j�����Y_���5߲� �_X�.�o��Î<W�W���q=���ט�*��ў��n_��s����#�J�v1��Yy���������oW�Ex����+?��:�3��!PT!����y��8��u�҃f'�G��qA�����w/o���K�Mӯ�ݼ��ӗ���|���щ�L��|��+��җ��5�ӫ�o.�W��������.��wi����b������j�-�C�t��E�Эc����
�E�S�t�uK��,������FD���Ҵ�A��KLR��@���3�<쮮�T.����J�g�����}�������l߈��m�����*��Kp��N�O�S�B�%�v�!a�E3d� 6�ҋr��۶t)<��*d���*J��%�0R6�y�91��D#�[U!H$viε&���~�������l�APupg7Z�YO��f��q����8|h�o^�U ���!��d4S�!��Aq=�)��$�s��bH��İ�fl��~���XѶ��9��6��*ę�ZٖI��9iNE[�f�E�E[.~X`<�`$'���E9�-݂��|�h�8������>#O�Z�Ѫ\�i�h2<U��B6����\(f�ހx�_�v_�c�g:�����?�2�    IDAT8>�8~�l������/��㐙��18pN<^��qfp&A��(�I����ΰ�vD���&r	?a�9�_�
@�(G��3�����`�ڊ����?��?;�y����kP���V��\=)��d�͓&��0
���b��ny�V� #L ���^�;
uUV�R CH)`�M[hn�*��/e��W���Sb�wo��!�d+1���*���XF YE�3�j�7�İ6�#?�	Lsk����� J����tU�-�MpNͺ��E�P��3ؓ�M�r�;[ق�s���=����{����j�}�]���!��[�}M�߆�A�@^�`��5�N�(;){�sz�j@96�֧Ŝ��̑�GBkC�S�!��\��.gs���a�Y[ZTc<�hH~/��_������ �F������(��9�ӛ�hRx8�(d����ٚ�WHa@
�3��|Ec3�D���!����.+~Y<dx,�����۪ZB ���Ì�:�i�^`�Y���K^bg?��H�l_I�C���S�Γ}��3��μ�<�t��QHQH��餬��KT��D�윣U�-�6�+ꈈֳ�p�g�c.q&&���R3��1�i�B�B�R�����r��M#$�fs֕Qn<+mK4��-	'C��K��t�B^�ާ��Yb�[F�c1C
��<d��1;�V �x6��v�-�V�l�	`�	r����6��Oo �4��a��Vm��Q����-^�u�j��\r֤,��01��i �TRxꁭ?�D�S��T��\ � 0�D���D����^�%6FҐ�([b�*ұѤ�	$'̔ˈ�=}Z��`�+�	�DO���o�󗕿�a3���Z��8W�-�I*�K�9�xxfF�^40f�쌲0kr�Ts�/�&-�]!TJ�*N�J@2�1�Vl� ��S�ڞ��_�D�x���9���Ќhb
���h�(���P�°�փ�H�T��Q��&�e)s�� ��ɭ�f� �Έ����&$Ro���{��<[�!��M0������c�zY�@ fU;/E�3r���)�?6#O[Fv�M�\���y�b��T/D��L.'[
�j/X�3�1���Db)<B3VʔfD����N#�a0�J@���caZ��_3�����b��E6�B��#�p�xJa�� ���BC+���`�ή:Yt�R���P�]�<��H�a	?1l��a�>�Vz��ŵ{|k>$~���nm� ������.�
����	�_�E��f�Y"|<�j���K�
�AC��LTz0Q���IrҤ�B�aYt�0�ހ�ԲVY�t��z���9��hѲ��	�h�~R���-[�a2�!~�A���W�@A�pZi[<$�n�B��)�S-l�]fCR.�9�ae��k�_�&��l�����8QUZT(p-��\��HyT��٢uΎ�恩�����'�]xֳt0��`؝�������Ф�f7YQ�SVT1��t~���,��]�H�������cf�0�����&͢Փ�����i�3�B�Z�zV��u�VE�� �H�wda|�3$0i��iH�>�0]��}���J�O��>p���[�r���1d��������}^)*���ˢ��ggH�m�}|k#C�EҐ� 7����нõ���Y���U��۟˲�"�~����b�jUȽJ�+�rO�O_Z�K����	~K{��=��E!�n��>�b�����޾��ysxu���z����M�gϟ�&ׇ�'�'n�>��yy�|}M��Z;Z�nUܷ��M��U���D԰�5�fq��S_�{ys�1�/=zztxz���.R�^��{�N����GnU>z�Gڽׯ��_>{��W�^�?�����O}E���7����o�����ťᆱ�y��;p�?#֋g@�z�5�������B�q����c��g�2��l
���l;IqAɦ��c�;{�.����S��gOo/���x�������O�|����/�n��^��(�tX����{�S�pz	��mN˻6��b�*����n��Z|����q�R���q��k#l��u4���6�:*�3��x�4���d�S�^�:pm�cC.�=l�"�(���o�Z��|�;lO�t�3 �s�rYh�k�(��doU4v|�,����RJ)+�e^������U*���f��C�IC�\W#]��9�ww��~�M��,�İ��e3TT����,� 	';6��uE'�"�ʮI!D�7$<����<�`��	I�L������P R@��-�� MMT��*��\�.&���Ւ�U/�C/�$7��� ������=u���[빬����[~j��?��Ͽ�����~����.�Ώ�c]���VT�+̮`;���Z�gv��4�԰S��Db8Sc7]5ex�Z��0�����Cco�	�={�a�,��:�l]Ռ���c�=�����9�)d��ɵ]�2h9�PN�_C�CahiZJ��Rg�lN!6NNU�[- F.���iVe�'�� �@g��`x �N���[K&L2$ZVu5fC��D� �`<*�E����!)�܍���#�*�\C]�0&:��^�Иh�;�B14�0�r�\%�D�DȰ��1�͐P���f1z�������H?���g۵ޤ��o�7Jh�`o�toƲ�:Qb�:F��۟�p��^�Nv�W&¶_=�\
��w��{U�V�fD4i��"W��C �f��e�Wr�C�r2H$��n�(~���׎��D�i(8~CxCڙ�6:�C�S��ҦS� ^�<R�H��gT]Tu�����,�s�\�QeФ�A2�%�!�넧�5�S�	�1��o]AN��*��¯.��m�l������]�c�c��<�.aTz @��wmK�n����)Q]�1��Dl�"  �$����BbR�N��ӎ�&�mK�a�y0�'H�������Rl�d6S)~f6 ��0��E9�Ka�E�d�)�'���s�b���NN��tsd�!�c�9k�~���i�' C!��N�B���\�A+����u�I��VE$�4?'6�P-��b����&�tH��3x6n�`�:��Ab8�B���[,�j�R{��e��a�,����p) �f�����cp2�	��i =b�O�g ��B؉D�R�S3�ؐ���u����#�/JJ	lI0:]:�iFeMQ�\�;ZQRQ��xV�������Z-)�I �Uf���F��<Ւn����<R�(����@T!a�\-$	�𰣲��dx�9�8UZ�.�����(X���w�ͥ&%V�P�a/��Җf�A�����B��Ěi��w��م������
ʙ-ԔJ�0@���a$����	�!�HB�B��	[h�`DUE<`e18��i9y*!j��H�$lNC�(�Ec �g�*dHIv$l���8���U�&aw1<�=,$k��B<��,a���ٙH�a���~%:�N���K�#��Ov NT�S��-�(-�z-��g�BlQ:��h��e��ޝBl��P�� ~�em!��߶�l���� C(���ʤd	mm�V���;<"���jU���J��lM⏶w�<t���^%"D��`R�Ӓ�pn���NQ�� :F���
�ST��M�Z$B+ ���MaR����pb+46vlC�*����V�r��Y"mU�Im0�ų;})�-�f@JS�y	�z��E� ��y�l�&�!��BK����>Y�[V�2�V�Ci��/�'g��+3y�g��P�����B�?#�!�c�0l�iC�A��0�+�nȮ��v�nu�B���y�SD���u0�Y.�D($ŰZ%���,��U̙�x�ʎm�Ԙ\����l�Z4ѪLѢB10H`'�aN:a%�c��5��M�U$-��]uTBR-&�U��-�'�!��Ӣ^Ԍ�֧=ӫ>��U�/76���k�_�,Q�rk�&Z��k�E �kҵ#נ|��A���>5����i����	��M:�*0�����]����n}�T�F `�v�u��A�z^s=*�Ο{�����g8e���(�1��p.̜D�ݸ��8zN@������iW��
x*RKR��s��?w{��o�~��Mʭ��ۓ�rv�&���5�Z�9�+�O_�_�G��+o���[�>n��~�ӡ�����"\���_�f�>㻯x����ѱgp_^�."_"{��o}e�.܋}�.�><��;~����׾����ϯ^�����<{���kO��3{���������KWlN<Oz�ng:Ծ�֦[�\����a<���W��;D�.��������/��&v����ʮ[��~���t�R����Wϟ}��/�_<��N�G����v�'W/�_]�??>���*�jg����=��(N��M'Zjaa�.���Z�mȓ�V�~�g�ov4�HN�!)4)*� ����q�#{�I�F�v��R�!r��#�LeY�ri0�)�LR"�� 4��uN���U;��>p2�i�p�:��H��
YjH��Ü�,
����P
�D��'+`CY,�O�%�4�n�>��00E�.'� ����p}���o}�[.�r
� �
3�F�0fp֌"�Q3�9'�UbF6Q�*l�a��M�� �2A)�4O��H��05U`vCEaH�t9��`Ն]�	�l�0�뇇����*���چo��`���&m��ލ�~�N��.<xx�2��_����y0۵�_}��?�|{�j��;���L����O��g.Y��(���`unj[�<�J�<���e������ܘٳ�yʒh�Ul�h�`6�V�����r�ד��6�\�^5#7����n)�UG�l8K�Z+�f�����9�c`	x���n���D�?�\���E��	r�Ģ��UM`�3���N k[	C�)��q���"pnIK�AHb愩.O%��J�,ʟa�8!� ~F��`�?��JC��*Ѳ��h�V�:��j�9ˊ���r4�.[J �&W�0)��0<�~���>��۶�g/b��<y⌉�>�J��Z��D��h+N��!0���K�%{[�Kԛ��3�i��^ȕ��+��>JHl�����;�M9�D�9E�1��&�:UG��u�w0��Ua�d@��:���0����D�*ɲ �h�$Z�H�	�P�����x�0f�;Xh!Օȃ�a Q
6òx��S�p���y+SKfF�TG��I��J8����y*�E-�p
)�MC�l��� ,�[�Hl~�K���Lb�y¯q�`)��h���&�]�O~�c𧏧���e(��Q��Ԁ?��,��ڐ���{���Q�D�h=�����-'�! �S��R��0����-��M.�{6$B�4��cX�$�*�3<d�/ϖ}w�qt>��C2N�Y@k%�����U����iؤ�\��3J�A�a�:�8
�����͔�dE;�H�5��г� �Y�HJt���HE �p�e��[!bCz�r�COSn8%u��]����,�H�j�(!�f׉� �ّ�"�C ���q�&d��Fa�u�t�S�1�+�A`:R��/��7ǦY��M��Ƴ���l�^jAv4g������� ejANW�u^�e���D덓g�d��Rsճ9%e�O��y�qb&���W�B|~F{�6�H�8aꟇa�Ԙ5@�!�I �w>G+%*Ѫ3j	Lz�Br�)��X�0�K�O��*0������t�R���
�8s��^'�x��Ì���`<����Z�u�S
�h�ڋҐ��1Ң%�3da��r�){Qo�P?r���S��9%2��pO��un��Ȗ���dCFˉ�����`�H�H�@����l����I �آ����� �ݱ�/��%e��\?b�o�&e	I!<�@���+T.~Ww��DO�
���&��E%����U���C����ϳ�l�am��G��9�0�E�lk���z�e���`���r�`����҂�0 �T�0rZ:�O0)`�U�/�9���!-EY�Rv�,�!�V�����3'LYU����&JRj�-��s�B�1�H��A���n6���5��@�Cs�e��s��I`M��4�v�a���c�$a���� +T- Qs�]h����p�ɝrC��(a�0��<��[E�����wj<Hr������4��~UHx0�߽��y�(��	���5� ̀�0�0lF�+A"J���1b��
q�I�ͫa=s�z��S0���	Ij{�J��d��ð����N`Z�	���[%��!πa�x�2�l~�t�C��-E�
����� �_?�_�8E	�!-�ۍO�]�uu�[Oה\�R��g���tQv~��$����ˡ�qo�S`D9q�2L؝��ϓ����k
l��TM�G���o���'`w��5w'��%P~s����q��d���>��C����Z8���9�M�#O������VՅU�ԣ�뎩�����s��_������u��ھ0������c�.��B�R���M������������N֓���Zד�����w�r��[���5ux�����j}.��M���7�>�_��+�� �������<��/��y����6�~�ߞ�?<~��4M�w�|qu~��?q�����}N_�{u��Jon�����п����g���r���=#k��䦧e��㭾��zz�����6���ۦ�����A�`�9lw=`c7z��re��$څ������o|�w��;N�^}��g?�ٯ~�����w���/�?�d�;��M�]�]�������o^\���?w]��˿ q�����M�Q�0�1-�a[1�i��'	�N.�pr!˥���"ڤ���3�'�>���P��4p�1Ӥ�uΖkM��c�|�%#W������\ך\er'�uB�iU�'��.!rxQ��d�W���M�Y@��[+���([-��萔���&�C�������pY{/3/.B
���F���nj�7f�H�ˍY.��PH0[;kW��&ٜ���Ha�.��F�-�ĎN� 5�?���"s��q�h0���#l0���M�h`��MD4�fH��_�Z����VK0��ѽ��cϑo�<e��	�ӣ3g�u��ڗz�{Q?�{�'��O?�����O>��~��O�ק_<����Ͼx���ˋW/�}�퇏�/}�b���I���.;����G<�w/��wg܂Q[֒�a��/Z�t�պ�`fͰ�Z"��4�1�~�aKC�[7�@m[������C��������E�so��*�k�{<f�]5�&,zg��kVEхQ��*i�`��C��Sb+2���4sC20�MH��L�� %Z��iC΢�'�脆�D9U��V!ax�(��n30<��,NY�c���.���r6)�3 ������Is��0y��P�Vk����UZ�z���r4�Ɇ�Ub�WH!N��)�Ӛ�eo(jky������-˦�O��|���H���D̴Z������C��������:���R'�5��P��l���В�~T����ʑ&�3CFH):�ެ�q0�8�h����B��a� � $��eyG�''��+�����h��L3��pz�+�:�
����IS!��ބ�zcoy���9�� ���)+�tU�	�00�&xiܺ�+ѭSY�+��Ҷ�ţ=��a�Bc(-r�����ŉ��O���v�m*+�A��MqcCv���醙N������r1�g\>8}�����<'1)�����5O��:
��8�N�JqO�&e^HHTqllR��� �XnN�2� ����c�����B�%��]W��W�ca Z]i!��-��s�^J����I{@�±sr�.�X8X=���=�Fly�h��Y!�u�
C�M83j�&�c��p@�W�p\����`�Y
-Đ�`;�l���P�*��j��*{XTh#X͐^G�@�    IDAT0l��*�lY ���T����KW1��!�N-iL�*i!6XFE�8+�f`%�Z�T4!�_9�fD�QvY�FC�$0mX	6�:a���#B�!�3�� �"'�!�N6����,0b�Uڰ��ӰNxP�V~���ft�kCT	Τ!]���V�'<a#� ��0�<�`y�.~�1 !y�� �S�� �E�D����$�"�Ï�hT���"���]�a��[{�C��Du�U��EC� �i��8I�d�0���uCY�1oI���� 6����Ey�+�p��CDy��fmH:�a�hL�PH
*FpF�, EEk5�,'�<���Z���R�bc�L�M��G� U�41�  �W	�T���Ϩ:��x������,d�Iإ��_?�h�ghˢ �D�0�٬��$�[C�R�V�ְ��%���#*�mF��� �jp)���<��6Q~�����"���I�[v<q��g�ʁΩ�9�U�dl!`m�g4NQ~�r��r ��1�q�g�K�U|K[����z)��!NQ���;'O �4'�'�Pz�� �����UɓS
QR.��R��_�_� ��������a<�7��c4�0T�N`x"���-�π�E#d8�ͅfC�R�Ax*ڐ_z:�x����O��Ey�(�ry��+H�CրE+ݐ�BW<B$<Nl�GΣ.憐 �f3H-�&���9#dL��E�4)F��:@H�x�D�Y�Rf�X����D�x")�O��Dh�.7�1���'$��Bߟߤ�^���[���YW4i��au(�P��ȝ	�XC~CY餆'+�3���5<��9g)xZ[gǔa��&U�O�ڨ7�r#�纼����{�熄��nj� �3~�w`��z*6�'f�َ��,���4��,�M8��܆4�� P�I�� �U1��N� �ڠ|P�_=������%���v�Bփ��~�{q��C�����=�^�����׏p��xl��]�f���z���7+�l�/��Aq�\qw?o�WYDW��m�����ƿn���ۄ���#�N7���p��bo}������l�XY	�{i��YK��!q��D���v��>���y5�G��-��ͫW/>�:�>�ۿ�,���g�N�I==�|v��\??�AVwa_�}xp�q�~��vC��Dnݪ�{�.6�������v{��M�=k|�wbN��$^^�_��^:�*&��N��?�_�Q؇���8�>�ðy����'G�'|��;o]�|�����_��+��7��t=�z|��驻�O��z��������g��+���Z˵1[@����
Y%!+�Ɍ�M�' m��gء��0 � �$<�j�OΨ0�o��	A��Ή����6H"
�l _�uP�2�4����q7��$C�.ٹf���B�k5�~����������!$ZYJ��*����+�@�F"��B�#�&H�`�����eɵ������c�+w�\Z��?��"�=��aD5ICb��ȋ�c�i#NO�U=�H~�2���V�Vj-ɉ0N�J��Qz!�t�h!EEIEw���Ɔ4�l��Z1v��-�9v�� 	C'`f��Ks�X���u��<���݆[�`�Ht{�>���7�|p��/��>{�����7������?��߯/n���|zq�����ӗ_:��������wv�t��
�K�Ҁ3�k�N�kحA�V�>�]�I�R g�fg
�o�q�1�7��$�HO˲>�+K	~�8ڵtM�g�O�c�c��k���z��VË���)�������|8�¥p� �^y �Ͷ	s6UC< ��;r�e5����G�j��
��CN���c^��N1D޲�z��F�DH[)Z-m��#4d$l����\E¨b���&r���+3�h)H�A�嬴! 9�0���U�*�B��Q柖b��dfW7rE���6���_(N��Je�n��wk4fw9o������^T�|�jI���ƧS�t�?�я�z�pOH:rY5��������gx�����N"��@U-嶫�W�KE���0By-8+�V�ћ�t�ͮ�5I���!���hv1kLQ!�N� ����#єQ�R'����B�D)����.�fa�`�tr�$G+�Xa0%�t��MJ�&r�#�[�Փ���<Ds��Ɇy�V���w��g� ����$@l�-��D�,`��t�D�?(�dmW��-�ӣij�ag�VF��� ��� k�)�̣�*��iJ1d�=!�zx�eѡ�a��5���E:���BI�3��n��*1 I���'dY��9��4�>�	�P�����%�R2h�Di��.���MHVsl��ɵ��͚�t*����$B�h�����[C��?@lHHK�d�i^�Fg��҃a��(��8�y�-u�� Jho5�� '�%B��p;�y;��0[.g��H��a���b���9J	��X��Y:f<����E��?k�b&`#�I�w�a�IW��t+��D�ɓ��й�`X�Np��Ø~vHLl�/�O de��c�N�i�V��\�0�B�&1��()Z39�XXQ�*:Z3:4�,�n���5��y�D�M�������!ZҊ1bːRE:$��5�C�#T"�\0�jV�@�&�p��D�0Hz��J��a�A���rɭ�!�l���8g�#�N2hL�S�<4{�u��D�)�=��D�&��h�B��J(T3<�Cbj�"6C26<9�`���>ٍ�
l�*j�r�d
q���M-%g%i�l����j�!d����<�H`��!L3�����Ia�Ix�Y�4�@%�X�H�]	Xu2�� D�у��?j�ǐ��Z
?O���xHQ��\� �K�	�����cmH��2b�x<%�z���=H���"�Z��j��[�k��g���*J�݆�Ħ��,�rq����6T��Sn�V>?|)Ug�a+�I��gD©�VrQܯ�.&$-W'�Ɋ�� Z�H�&CCZ�����$���4���٪�L�!N2NvTs�!9wg��G��D�ᜊ���U&I�	E8MeT"�E+%��![E�"�:<a��o.l���6�_o1+� ���FQ� b6���Bv��5���x���)�G���O��-J�0���4�n���;�i��8[@�f1l���!�ʀd7����G&f�D	:���y$H��YH�(�L���1��C� ��Q-�P�&��O~�Z9��&qus��Ӣ�n8Q�x3L�M6��9���G���3���,u���!�1ZI$�\Ѣ�$��֡?0�!��YN�y"6�1�ϰ�Ӑ�d����Yd�i��v� ~����'r���곕����>ڻ���0T����ޤ�yr��p��J�!a ��:@�#��k�ǰE�[�:�'�aE�x�
w�y''��m}����|=츝|������*�nAj@�&p�3��xݜ[�¼����v��=o��=�#��7�:6��el�)�߹~L�
���ɕ�,��#�9�Gסlv�s�n�l�n��ߜޞ�������_Oi����˫����ZX�XO�7D��#�{��wC��T飃��ˣ�uo���}΋o>|x�*σ�u;������O8�{
����o>~Ӊf�	=�>a��Z��ݨ����8�����݋�#o2d߷�Z�=��_���P�q^�.�c$wo�]��*�+ �~��������}����ɓ�~��<v��
�����|��������������Ż�����o���_}����qz`�a��g/�^����5}�_����ڢ���fQשl�J\}�����<��n��;A������_F�T��$��	.��ra���r{���$[�:9s��-ʃ$���=��lU��z��!���eF<B ��-qO�vq��Е�������:!�G}�_�<�%� r�Ѳ�kSH�Ƞn�_)�"�鰩��ƐL"� 攈�Q��Z����рӔ�M�7�zE�����L\
?��a�(��!��� �H~r=�RQQ��a����0��K�VH-6�Cl��<V���	�*��~8KA�6�aEE�.�t��*�F%D�mx��r�`���G��vD�/�O���N���tk��8~����r�||r�߿�䷿���������?����㳯|��Ggo��E��}��c��.Pcv9�ɧm�%��^u@�Z���N5�&��,L������d����mљ�C� 2,]��#�,���3��ļ��e�9��h������9}�r�Լ�T_�5�c˪v�
�L�d�r�ꀡE�Ot`X�����x}�L�l��1�/��y�/���dM8-d�*$�:�!W�
��`��*�:�'�$*�Z���9�����s���gY�zc�j(��ᐗ ��@m��j���&���Mʒ�u� b��36�P%b�[:pK��PT�`�ߥd˪��!��tњ�g&�!��kIޭ?��K�o�6�Iy�|���h�y��b�;S�9���oڊ6����o�����N��qg�^����ޞ���S�Z�6m�K�@�����/�B�E[1�*�f�f�����-���� �����Ӏ��tK*$K	)u�,pr��t��R**�!�F#
�0�uB c�
�O7G�\���xD�xTa��K��9�0x�T�c�*����D� !��֭!���j�$[T	6Cm��c�rc{_���^��aE�8o ��V�D�W��m��ر����?��d�k�e�Q�����U%U�bYF���nLs8A�CA�"�����
� �+����F��_$սj��o����ju��ʑ��9�k��欹���{ ~��;��l�����?D➽�l"������`gݙ�t�gGs����)=f:?�h~�E���W90Q�)jH���4d�)�*B���c<�!�(��0�� v���2����Q� ��.ud�ؽjC�������#3~��3`���BlX�QK`e�	d�B6UH4DR9�T"��vīHkO�d`ӑnOJa�L�z����+C��s�Hf�����tx�,�Sqӡ�ʰuP�)��0<r�f���DH6LF!�� u[;NR"#¡��4_�/����Hx�+O�a��r�9�el�Ճ!	ӂ���O��d�͂�O���l!�f(D;R����������d������Hx���!��r�yP��㯨(����#�zk5صa�_bF�e5�<��J�lR9!�l�ʩ>Q��Bl�8��F����YyT�q�!����N&�a�D"��KC���M�3�=�ï�q�I	�o�扐QE!v)�HZG�p6DR��?CJ��#�\��8�- ���L��0��Ԙauw�J��h}��C #Z��wdy*�(�G(��(DL��S�S+?��ѢB2�]�Y+��P����"�"<g[F�P�c
0S���:L��gl�$��pz@�S��:tL��m���n!k�,�������(	ɏv ��'�3�*2�i2���ɪ��V����R(��S���H�1�b�E��3?]{����	c�U%��AF� !�r�����\�#*7X�0���D��	��¨�h`�!�ު5x#X{�&'*�����t!N�\2�<��4;�9|~�z�_��y5�`u�Z�_:#��b���JF�`x�L�X���_�#3�б�U�Cr2 j;'��q�b�V�B���;��k[7H)������h���u*]ʆ]`uц���@7,�=��N.R�<I����Yg6B2�< [1v��y`��X��*��[��� Yuǥ(*��!�VJ;;������䡕�*����0?�����ܚiRl�_9vTR!	�&x�C2���<S�S:'��9�+���O!�Ї�nL���׎a�����٥��|f�){��|�h^&��4��X�S����(��y�Ha�
�߲���yA���1�  � �ИtC�C��s��_Κ߾v�n[�Y��G�v-ݹg������������M�c:��W���\�rd��Q��,<�%��?�^?3ysV���X,_��<�V�z�q�`���A���}uq�n�yxqq�\y�n�ý7��K.��(�Q�I��^���[�W�׾GV���2�X��C�#��q����W&�6�-7 /���΃�����ݳ�W/�N��O��޹��/����.���{Ӯ��}�kݮ�|�����Pwn׷��"Zg?��ʱ'!�2쭷�_�{�d���_jϲ�5�[����ǉͶ�y�����c*d���<��펯+���Y�آ���;���̳�'��~�΃7������އ�����'�?F�����x���|����^���/^��헯\<1Ҡ�ubǶ�$��ۜ<�]���;d� ����N%�Kd�ohJB$��B�0�=G	Jؐ#�'�a!C6Z�6?�� ��՗�khR��9F�ZaC�B,���gmqv���9�.�Jq�����k,H�s,`ڠ�҆�V��Ԙfh��R��t^VC)*� כ��G�r�F�P��>
�c���Ó��S�  J3x��2dA2�"a'ChV�<�0���fК�� 3:?�F�[�����)]T�!�7�0R�aIk ���W4{˸��n�D?Ûo�s n�9�oD��O���/_]\�ܲ]�{����_�ԉ��o|tr���WOO_>ٿ�xk�[��~��G��/h:i�>a�]pVڂ��{���G{�sX}સ���FKg�l23�Y�m�0�hӢ5qC+o5 �lSV�-�}ȶ����UK�0���������tz����o���d{�S�b�`�e�0�^Q�h��ep20�ϓ��$���C���8'� �� �Y��!�OxZeI�ya{GAe(e���8-q��QKuB���w�C�B�����U��V���6���Dc�����By�p��أ9�H����0�*���@�pV�'z�c�H�+x��y/0�8���H`�lh�y����[J����,�Bx [=��ǖ�˽�i=��B�
���,ZQ�̪j 9?��1�7x�<5i^���tQ�P~!�s��
� ��b��:��d�]0�ꂩn"qֿP;�Fn�OY�4{� lS�Ð���n(Q4��%�H0�T�Qore��Ͱ�'��2_�H�X]��`�Do<x�����B�<tT0� J���7`K�#�R��s�ΓͰ�i"�}ȶ�����٬}[���;��;��=��_o�������?���(ac�j^lo'^)6�����u@ٖ�6S���(�l�4�VL�6��O�� ��)���i�R����(*YU��* �5Ґ���X�P�	5�� �Նw6����������E
����9uLcTre9��-�ŉ�м�k��P'�%����r�Hhx �4?]�����p�-�6 ���-g#�'QE�f(���U��;@#v'mS��lQZ-�0�p��1��#�('p�j��;���r�#}��di�r$f��!�����hϠ!��n
:7�z�I��T%N`v<C^u:��6&K����aӢ���S!���	�O 	C���UfK���9!K@K���3,4N����yN+Vo0%N��&j��[~�!��G%�M��D�d0�<��P֖��9@��'tþ�"!!̨��13f}�i�(��C�@����
%��i�<���ɏ�6mH~���J�!lz�(���%�u���?�9gsA���+�~İ>y�j�l����GX�0y�#���p*����P)!�u������m���0;� �Zʹ ��=Ö~���y�e$R��a)<Đ��U~�-r��83j� �!���J�i~z�,�ٰ�6�]`�sC�0x���B�2j,C��ޛ��y��W`� �,d��1���S���i?C��B��J��p��R)���Z*W�x�V�;g�i@!�]fCQ�Hh��M-b(�;��-C32ddg�ah�Ґ���I �P��BQ��ΐ�����aԧD l�(]F�-2�lS�զ�Y-!Cv��R�1~â`��D���`(Pی�7� c�<B��th�lJq    IDAT�ͼD�����/�� ��5@�R���E��D�0����G�C�0�)�Ve�!p�#�y����aF�֟�I3��U����7��\%��e�$�B!
�w���'�I�$�	#M��Tnj�"�J�:aG>���H�cC�vN�$;�*�5�?!	mXiZVs/=* b��'��|0T�?Ð�0�P�qN4LE��Ms~)�K�ֆ��D!�Dg'��6>�Y4bXW ČbȂ�i!y|�g��9�����O~"�I�㑾+1��F�P�} ��jq��*^ $�l�&��K��(Z�4%��t�3??�"�t[�5-�趍�H�_��_�0�/c����u�m���nK�~�rݫ��B�ru����-��놩;���q8{��s��M=9�O��շ⦺u�����
��\���3�"炶{�'���N}/������[Mn�_7Vo�����涷iӟ��Rۃ�뾦۪Vբ���}�~�������.����}{~y�����>��y�7B�O����{yv�����v`-˕s��gg�}y���ux���9���.�ę���:u'T#���J7ZL�#�:�������SW0\�����O>�!�OW��}�����?�B���.��)�w�w��O���֭�{��mݗ���Ͽ�o?����g?���������x�ԁ�-�6�N4�k�L'B�! ���E�t �e��7/!)l�����p�q�0DXQ{��h<t�Y3t<�50��[d!N̅³��V�y Z��P�:�=�^�<��*�����^������S��3�S�.���"!r�C�6k���HUo���`�!�\d���Xt8��g/��|3�k8�t��7%xl1�r�@��)�r���ڹy#6�!�  ,����	�!��Ll�K` ڒnT ���*�OC��<l�;C����ó�o�I�j��C�� ��pT��MzLԲ{������.��N@�n`Q��=�s��r�N�ٳ�Ǘȼs�����]=����??��w?�ѿ}���g�{�����_��׾rz~�������?���W:�v�M���}�El}�s�R�7����o��oy�@��[�ݣ<�ּ`L����d��!���� ��VB�y$V�Ͱ\^q�i�����0s�4�<���͍��*G�a�z��@�JN�M��W$@�����&��_���ӢBk��e��I�Ѣ�8��R9	�B��
q����P��P��XG�����>|h8�VЩ�D$�R�4O���hR�d����Fe�n�9��Yҡe �l)��V��+Z!F�篷�1W��s���*B�a��X�ґ0�KH����GV�ڶe-������_m��:��Ҧ�ܡ4T�k�����o�Ʃ�,[�_�**��Ў��m�9����=�L:�[���f�BZm"�p�m�l3SxT���
�=�U���aӴ�U%<]�y�B$�M����D�͐�n��#�Z��.˰�����D��EjF�k�x ي�8�h{Q{� �*�6r��3kY��� �j��� ���z��U��bN�ij*Ʀ
$Ns�f����J��(�n���Bv���~_��������:�)��{��o�;@B�Ɣv��=9�����)
C8�ad��!r���I\<`u���uL�dӢ<x6��CN��Lӧ��fe�-�1���a3�DC�����3���О�53�8nN��cZ�Ceh.��tn���W LE-`o�B<��e�p:����-O�ωv<lT����diOT`��`�H�́f��D��X��\h)���!+6)�B�B������P
��9�S.d�<6��B��i�a�\n�Ox�%�l�j�0t!�!�,C���z���2��Yɯ���M � lH�8�-o56�3F��a�6O�Z҆Ή�]<��hF%D�l��p4Y�y&�Ӑ?8;��!M
uX�1��x���{��0Y3k��&ِl���n�չ���qʝ![4*�ptF�r�D	j�w�l"�0�B��:��*`��7��,g!�p�z"H�H��xl*m0�D��lx��"`�P��B���C!�Hx��[�O��4O0x��9[�` &�I�(��&�����o�0 �R�-�F5,�rH�����gYZ�AJgs�i(����C��*5��C�?E��RV���Bl� ��)��r� �����wsR��nRq��SJ2~C�O+
�������D���<��ӿ(;@��]ɯwl�b�f׹m �L�Ң�W:-kc�v�"1#m���*F��~&�'�a��vRc�(�G�r5-&�h�5�Bt̲zE�������Ib㌜S.Iuk{���n� @@��kH����S�!�T�m�a+7$gs,�~���hI���H�q��Y
]VF��^��`1�$�6˚wC"��aO)Q�{-�P�A+���^3��5�FUV �dJ��P���0��&*@�����5G����0iQ!T3d�Ѕ�$�Y���DkF
a�5�����{e���3���L�D"qw�	�{���8y*7���0�-��J���½@�2lv�j�`H`�"!�B<UW��hQ��0�%��m�Q�g��=Y��tU0s�-Ѽʪ��jq��)�0\MllRB�J�,g�tm2䌪h��	���H�8H��<q�a��䒮b��L���ه�
O�2D�?O���8��PSNb)�v�h{�i���C�kUz!$�W�Od͎��)Z9�q��a[���ͼ�.�7��5��N[h�a`ޜ���v�۞�\Wu�'�`������ݸ�Ĵ����#�5�>�G8�.�n���'(�}�+̩������E�__����M���%��x�+a������=:yu�����ܯT��� �_�\T�z&nh����<{���=�����W����nC^�����G��:<�zqq�����=�Sv�{��o�==>߿4�'�|�����Ϯ��煷�����C3������mog��erOpjã�{���SOr���H$Y6������ud��X�KȤ\rG��s����໾\�t���>�4�#i�|�WH_i������y��ؗ�^��,wT�"��g~����������K˹��!����ĺL�%�Gxu;���������
��v��Z|�;F0B��)MyI�Iϣ�,4@�f��td�`���50�z+�Y�����0`��-`)��N���y~��G��kM0N�s�㰺��+�|��'�$�X����.�(��"i����B���dk�ZlǗtI�R]݊��9��z>OE���)h���3ͱ��Q��PQbH6���*���Ȗ���&aD�dہ������b�$2Z��1�Jģ��aú���%�!�6�h� t���ă�04)!�d�O9^ˆ���羬���w��現x����n+�'!~I��[oܻ{��<�xy|{�� ����b��������{筗ϟ�>��������������/n��O_�8��n�yL�_��W�L��c�hCH?��D�}�s�pv%�_��D��y��4BH)�mH�����[%����[+Z���j	@EkR-��Bb`����e�<N�|�2z=�t���KL{�*���G%��B�<�I���>8��kn�ߖ�<l~��' �(�5�zl4~�^�5V��10Nx<��Ɔ�h��N�����0�ZM�J�)m�Q���Kڍ懩���5/�r#��e1D�lx")�� ��8�`���W��3夳�j�Gī�ޡ�(!gO�½C`N�O��Iɵ����w��xB����n�9:�u�6�8�:�c଱����
u$2h E�mG����&K�#�z���h^Mnܚ�&e�� ��Abf`���+�)�.�q���lc��x��<M�U���{��Ҙ��Sa�����IYRf]3�N=�O'Qm���LW����V�y����x��7/�f�D"c��Bb#��G
��Uo�0M�ӝf4mͰ��P$�N�����ԡ�Q�+0H�E�@�Ηh����@����O�2�We�(%yb�d��z�w�
�#N�j�z��& &�=b8:��BI)<`�4<-Z�;@̆Q1x��,|Y�PuC��V���Eɴ4� �
��Ǭ��y���Z���_����o�~�ҁ9 a[L��T����aвL*��*�	�	����F�):�x� ��920p�1�ؕS�3gȩ(w��S���o)`�N����1+�-)��]����S�δr5�J!��$'BF�,"��\��m"t��Ŷbc3�5������+rC�t�]���M��`r��6�E���>�hu�!��%j#��<��X=KV�6�5����V�MJQ(f��g��Y9N�ޛtS�S]6�!�P�E@��i� |�Zb���2�LDeUH�(�I�0c��!g�����y���a͂V
';��u�	 a�G��9���pJ/�6�Y4���a)e�@�jD['`�]@�<B��!~$t�]B�0�0ԉ]����d� +Tn$��*��6	V�Hڙ�m*�R` ���B`$���	�6,��l߲K/S�a��0�ah�Jӽ~sB�/9�N��̐�ԉU��<J�dOE�G�Y{�(-4H��5�0��S�� B�3 j&���hX����v�L���n��T�&:�`DiR�����X���k"1�D��!w�a��3Z��.�,�6$��%�sK ;f6�)�L�ą���2����x��!��h�%R���e�gL
��s��^)#Q��K5Na��ܐF�I�ʐU�!�G]�d�28E��[6���	�$�d�R<��l��f�A�b��T���n�����\�::�X���R������|K~ 0Z2��-�ؓ�\60�����)����#7�4����Vzr�^��3��>ws������*�֊&$�r<�5ƨ��z�F�͉-� ���9`�)�O����Va)̅h+�hT 3d�@M�1̻mΦ *D�Ԙ(1�DC �g�V�e��k��a �9�p�E�RJ�����0C��#�I�����U�di��c�O���7>|���E�U�0�	O���nq��?��	*�sb���CvM�<�k����OF�Jl�A9��%D�E#�˓�͙�1���r�hWjò�7������}侠?�nv��NڛS�j�w0�U܉��Y^��f:>��G���'�?&���NZ��c�����P�ۓ���}��T`Ѭ��}s���f�y���/�~:ӟ�ۋ���������Wg��G
y�S�W����g��I�m��fj=�sۍ�ׯ�������յ�8��p����Ş���?��g�{w�_��z��\��8w���`��z����Kw4=z�������
܋�u)�s�ޚ���do)��v=����]a}�-9rvm��<�x��Z��s�����0G
���0ڑu��1�D�cO�����?��?����'��~�Ǉ���?��k_{�R���_�8{~���[w�#_��-�Ó���q�����G���.�z���:�'�>|�u u5�f���_ڙ<�γ�BN:<m.慧y��*e`<d ���_K����T����3ZOXl�0�0�V2�u�H,P��0y�x��Z�:���u�*�&�
mO�j�d��o��gp���.d�m ̪�����`�����M�B\'�\|��_W@9�F�2V�Z2k!E�k�4I�@~��0)�s4M\� LCF6�B�D(�Ѳ����L
�bٮG�;�ը:X�8y`�ԕ[�(�`��ƞVٜ���t��p��-�T��&
M{�nB�t����p��13u��A?y��p��ɝ��~����=������y�����zw���_�����_=��������~�����޳W/�>x�g?��g��p�}��?��Sf�������߻R�FRWol�h�{"m�k�4�虘Q���~��LpVǈg�CE;L6A�4B���*��E�4����_��_BJ1;+i���Ӗdt�$��T��:�2��8a�LC$�<���<l�2j����&`��#
3�5��==�qJi&��U+���E�î�V�!�O,�R�k�������O)�RQ�8K�Z-T�Wt&�HZ�4�-v�	�9OY����������CE���]?��D�0|F�U����	ϣ���s�ǍI���G�|�Tk�2'qGZMb�h���������zS�����ˉ��n�h�K����n��Ua '�^�<�p��h�a�����b��>5�h�C��;�*���,����n����`  �;:� ��4�/�& ���,Z�h�
��|x��Y���l<Y��'@����!0??ij�ل��p(a��at�˖#��i�ï\"�*�DW��m�͎�eQ�p�[��>�Z<�%K���SQ׌VM�8�V��Cǝn�d�hF��!]>�}�����OS*zwA���?��w�8/��I��9��� �z�O����+H]/0���ͮ���B��6��9�%r���C4*,�֡�D]��1�@�IY9�h� 4�VU�����Q�@�`���4��EVÿ~h5 �[�	AJ��OC�1��+�LQ�*��4,��.T�Љ;��&R�l~x��(��}�[�t� ��� X	�SR!}B�0]�ք�!�ހiu+�_$��0;wՒ&��j����$,E?������jF8�&n�?�:��6��C[��U�h!��8�5TZ�*"�6&1C�0�㙨D+3-U��2Ț�D]������l������C��I`� d�ss��bQ�0���Г�n�9ͅhi��篟��I~3���su�z���5�0�0U�����	�\�D��aT�$�!��DTl-��3����3[J�d�gB����d�&���rI����	��v,��m)�����m.9Cʭ����I���� �����~j8{Z ʟ�16����3��Vb)��k)�4���B��Ν�r�Pv�*y������U!Κ�� KI�����a1[�E��<��#��/=N����n��dӤ�� �A����)CVζ�%NKu.����jЕ�%d�I��f)Y�*t�q�Sn+��0�h	�,�״���eQ�� �lR�ri!��a�;�S��V�oH�+�����<00ZՀ�<H�a��>��⤫<�v�%X<�'��`�� �0�D�b��aF�1Ȅ4iH�<�F�M��D��	|�"��°aT��rr�B[c�5)�-�[}r�����O� ��[d<3T�S�<[Ƣm��%Q��jXn�ɕ�(0?�d�ϙ�o)Ã��&��ٲ��3�hp���&�#�[դ CϞܐ�-4G6'B�8i��Cŉ��b�0|6YMS)��Ҝk&�.e�F����>[��43����O~C<���PC���	\�`��3�!�Ӥ��g�g���aȢ�����DW��Hsa�ͼ���1�Vt�h�8	g�h�l�8�՞� a0 �l�<�<vs9�(�'�ed#6H$B2p�N�v��f`��@V4���m60�YV���a�?��SC[|$)�SKֳf>V�qJq߈90��><��6��0 ��+��)��۲8�RW��ya(��cȨ\!��-@�/1�\6�a]�b���r�w�܆�Vu�m� zd�ҝI��y#��o�=��F������<{���5�ʫ��I�̼9�m��E�-�V�]�*��^��\?�yu��)}K+'�Uk��[�v?�廾u��ء�e��nC:k=��T��3�ދ�;#���*��fЋkہg�[��kQ�x���-�Rzrԗy�Q�Ǐ�ﻉyk��<�88<����;���V��_qq�}7�|v��?�|���=�8�>;��!̳�ۇ'�0�ֺ�N|����D�/�.�d��þ2w�����~Z�Yo��j/�X&N{�0|�Y�%�����:�~A����w^\��~�������q�ܭ��ȝ/v�����{o޿s��w�;������������y!��˞])[c�I�u���y�͙���1�q    IDATۜc3&���a;W /�!�#��%���D�!�Beǩ"����j,=-��\������0���*�4d�)����r�Br;�``�N�� �����Ŗ�}9�~���H%��W�������_v�����]<v����bӑ(d��!*Z���&�E��PS�g�3U�f$j�V�&Ma����P6*C�(1T��j��I���B�'d�iH)�n#[����O�-4C�i�3h�@L	!6?c��c���	\�Qp༅���w�����ǝo<�����ν7��]��|������Ǐ�x�tx����O��?��8~��O���gW��I�����G/��9~��������e��ږ�s�I�"����Ӟݢ �m@�nё������KӡI+F�4#|�� M+��^[�R��Ն(���m�b�������?��?1��S9��rXߚ�c/'s��E���j�!��Š-�-G��q4d�%���0h~����� M��YWM��������Ƞ��%b�$l�e1��9m���}��G�qRf���Dn��
m�nsɮV���@?�=�!�J�����ɕ-��xr� ��g 3�ch���C�S�Bl)B����+�l�v2;�+�K���i�;��o���2lM/!ڶƦ��:�w����j�d���'6q�P�Y�6t��1e��Q����0�|�������N�'��&�MK�l`Z�Wßl���Z�� ������E#�Y{4�C��w;؀�F���G�5��&���'Ω(1�Z��� ��81tt 9���)����J���I���B��݀y�:gT�A󨎖��3Zڐ�sC`�+�_۵$��cdc�x�\�̀����
�6����~��k��+�aoB�n�y�P�,`S����_Ȟ�䱱����{�`h�kFj�Y-H�>�� 6ß/ J�P��m�[��>�45Q`��4k��QY�1H$��G�����Vy� �cY�(]��N`�O��l2��28��F"򦦙j�ĺ�	�Sc�^�Ba��x`�H�H*m�;�ͤ0��Vӯ_�H�	N���̖V�*[�R [ٛ��U7Y!���K4�v�D1�i"���**����;�Ia�*�9g�aP�)ثʅ���%��b�����~0����/
V�&�O�k��3h=1h6)%@v��f Z"+���lE��Ӱ��#1�`�Թ(��xjl�B�?1Dk�&��j�  è7� �X3�R�9M�d1DK�[��f`���D����@��P�Z��Ee��h�u"y��u&�!�
��S��ьD�Y��r� �bg���YH
O���	�mN�Ƃn�`R�_t���l��?)ǯZRE�<�S:�J
U���hYi�
,?ͩ���6���Jݲ �R=�ˊ��&��x��9g"�1�0T���H�X�M�O��3)ͅ'�x�Vi~x`�s���r�vr�ZZz:L'���9i�+�Qi���-H���J��=����z��&�)��ΐST.?|�y��B�J[-3-R�솢٢:����Q����]
N!)�3�E� �������L���ъ
ykF�!�<E�y��78O��4<0[H��x�����Ϧ�%f��p
Clt���<9i�p���sTV���(�Ubj����͋�&q2��3�7��@c3���E͠�9�i& '�&�`�&�h��Ǧ����wds� ��6h�I� ͢(-K(|G?]3R�a`�E�`�uȃ'�0�$��uRK��hΎ��<%�gh�x0R��u	�� ��`�	���XgCNC`M���K	�[��y��=���Jd����`�E�ϰi�s�`O9M�N:CJT�Yl�-~�D������i�(q�ܶ�*�+C!v�˟��Q��
!2�'�40��d�Q��t6C�i�%*1'�Nꓧr�8g�`13�?�n�B��I���؊f+�'f��0d��0�d����Ea�:�,�'h[���ƹ�_)�8�C���%>הd���!>θT
�gC$�{��|�^GZ���}��Qi�S.<�7K�!��$�R!F���!?f!>^�<~~}p�	B4����5��oW��\��^_��#����\���^\n7o]\ٟ��JY��w'0�}ӡ���{���y��j�8��/=�x*p�W���'0�mfjF�ח>mzR��Բ{W�G����n��T����z*�c�
���������_�H�o��8<��?�G�w�������}_���������G��Gw�O��_�?�{�����'�����[�/>�����ww��O_ݽ�Ļ���\�.�tl��N��|��\wN}��GV�%u��:��;�?�<�cvۖ8_-{�sߝTk��Ŷ�Ҷ��8�kF��]�C�9}��l��>:��I��}�o����������yہx��Ͼ8���յy~Aԓ[w�q���=�;O�Myxp{}�w�{z�ʥ�v�%W��eӪ�h��z��C�vr[^�ް7�� �:��V�6$��l)����J�vi!Y
��C0�)�V'Zu�8�!��f�j1x��!M&E��bKO��D�^�����W-��Í���v�2`���N5���l)�8K�-���n+)jH:gr"�S?��Sch�@9��m���$�h�i��c㯐D�����0ԡ��49Q�� ?��	�Y�j�`�̰bR��0�1$!i�t��CX.?B���=!�DT"6א����}q�����[��x�7~�}��}����g/=��'{��^<����'G{������ǟ��������:{����ˣ�|��茶<:y㝯���~�uD�\�;ܿ���?��Oj#�^�ݳ�4�%�?��y\���c��ק�� �K������H�T+�,�4��Q�el� ��$;Ł���xn�����-��O?U�����t�M��$�J����Ç|��9p�:/M%1�"ML=Ŷ�V���:` ���BM�S�<mq6�ui!TaHa ��b[֪��3C����L�?0?�6��ʁE��6 ��[C��x;𢎢��d��DvHiH�L7Tw<�4@m���k�<��k8p����&�VCzj10�)' NF�Mp8�Q�B��r']�.��6��	�FU<��������}�	����� rl�=	7o�O��ٟ�m۸������K��wtQ/K��j�00��z`(Q���g�c�VްƤ 2xFlN;D����ِ1s:}ԕ���s�A�����H'�8�H$ �r��W�? ���9���L��h��Z�G����`��g0Q"d�*'1ZF)SKo�3*�7�Hfj�P"01}NY���!fS���x-;����,f���]���;:B�!��tT�SZ���ܬ���󩝬��a��4-��qzE��e}鄡w[�[/�&k6�$M�+5�����������O�T�����o������ꟳ�� M̮c�C`��o^~`�b ���.$�*L2��̮�a�aJg7�\�r�QM��C�8��Y'�B���%�2���H[Fx��P7���V"�fh"ت�Z����UHz�aC�� ��/%??;i����EH����IN�:1�8ͺ�*M�CJ����$������t�O"�0jƟ�Q�_�����8[��ˮ��q�_3��j8�=k�b����D��1�؂�NC��������V��`	L$�:	FGE�,]Q��N!0ZB�#a�U��J�jI,ʙ����	c0m�A9f��+���7Z$:!���l��am|7/�V�S�aF��T�ea��|�O
�hY[k7��
��"��9�m)CvD ��dT�V6d0ƴ�0,jYؑ�d�7#F$�]���\ʥ[^0����Y�--e�k�j�Tg��� ���;֜qV8�(<A����2xt�������+5?��ۀ*� �ϖ�P���Ş���0�tz����\�sB��muy c�)K�MUjO9��MV+���S�|1×?rY�	L�z�0��E�R8#�"'��b`p6�ͽ�B�����NpXK���tlS��:��<5��X'��0Q�C��Q9v)2[�tZ�.�N`� ?q�E(�(*1'L�0�86Yt�h���!#�ݢ9��(�,�i�i���DH� <�sCM 1��D~�t���Bo2â|�0x*��&�İ�w�j�,+EE;�M�ΎafdH��f� FU�Z2̳��n���k�P��~3���LŐ35�V@4�Y���j���(�aL7�f�&񔕧ҵ!=NR��STVC�Y0��.1{r�:�(Z$4���f��\0��T���qn7$��bfFH��(�I
G��_�� �0��UF�t�J���g�4�%D�h���0�����,=�$���xj�&#�4L�`DU
���iFbX0�dp�hy�%YD?y�0Is�+�� ���FHe�N] )��`��ۇb�!}����3<���_�4 ��P��s@}f�,=g�����( !�ڎ�B������H�O^l��4ku1�&��ӆD <<����]HV�ώ����ز\M��q�7`ܹN�<�O��P��>UO#^�;禢���pCq=��a�#�_�z׭���,��w���8������+_���-�i�^�IO��ug��NG�C�k/i��t���<:X�E}]��
���*}��֩{�.7����'w�k�ѱ66�����`]7c�e��Uv��T�.��>�ZY����c7S}�����۴�'w�}���g��G��u|����˵4Ww�z=<�� 遻���4�'v��*y-n/X�n�m��*ߕ��yV���_�ɥ���������{}�ś_�o��Q �c/9���Y�L�6���&���y�f�s�~�{p��g���֝[��^<�������8��/_]��?~��A�8|�p�#���x���~�<x����]3р��4[A��E���h�3H�%bó�a��%�T��m�f��a�X{ް5��0@)5&�d9$]�&QJ����- ?�qt0�p�ِ��	�h=Kg�aZY�w��3@'���0���Dm�dՋb&��͑���I 0d�H�+W� �#����F��V����b�x�Ig3��(Z�~�u3���㚅t�0��È��t������j�����P�a�y��4S�r��͂A��p༕���.]=7ON�e���Տ�����m�~��X���پ'�/��^��2��{�ί�>~�p���g����_��g��ֿ�s����;{�Wٯ^>u��@opf��^�{+�7Pר�Cq6�>�����K�&�2'�4d��L�j4�m�k���M��,T�,���M@�` �7��9���gH!� �I��r������k� ��;�z���0XH!���Um�M�|8E����Sߢ�E�Zbݜaf%��<�+'�)Ti<ZToHD�%*�Ϟa$�V���˷��m+#jAZ��%b�����P�N84��<����
�7��3vu�t��\���4@?'v!xRۢ�x��r��I�E�U$ ` ����NlQ�_�[��o}˪�ޅx`�hI���D���'��hn˺����(i�73�
����� �S�▷&�=`C����ѧ�0�m���@� ��וm)j�m�2l�� <x���0Dː�0��l�GO�H<��"Q��[�=�!a{j2 '��VEh��Џa0�%2୆ea���%�[n�Hl�'� ���;�i'�N$bCE��V��x��U������(�]�Y���`�$M��Ħ�\!<��D
Նl�t��δ�RL��i���w(����:ԡҪ�@=��#�m���ȵ�+ Q�Ho}豋�z q�-)1���KZ`6��A.���c����Ϧ3�2���iex�4�ĢV��Ǒ����%��]�߱pr��-��rN,�KM:�Ud���m~�iv�;(���>�e���ak�<`��K�$L8�:4�NnN��c 1k��ijr���Z�礽ٷU�x�;'<<��ج�?&�IR�R,�}��D~Ȳ����:� ��ó#lY��_
��,ҢC������TBO:���.OCxE?0Q+��p�s:0g����D�aRŲ`33�2�6���t�W7� �p�<`l%���a�>MI!����uR	N�QeΦaD��1x�6�T���x=#��sJ�O�hQ��MJ	�g����2��-[z0�a=��K�):��DT(L��I!�N�Ӑ�>�5��޲�����l� �U��c������ [�!���zH�i�sJ�V�`4��i{��aYi`E�I�b�ώ�D�zȈ��Ad �l��N���	���,�o�7�[�r�W���x`0����i^t=0��a&��@V�q�7�_�es����aW+���u�� ��U�e���ac!� �`ͅ��d�Z2#!��ZmL����8�ɪ�2����6lń�f�\x����Tg�U�Z�O�JK�:#�!��&^����7��a��Q' ��՚���8��'���r��e�有ۭ�C�O��T�hUg����;w$�-1N���#�$�F�;伲�h����4���ʹ��Uo�	F�������-
#D<5c�Vb)�UL�D^.8�4$�kRgl�jI�Ynl4��{�P!�+�J��2n�T�ʖU:� J[�H4�u
�*�Y�|���;�x¨[�ֳ&k�-���� ?m8� �pf���38�y̮"=��b~���P%�&����4@F���yoz�'$�Y�HD	O�EyFLzG���8��ǆx�����a&�P&�!������ʪ+W&}��ل�g��`)������Iǧ'�|�A�����>�w��]�����0��un�L'����j���5�� HT��Va�-�Z%�t���\����Od��Z���[��+b�S_���N%c���'׮��N�۹k5��I�n�6�jF�~��s��v������l�Ozj����mK{D�o���&�7����=r�pMb}O�����\S�����-��L1��"�������,t3�×�#����.�/�5��p�es\Ϥ�N}W��5��g�].�W��qW�������o^_�T���[������]i�w}S�W�O�>��~����W�?}�?/._]]\�ܻ�-�� ��V����5��������k������f�i��+�<U���v�������UC��6p��?����>�;�k���Tr���~���z��ûo�q+��m׮���������Z]w/]�{������w/O�����??~n~Ǟd�s�k����������o_��Jx�Q���Y�<�E�	1��mk-���gj"�lXʤ�� ģt�FgLn0��4�܉�CÚaG"�[}·�Ҕy�4̈�K�	����EJ��r)09���W:���!�FR0ai�s]�.x��1 �$�B�i���AxJD>sfX] ���R���R�S�,0b�4,TQ`ÄMT��ڷ�/�Os�6�s0yh)�V��U`KϠa��̮��I�$=�:eHAE�%�!��w�o��Os<��4���]ow�o|�������O��9?�z��g��~v�|������z�����{�O��ƛo?zv�u�/&<p�_w=�����z��������s�����-ɛ�-ԵA͸GCzOѭ��|zs��>�c�8fd.�&�3�m�9۟����DJ���k�;����`H4��iUo��(}��.�z���O���y�T�Z8]]?t�ӗ�rI����4����� �f����"-28f���Yߚ� c4C�Q��y��z�(�O r2��f��f��q2#$��'@݆��t -���I
�@�1HlYx���*��dh��08i)e�3rJ��.��\��Q�BR�m��?��0�� �$Q�aZ(�8y�)�Λή��HlUmo�~8О�z��M��Ul�ڑ]Xn��*g�mE�!亩�����:�O	>��#����Օr�]J5bS��]{u�"7�B���+���bng�u׊a��B013����@�4��+�~^&E[L�h	 �BzcK7̀�f %3��xD(�,Y|�    IDAT$�>�3TN`m���A��^�<����dٲ�t�� Lum���V�6x:7A�nc�� ��ɖ�/���p�4L~��ʅi�LۢB���(6G�!Dc�a8����ZJ
<0N�E!� �
���)��^ }Z;�w�w��~�;���_��_cS�����'M����J o��J$Jx�Z'p Φ�S���Tc�M��&��qB�;
��NLbR�)�Iğ'����r�Q	ᩜ���u����Kd�i�,K�ާy�C�B!�� �t8��˶�
�#�٤��`���ј�8�������'N~��d�2��ڮ<`�	N<�55ui� *g��[�cQ�����HT�e�����au5@dсq2b�GED�&�,c���k�0l�x���H*Jg�&%=���$�[C=D^����l�Q!C������nTz��O$�D���ĥw��vz  ��f�O~�<�uH7M~ Ȫ�3v;�1�,�`t�t��A�yx�{@ݖ(��#��&<�j��g��5�{D՛l����\�����r<5�A'��$����3��ߐv4��ɖ�����Q�)�������1�Pb�D�H]AF;Y��.�D������I�<��$[��d[VN�`e�u�i=�)!e���5 ��a�I���$#�r�ц	/J�70�=���� ��H�hi�J�3�R����̂�sA����H�gďs��)W	Y�8�R�WAk۰ƆP��<���9��g�3�!;Z�$�R0�g�-$� sZ�\<f�@����Is��Ӣ�[��P��6��B��%S��K��!�g`):D��(##
�?+6�,Q2� 5P��	'�Ϛ��8�:����|7�_�g�SJ!�Z
"����B��
6)��Č�8;�<B4B��>�0|C��'<��1$� �i����w��E�b���Ӑ�̐�[K��)�FeXK���~mNs���ͨ�d�M?l!CTll� 7� q������p<9���hs�$j����Z�YڨۘEK���RT4���0pӇl�{��������R)1��y��>�a���[a!���P�03
�*mF1 3I%�Rt�?<�YK�-�+�i*�L'U/�D�l2Kں���fr��+�-���=Λn^��� 8è%TBͨ?̄⇇i%a�!�5����(��B�tFEg� �$��kX'>5��̧?��|)���O�1��I��B�}G^ŭ��fLv/O�SW*C<��o<���lyk��;�({ T�	�!�!����fm�a!�>E�9^��e��o<2��`�!9pq�ϕ�4<�8���Z�X<~�5�Ʀ���_�H�P�=���KF��/�f�<���C=���z2�����+7��w���&�6��:�{��{�����(9�~Ww�)Q>Ql���/�.օ�_�������;k�-;�=}�i�S�JJ%�n���3�̊�[���`���to"��D )��FĎ�~s��6�&��9|�p�s��v�^g���ۖ���Cq}��=l�W���o#\!�|Ga�?��Vu=/pyw��[������o�~�oW'���]���F��/������������S�����2;9=Z��_�<�?|��7����E����h���*�������?x�j��Q��Zj���׎l�:����E��g;�D��	V����7��o|��G�G�z������GG�̞^��`)N ����w�}���[��������9��S�G��8#�d�mKx8'U2�I4[j\MlV�1ȁH�N�E����C�G$�:AMe��D롱P�8ь��'���;���'˅���B�6� ��J�H̺%Njr�!`�h8����L�fbMk�k}
�[/��y`H
!�95�ɊR�=0�)�$h�eʝR�U�c*1�ғ2
�G�C
A�|�Dt�Nj�����r#2��B�����u�/dd���.����޳�0�h3�f��h�
��z\�����]v����w޺�<��x���u�����Ǿ\����ӷ�::۽z����o��_?y��w..|Š�7X_0�ڴ�ʩ���ۓ���i�du�؃7�јK����>g���D"�m�Bc����F#e�P)��M.��i￪��	��&Q�����O�ڛ���^8�|�I�m��:P��fJ�$L���,��H(L��qj�C�H�2j%~
FH#�Ia���t?J�tDԪjB�*�"R'%B8��\Q Zu��~B�����oܮ���.�JEÑ	V�,0�#_��hU�)dʐ�ӡ(?nJ�E0)n�����#��-�>'q��X �lNd���Y�#�\4:C�:w�l�:�nj��'?��~�t$�,�ѧ#%���c�������:G�N��f�Ҳ����z?RÉ(
tuPB�4;���ZQ͛�,�x�! /@п�%�VqD�l����@�P��[;�>��F�t� 1�����!l�� =��i�Z��Y'�0͵_oްѤ׿��N)Q�FA�(�\�p��@0�ʸ\�l�Z{�M۶��W��J���C�cu�L��(#)8�J�v]r��*�H��(��BL M��!0eR�J��o�s3	G�#��%ը+�7����w�PN]|/��:�束�T,P��Q�;�U�$�m�@+ŉ&E?�iBe�]�[�����+���R3���Ȥ @�b�aR��r�|),�Ry�X`�pjY�iMS���ц�8:rq��s�m,���:{�����	N!;c��|G��5���!���sU�3�|���Z=�ju�(wԐ��`�4~�tj�A�~�!-D�hR�u8NQ�ٶ(}����!���
�!���1�|�4�#��f�|`L41���r���1U��)H02���p��'�C'���q�D��@8z���W��J�oS0�i���+WV~ ��j����*G��N�+���Il&Rs�y-�� ��$rL#�q�}�LqX��3�R h�VO[W��
u}ű�B�S>�q�2{��|��j1Mg��V�U��U�O6���
δA���z�@=8�h��3S(&$��쌓�L3����Α��Z���#�͙��(��S��*�I�P0RÉV�3�
.¡/�!�؋(�ZY��/+�pH
���H|#�0���8�4FY|d�B-\�ˡ�Ҍ�:��H����qu���) :�BRBb=7�`�I6r��֔#�,�*l*�)�R�	�s��ȏ/7���1
i>�)#O!��FQ4��&�Bz��W�V�s��U4e)Ԁ��R091�U"���� �0�1��M�,*QT"������I߸kPHhګ�e�||����o��J�X���88�k� 
g8�Պ��4c���������&�pv%��Œ��9U�*-'}%��J�R��6Q��V$�r�KR Bʅ���1-}J�A��F4d�F�g�f��5"Ս��\�)�����߆�2bjB$�D���IL�D|`}� LH|�T1�c��of�vU��!%�2pr�Í��8�%B� d����*�+���j�ik��I�h��(�2;���k��%#p��R��g�C�DYd+4�zAf7�lD�P)���#�nL��t4�}�^�h	����1�{xR�f�E�@���8�8D��ƀr9U�'O�}0�$W�,nJ�VR
0YN�pF�q�B+h�C8�ğ�)4j�Z)V1��#��|�,��BR����p�0|�~�$D�,���6MT�(#b*��Qz��	Ʌ�1�,HW��>�A�O��W��c4�H���~�SE"˭����|M;y��.���e���̭��nu��ÑR.oV�'�\�z��d��:Qו������������7�*�6�Mw�������S������O���{}�;]�3bߧx{z�;��������7��}|w�z�v���ŷZ�L~��o�=�U��[���ֹIC�s��W����wg7'�O�x���/}3�;S��p�;?�E�����ٯs�z}�سg�|����������b|c��6�ʻ��z^�c��;y�:���������Ӥ��ږC���]�)�P��	z��[�en��2�������?x���׷������G�o?���O�O/l�œ�W��l��{�u�������7����ˆ_=���rT����9U�UT���>\~!LK�Ι����)�i�9j������6�E#��Ȕ�3��W(�^��J�Oʁ�����z`Ӷb.}�"PPE�:	�"*w.5p��҅��8+ �	'KM�)�.�&L3'2�������l��^3�Gk	5m�����͡@��2Հ�-��g4c�Bխ[!��~��mH�	���[�wIa!��I
��I!�1E�|�|�q���
�J�6�s�|�FjJc� ٵ��EB\��Ӑ����{ߤ}����W���������ի�_\�x���WnG�>�������/���̯n�������������~��o�^�������_����7ͨ�웮�wS[�w���BL�v�տh�#�����rp����,E�mj��R��-�2og>��t�&b�^y��3?n����sW|KAƁ�	�c�*�$��z ���*���!�Dmq�r����d�Z�XvLkCf�푬������n������i=��f�
������DU4ńP(��iEB����fs�}@�%���ˁP�d�LF!�C��
�eZ�!�e	���BKtkCnc��k%�1%2��Z�a�µ
!�8�˵-�˦��jg��
���tw�ǟ)�����6P���h�Թ�
#�+jm���w�w�z�\�<qS�+M-L8@�
9�;LE�2���[ʽ1���	��ǔ.��VgO�:��I?��5�VcB����% e�r��J�T���a�9E)�ɪ���)�K��(�*@N˗��(Z&Z���EViV��r��C F>D�h+�ͩU3hL�*&1��P�c��VE��&]�Z+5�V�Wb�h�\d��s$:��!L4Y��I�aE�
�D��l��A "��� T��h��Rsz{��A��/~���B�*��w�]�W��3'��G}��������*DLq��m�Q .Ŷ#�u�k)��yU���!�Jm2{�i�,!�QbL#��p�E!��|����4�O!4� �^�}����!R��	+�A#M�`Ĕ���3���M��eW�^8�G�&_T������Q#����Ϻr�A���*�N骤��\S�(?����ĩ"ݑ��w�㰺��W�DL���'�'�R VS�Eq:�lQdH)Va*��FH�b���F_�\%�L�ȢB���=���_e��؈��u���M��F A��%���J6<�>8�hF�Mom�)#�7��c��1E�bD�fk���X��~�|�T�jUTzu�rBQY�41������)�Q]nE!��d:EkOQS�����8�ʐJ8����@���Á�U��1Y:�䶷�*m����`V"qӖ-&�����@��Hv���FNn�j��H%����8@���G�M�l��1Jߘ�6�		�U~�L��O�)�3#l�=4�#�>�e
�9��s)p͘&U��`5F�S�ν�DN�8J(ǡ�lUf�IM-c�!��s�r"��q��6��Pb�p���M����%&'ec���B���*�T]�s�|6d4�����&�XH��fR[*o�Z�3�N��i�z�#nl��P�d�ͩ:)"|�_b!�h �#��DuG6N��t�m����l:��פLk��h��J(�8p}N:N�rfQ�z�<~
�f���b!����c$������-��8�y�1e#��I�NS
�#@����E�ES�����(�!��N
��Z'��J�;?B0�!F�d�D⅌���k-}:i&'eLYJW�DfH~�Ԍ�X	LN`%d!�t��!t��R���>�V:Y��:�ɖ;��,D����`2"�d�S"��h_V �\N�`K0v�ﯫꁢ	�ŧo�Z]�C,\k�h:]�k	B��sʉ�XJ�mWY��e�JU̗(�g]Ǆ*G�M�� �Z�h�U\{�\>�;�Z��U���8�q�q*!7��9Y�	B�~= S�7[M�9�8�3+�TZ�/}��A*'�r��Z����;���ԮJ,4��!�JG��J�bF�S+��ҝ~UA���Z5�#�(�C�Ħ%���' ~��K�_x��)���/�_}���s=���bo֏���:�>�u3�κ���x�1���ݑS��a�:Չu|҃b��[���ݵG#�x��D������߳��'ǻ����U�r}��o����~���ڰ��S�\��4���aJg��4��=9?�g;��o�^t�s��	uX|���zd�s�kQ��P��y�������һGK��]�������ӧ>/{|p��?������_����թ��6��?:?;9?pB�s�ۣ~��7�5+;ڝ����!n����u�؊��a���������q�ӟ��l��Z��댽��X�[�m_����� ;kyo^�zc[�k�W�g� ��Ջ�޽<]ߚ���x�>e�K�t���=>;w=:�w��l�N��u[�����/��[z_\��=R�Jtv�kl����g2Ef�Cج�c�h|Py��`g���.m����J�C��u>��L���T(�}Z"�V�DM%f�r�ZU�ִa�I�J�8pp/=H!�h^��BP�(%�f l��d��@j	��)G
��1����p��z3���~sm��A�`�N�-��/ǷLkѕD�P��m���)G�1M����pr�� ���� ��x�Eh�8��ɂ���a8��8�p~S��f6�e"�]5���E��.�N�>�s��%�.�}��o���|q|p~�{vs���}MO��ߺx���<M��?����={���_����G���گ��3��}�싗.�z?>zt|����r�|��ۨ#�oO,��M��^N�mQq�Ғ5�p|2�ĐNV�m'֙l�F $�׈�
y;�9���Y���S�"�%OItw�'�t|k������ �i9q�N%�^�P�kf�RR$|�#Q5Z�B�N�X�mSA�R	"�Y�o�&-���<!Y�"��02H#B�qW�]����(��}��!�vy����'�������NL���R"<)�p��AB�>K1��Հt=�!p��2p?ʟ����e��rL)�44��-��(�˙'݋֝�>� �}ugm���l�t�����+�6�n;�p6"(�����I�M#g3��R��X��BY>_�Y��Qm�C�I��R�w���T�S3�5U��8���2������b5#ʯ�?hQ
��,��\�th��JW%)�t>����B���ES�E�i�@R+d������b3�ki��#ZK9B��Z�,��\������;�@��N$�[��c�#H���d
�*Z����o����=�&�O��iQcY�p�2�_6�3Jq�Hw��rС����}��߆�dGV��(���Hу��W�N�+�}贬[dS:��\����޴����YM��o�5��̏`��U8�~E+'j!¨1S
BNHQcY4��ҶW��]޶����nu�ʞK�o���/�	J�S��<T]�t\S�Ѵ�Ն)G���a�[pX�:�+��1Yr1�T�rL�J;m%��Z]E��L���1qg5���Z:��(�ԭGW8�2��a�8`k/.�(ġ��A蠵�����g�hD'���W-��
�B��B�q�K>"�3Rh���i��L(�`��
BC�Q $Yө%űh�Ӻ8Cx��5�Z:�H��R�2�S�<�UJYpj��BӀ��"ǔ�('?����ҙƟZ8��'�(K�*�B��5}r���
��e��@�4F�����3��o�0�.,^G8�&U�J���n���Bgh�}H� �A�>!��J��,�h%�������}sѐޱ�Z~8|@V��B�8�~(3ӎ5�*�)2��Q�#�jh�p\O
)�0�2����08>NYp4�V�"�i�妜T)��dE��2!��45;@<����Iq��R��Y�˭���8l��G��cl@!S�=lj�r�H�U�&T�y�۩�O"��7_�x�Sk7�JL�n��f����    IDAT��0�X?@�* NWSQ)��ʹ�����h�T-��@�@��6�J�PT�#Bc`S�,�ܔ�BH-Y�F��[�!@��_�ь�C�L�ȍ�,>'���D&Ą����Ko�τ8e	��!&1!L�C(+��\S�P����@S>�a8?����TA��A"]�eq$rT�i"��ɒnJ'������p��9�|�6Uh�0�1S8B����s;.eK��1S&��F8`Q��6B�ě�~�@�&+���N�3��o:��I���$�8 N <�P��E�����B]�FHjF:�::��Vm�J"K��*R�Cz��"R�|Q>g�Yb��Ut���V$�?���������3
�'����DcNQx"N*~���Mo�]���LsNg?$Z�
Q.Z	~����fl�+�>�Յ��̙�hF8+��w���7V��t)�
�Z�vq���8μ[E���ٹ��@�R`M!tD�PQ?���̇����\���|���I��)�
�G맻U���m-���no��%��ܶi�q��]7ݱtOn�мs���#����>i_�ݼx���ur�H��m�L?�l_c{�/���k�,�H*�;?;|��#���{l����I�_���>ޮ���J�v�ѧ�}���n"��︧T]n=A�W��}tr~��pO�^���g=yzt�Q���Ɀ'���'���S������n����O�H��3J����۝��]Z���U���ח������*� �[�~κݝxb�����U�^�^�c3����9O� ~���}�ǘ�H�-m-ym���_}�O���o�ޓ���������g<o��_]ݜ��tSd��|;��ݷ�y����K��݄� �����������Ͽ��O}ʤ�]ݲ�4�j�J�}�.қkf��=�8��čYY�%�4���rX!%ʭ���`�g����rqʵ�^h���r�W���_4�����S��#�Ũ��W�i�&RB
A���k{yr���?<G���d�|�m���>�/�O��Bp��
e2���Lc��g]ߺ~�=)MpR�s��ad�jL3�Q!>�T!�pZDu~SQ�G�t�Q�̷��L��j�[�O|����#EtUb�1�H�Z��"�D D���qT��zj������u��|���ū��K��ę��,�����(��<�*�{�������^���~���=~�?��3_;�{�|�rw���-O���κ��п�˿$�Du�|R���[���C���p����o[8���*��>���XfQ�5�j�ҽj:I\��6.}��qv���m����?�裏Ⱥ��$sS����?���?���<5�^Z�$x#�[��E|%�j3�5	�HU��i��.��-��T.�(d��D8����� 98E%"3� ��Z%��7��}�QcQo�M�8��g����+�&s�Ɯ[ӤJ��fj!�q ���No��9Ǵ���%X9�NF��J��.�����H!R�@��9,�ȇ#�4�۷@�n�w/݉����?�VS	g�-eN��f)�������=��V����p�:�<�֭eG�Ɇ�b���}L�R���h*�Y= u���vI
D�2������GR4i-F��;�
Rm�)�>_T�F�����I!���px�+��K��I�ʅpJ	�V�(
'���0�
�t��(!�A�HdT�&j��B9�.UhJd�!�+�J�q���(M!NGm��Ԏ�	v��1}Sp��L�ZLe��[/k@ps�a�ӊ��u�TB�v@.[�DnN��%d���<w�tR��^;]��D0��=���u��=�uY9o6B�Y�����wM�v�vRTW���Co R�zeA�{�������7��[B�FY9�tQ�r�md�#�B�-�7Aȴ�ᧉ	�����Ίt�"b�j����!Y��B|[�[�D9�)�����\�D�*$G�n2���|`��:���|ˬ�t���	��BY/U��j��R�b값u��E4��M��b�0b�:QA-#��{��!��J�-o]�I�vĉ��pF!���C�׃����/�g�($}12SmsF��EVH"�ځ,�*��8!9|"�5�o�SSژ�1��T����i�T��{�Z�c�D�V���q"%�̤s L��(7����f*�`j�#f�	&�S�XQ%���v�?��_iS��d�Bb*1ӹ�Ț=Q����,����+%�s@2R|�l��@%�v��A�O�D+ʯ���C����w�G�d8@���?[D���@�bj�Z��Z� �2��R�V�(�T�	�!�����N�,��D8e�t�R�7q"��N�)�Lu!���7F&����i�&0�*�qV���VBV��Cf��s���E<ͪe���pФL9�C�Ȧ�>k��/Rݎl>~)9q�HQ�Ț�~�Ŕ��0�Dm����qݦ��5���1�V�a��!���R7֭,Qcg#N�)Ga�P�����2��X!�)ӕ�vt��Xj�čv���� �q�� 5�&�f
Ʊ[T��D:����U�������E�jn��Q�TZ�eEK�N��B�\�F�D&kj���mjr�f#3M��6`!��*^z	V(�/�L)�'qSS��z�s�hu��d�U�b�pD�:$�4��Þ��,2&Z�YW�'�A0�����k#fS8�Q�4M��T:#���D1Y}����ۘ��5����
˪��ӎ�#[����),ݔ�i�v��)��F�8���"���a5����	�B�̢�tX�_��{ES@��ʛ�i[j
�ꦘlE�Y���<ǔ_-��+�2p:��Ϋa"W�f��r���R�R��"3�7�A,�Á秏9��-um>�p| �D gR8�j������I�!��q:^U)��m��R��-rY��[E����Y{�#�xS���-��-ɨ��Q!edN1�&�����h�[�2���V���)�_3�_uܶ������!zӑ8�#���$��C�k�ס�I�����Џm������u�9L���ϙ��<�y ������K��[��ym΁���t/tw��TJu�=]O���<_���橿��V����w����\�-�g�ۃc?�o"ݝ����v�ѡ/��^;)˭���ȹ=N���]\��|�wup�o�z��_��/�u�;>�]�>:�w��/�����ӣK��������jݒ�=FN?�K�>x�r}���Z������_ }�$AwpO<�y���3�Wo���+7�
�z`ճ����r8(F��pq��)����,a-y}\}qv���٣'��<9��[��W�G/_��<+{�����#-����'/�?z�Ζ��������ݭ���}��O�z�]Ϩ:R�X����{��)�_���ۓ����M��1�@>��HcN�I"�f�L7���h`��HIS��j���r�,S(�hd�����_�6�I���J$�QBfg�2Ƥɪh*k��O
5�,y��#T�#(�Z�P
�+ј�8I�kF����	}��D���&�
��ZFg4 kc�**��L�!���["�D�0H���4�6gJp�4N��@�\�ߔ~Y�L"P��_J�t�U[�`m��ۧ�g�q���=����w�z�ϭ��h���?�pAZϭ�s5>;��O0����ţ��U��.n�w��?�u~�|��>������_�7�щ�L3r�}����V���Ah����9��@����4�r��J��Y`���"˩N?>��k�>�>��0e�{ۮ_m�s!���ۿ��������6������|��7��Н��X%��I1�;}׎ooϘ-�e��L�JZ9�D"�?!��ZL|!��/�
�Z���Y�I�6p�H�@j�� ���t�l([�N��ݢ�ᚧ��qZ�H��H��7-^H��O
�fĴ��ׂC�
o$�a��G���J��2�Z�6!�-�p\�q��C�/d�yQ�����O�����m*�>���p��)�л�p8��������{�w;��	Y
u�;R~�#�7�!�f��[s�PfJ��#Hi�R�Zhr�8�u�ڍ��rFȥ�)�������m���O-ߨL��FR�؈�4Vӈ�P�K�a��VkOJ:��I�۟�X�hՒ�F��cʪ(&�hZ!jR��PY��p����[z-�/�]"��TA	:B8,���㦑���'����B|�/���p�F�)gO��NN�e9���'6�:�1]���=�Nߴ��+d%�������\!�f�Q�;k�M�����ƪ��p�̗�I�1pk���QB�� �ee��FLYL��׳t[����Ӕ�,���HL��1�d��%&(j�6���2��@V��c�厈� m�HQS7"�VG'�T�$B��A�8F��@��b�Z�IA8�*FY��!�"�_H�P���N��%ҩ��4�em-,��%8qS:l!ue�)Gk�p��^
t0q8t�3��z3�F�j�#*ݘ��@09�!u����D���
��Z�L ��@>��/�(=#��h>0�-�MV��Z��M%2�8�
M��Wn���aL4dV��t��RV��L��9��
�M�ںD ��J�Ȓ�-��V	~N��O��S�X4=�V�Ndq� ��^�B@��@���/��M���� �EA��L� �TX��u����I5vbBDqXHQ�RF�(����c�d�� ��Q�_hZ�FH
�����Y��#��ZaZ-#�ĲJ�[�h�c�8DX=p�sXSQN4 B��(�����kc�B���da�Y4��<Q�}f�D;���1H��S0�L����JL�M�"�������"4m�X�U:�'-ِk�(|60����p2��^JB@R~j�@�8@r��-���)�h.�MuN&�)Ԧ�Vq��ng�i�e��3�D�z�F�qo�h��?��
�Y�(D��¬�iA������Զ���ÙZүh������X�b��Q�\�!m�t`"-ZKF��ј,�	W´�z���Q���\�1HU��S�t����$iW�LGǈԳ�k�4f���2��*'A%�ā4������l��j՞�pZr��-��6|8��hԌ-$e=�)��8Gݖ�r#��DH|�~�����s�����cT2c�!0��9�����b�aUe!F
�Z�,�@�uEزWz�4��)��4-���QnuB,~N͔�_kt$�ڱ�+�dqFm��Ul[ ��!�����/���j�,���1���A���9:9~���QK���:�n�bOi:|!)��m���J�rL��C4Po�~Q|d�FQ�F�W�0���6V�-��DQ�M��)Z�h@:L�>g��п��������.�n�^�ɺ���,-؝�^�t6�%��g:�0ݮ�u�'��X�fnO�|�����%�ILG��_^���x�μ�/�����cσ��Z_�zu}�[���[�j�����k���n|��Sz��U��*qwz�;h�}u���;�_]�Fs_�s'n�p�c����h�Ck)����[����|�����V��>��u"���������W�O}v���gO�q��/Is�r���s���ӗ�_�xh=(���ת������~|rs�s�SU�3�q�g,=�z|���PwD]|%�X��(8����.���v'����v���l�?�C�9;9��7���w��{��h}	�:C�_y�u�;�]�}���o�<>t���D�nv��a�p�z�O]��{J��o6��d�4�$M|[cjm�k�۫{���7WZj!밾��V�i�t�t*1��f�1��A8D���a]=�i9�ū5GK'�(Q
}� �����Y�F����,�E˭��H���B��'ep>���s0+���I�b߲~���X��%H��*�cL�B��tR.q!|:�'}^G��=8Ǵ\�ZmԪ\!#r6mԃi����d!%*T
$�FQ�h���3�Y�ф�uJ��P��p˷|N=H�[xMV�M����㲩E���Ë׷�_�x���ճ�'�/�<���;�x|��������ũo�>{��
�����/������G�}����~��������o��ߝ��λ����_��3�֢�~4�sQO���p���KP�'�&d��L�U����0S�|)p��P|�p��O��3�7��D'�QB��L��c��������8��'��4�9���)O���+�a ��vƱu֪� Cf�Y����HT�H���L��ei@	 ��ah+y{�qRHV��uh-|gp�q�jp[��rZJ3�T��*.���n�F�!'�A��9�(�0�� D��c�pƟiU0%�B8!�t&e_-Z"5�n4u9cnj���F·~�$�P����d?�c0���y}7)ݿ������8ǀ�>8A��0Y�B�~`U���$n!��	�Z�'}S)ej�0&�b����T4%����N�V�͡��"���1��r3YH��P4隁�*j���EVQoȵ�*���F)"W���`d�j)���$�ܜh���*���h��	���┫|r��gGJYdR4%+�aǋ��*�]��K�qtS4��WQ-!g�6*�����,L#\���:�<OJ��,�9/J֙�f�3���l�^�ns*�����������}}o0r=YH�ԧ�~�u�m)�:�*�+��*��~��OZ��ܶ�|�im�;@rg�2U8UG�)��.}x���Fɒ[��?&E.SZ�aR�6�G$�)�P�)]��S6�88��S�h�쳋��o��5;��!V���K�T]z倦u"�ޒj9@dLY8�53�1j̉1R�VZ.���_�)H���v��#�*8v ߺtb��
2ШgS��XT��8��+�f�R��Ji�I��)HLǴZڛҢ-G:��ɪ�	7�/��N����2����Cv'F:�����6F��:�|!�K�_(Z�t�Zלl�*��~�5Y'FR��G3�y{�a��rB��ukdMsT4-Tz�RPEEFM4�����A R����adV(AS)
1"F�S�U��0�H�-}�[���'đ�4&��g[BUV���ޤ�J�iʩt�ZiK�:��H�қ�ꐳ/5���<�Ѫվg�(�e��
QRQ`�1S+%_e)qF(j�pX��|�R�@ ��g�,*Z�zKG�i�V�we1 �,6~ˬ4��1�"��(ʖ��"�ۄ��K�X�e�AJ���.N� �i���4�ڃ����3M�tS|u�"�k�$3m9FV��¬���#c���/�Yz�2��L���Ò2������5
E#±��W��<h��t��F�lKx�T��3��J3�V�ۻ�9�!��8��߸/��&���F�N�e�S�$ST��r�F������%Zc���DxO�NTk\c��r�I�U�RL���#M"�/hjluM[E4�)�j�M��@�N>0N�R6�j�9��I�EYQY@p4�����[鲄��h��b&����#.��>���%�7�V�Z�Y��,�A�I:IA��Ä��l�d�s���F!�����)�f�Ѵ��q����*F0�c��k�?�*V>M�M%rz+�D3
1"��j��r$�r�ږB��Ԩ	�� '�ѩ����q��{!sԭ!��$_��"'"�i[���Vs�i�n
�$H�i�*����"K�tk�w׮�9��
q����Y{��cNj��h�B0E����?��1�㛲��ˋ���0mi���j��\���<N;l-���r>P�ƌ
����8�ժ�V��߿�j%"�B���?
!��o�oT�H�o�~��j�O������BY��=�����m7��q85��zѻ!���W7w>.8���o{R�k!�ֱ�������+u�)�v���؇�nK���yz�;x��u+�ӊ�=���+,ө{��G������Z��W�����y����ɵg�|ht��A��rS�~!��Q>�lm�?��o�Q���\��_� õ.O;���@���Ϋ��w�]��|�~�[��?����=�K�9>��n��V�yM/��W7��w�>=>;q���_�fZ�ROl�o��>zmw������>��    IDAT�;�X���� rX�ӣ��-�a��bݎ�?/��?�8;w������~�Hs�0���=�G�����GO�~�_�}��Z����8Hچ�|����gT���>���Y3kG���j��*�1M��u���@>N
�3�8�8e�C��19�E.+����@�(�n�x������.ˈä�����p�#��ԃiѦр�!�.�ωFY|�*_nc��A"�ތ��!Bz��3	�BN��"�G6�P����8r!|���	Y�PF�#�T�E�wz[)��� �(�m�-�(��5)Z{���I�߰"�J�hj!ڧ�[Rۘubu�P�A��pQ�K�����o~�_g��v�S��Ův��:�k�+���[�O�n/}E����������Ƿ/w/��ׇg��������������Ͽ������__^?{�ʁ�w��_��sfhƘ�g1�D���3ms��hO��t}h�F˴
�t~`{�')d�ɟ\Q[���KW�^I���i���K�{�F	�L���;�����_��=N7A���F��}������-!�T�v��\NM(�� t>�ןNk�+G�HS
�f~�xL�iH
rE�
�ӏ�G��&;-��O�ni~Hrtm����H)K!�Ħ�ȁhUȘg��eԌPY�B겘�@��E.D��@C�im����	�3%�B��F�)�?%��	��)p5&�٫��0�n��@���t���˭75��zP���f�=��t��MM'��[84��v\PY���a:����I�R:i5�L�;3�����U��C��T�cJ�:S��ZS"�a)m/_u8d۰�cR"p�M�t� ,wtB(�1�)G4��Wژ2��m�%`�A�d�
�CLS�B8�LӲȦ�I!��J����/1\�Y��}�t����<�	��ou)�)GHi/a��V��#3Qիb$2��9�\�����*MP�C/�O��JD?�h�K��,QS���ܡW��׫���@A�4)x�x��k�+����b�^kɫ�TK����t�r��Z�:�"/�J�j�l��)|H���$�@m�r����AX)K� �l���§cc�	m�Lc�IL����Ê��f�f����������ml$+%)`��K����ˡG�CR��H�9S���Y"�Nj��T��;?��i(��+*Ѵ�kx���FӤ�8m��Y���t:s�ԅpDW����y�qL��C�t��d�#!�����Bv�&)c�\�LT��r�0d�Q.kueMTJ
�M`Q��G.d��!6�=Y�Lh�ʴ�j�ҷ�M����R,)NdQ����$�(���χ�bRb6ZlmB� Ӛ�t4���� L�hS��X5?#�Z��i��������9��4!5�ƩOY)J�تqX�h1�2�>���Sko�lB��kUt��%TW����k	�6�mZ���o�� �m�)M-.�Ģ�'��U�V��`L-�ԕ!e4}��)pXU8i6"s�քƑ��~2I
(W����9ZŚj���PF3Ư�,f��w�����Vb�JQ���[Q�~�����TbWl�\�1\"qkIAb=W�^�@�h�RDi�Fʢ��8�评�-"�B���)~�B�JL�X��hSc�%�wSS�IOӨ�9�LuK���T�d��'n,���YY��C��o�`�i�i*�U��<"�)�g�A`-Y��8� d�Z��s&
Ih԰�jE�9F�p�)C3�W��1E��&Z����nM=�l��r��-��\�U��1��kZxk�.N%�k�!���q�kcB&Q"�I������ï��֌B�GƩ�P[����a�D�\K�7����3Du;f�$n���B"(������0qj �ڛ(0e#S����)���䈲�R�9���G���W�&���4�W8@͐:�s$D�7Ms�妜Ԍq(g�s �l}=�TqLc�4�B�8� ����d���3 G�r�Y
�#��" ���.�
E�n:)�HϗEӔ�,�c�&wx�&Z��hZ?�%;����$���v�a�,���d?�F�$�,΁;�L+�'.~��	emT�4���$5�jU�M���@����J+�a@��a�){��Nh��7��!��>@������o��f�����k�nw��aj�w��κ�צ;�nV��X��yq��9<<��f4��E� p�uOx��5�]G7���J�C}�u���v�_�Q�OL��y�[^ݚ�޾�`s��`7t��'�;{�w�;�������?��݁T�܃�=���qkQ�ԧ~�;���@K\����T����,��z����Ӌ��W���/_����ׇ�w϶����������\�����͕��~�� ����m��_��q��#��K
�|��v't[����_�}����u���]_��> L@��s3���T��:�^+��y�g|���''��?����������?_���_�ׯΎ�Xғ�GO=�����ͯ����ן~J{}/���Yh��u�'V�������`u�QE��n!#dk~�� d8�����B�q�<Rx�(g�g�^&@Y��):���g�bҡ`�*7 &�&�_9�a4`���i&��������L�dK7-��\'�q���T(��B҄0���TZ4BS��qd%gu���\!;��a"�Y��z���F�5�p�n�M��9��JA�=�T"�*��HL����F8�h��z#+���t׳)�~t�v;c��4�@c�V.�P�+�3ٔ��Z�:�ޗ������{.�t<������z8��nw�n����'��^��^�_�����_���nmz�<l����/�/�xv}w���K������MKz�r��W�^�x��_��_y��;f������?���>�v��&�m�D?p�MJ�[B�bg�Ţ�g�h�8�e�h�"�}���HV�Ͻ������h�|��z��W.)��rV���}��D�'?���+�6��S��'�x4��K�v9�9�JhJΚ9Rt��{�@�@�}:�lS���b�S�0���iwL9�Zy)F��MY�D�FK��E�������W�"*]�iu[,����稒�ĚA?0��dq,�~Q#B��O'E#�9F�rk/$��1�?�������C־�WKϟ�8S��Ѽ܏q�Meg�{��{L�;�g�}f�z�8)�iNP'���x/'Vӊ��B�f�s���#�X$�V��%��2�N�q�VQ4����Sj�;���i��#Ҟ�K1%ŗ����/Z�*������}!�!:"�3�G�S����QEK�v	��fʅ��W�iUG�nJ}�n� ��F���,MF_?Ƣ9r�Q)�i*Z�kk�.+<5�Pˁ0�t�r[~��&Z{����*�-�XWh�Z����G�2�A�,N���Q��ׅ��cR��e�8F�8t�zQ�.���w%����Z9g/����l��;�?�����ҹ�cj�<�^5
)��j۔k�9F@" CH�YYpQ)U,�m��J�\`�BD��/}Bu%Ǣ��H]UQ(S�ß=7Ec��*v�c�.Q@`u�9����Ւ���*�._V��q�(�STn��GJ�kX'��ⴓ��6y���F!F��1�#��s"��D�7"�ߙ��L��"E?���t~]��6�X���޼��F+Zu�Y��2��#�ͪ���%�隚\�!�S�nј�Dp)��GM!~��z�)9�Z�?S�������N��2N|���6X���)ь�����4e8���m�LtB�lW%�����pd�J4"@"��2��>��-�������ϟPVtZU����?�I*��A9�fV��Z� :"r1�[�љ�éе"��?��+�z6������s*
��r��V�8��9�SL��ODu1Vh�*j��(���N�_����,d��G��%mp"v�"Z!�V�8B�Ţ�k�t�����*%rj�'\�D��rG�Q3Bj̘N�+*���ș��%6V_�Zo+���e�t
83&U���5#TK��R �*Z��tx]�Ge|� ��"���lZ���Z��Ё��q��()8B"���t8�9F�D��0+>��H-���7��M-x���[:N�Z��B�w@�ki8��D@�'�g�a)!�8�h,�ω �N�O�hSkMFS��t,Әr�X�����i��������Ff�	 ��8r>��f�*
�@
�t*���s�"�ڪ��c�^)m��ȗ(��1�+!�Tv�,��RDɊr��M9�pX:��"�Q�W��&�ol�HPEQ�q8��J!#�VY�K�T�Ψ�l�	vhR3ʅ�C�!�
A҇Tה�hM�t�ҩ(�*����U�M�@L8&
a%v�7�܂k05��/1�Ғ�9�%.�7����6g�bΘx���(�p
���9i65F�����dmL�*�������k8���~�kEFj^GUO܈�j5�A(Ki!���8mґ�Q��f8>��_���&A�MS��ϵZ.�\x�uR�ri���k�5'��
%R
���>����>$s�f�����Զ��Ȧ���~s�_�\��Q�}�q�n�:9�^�6dk��ڷ����c�5=4y��W�������z��|������b�G<�ŷ�����)��=:���/�}����wǮ�Y��⭛��?��6���ѧ��Z�=��E�[���j����1�89s_pi��]�O0�]�n,g�qqPov������G���/�^��zv��vsx�o��\^�]�ܟ����/�t��Y|}��Z���@O��zgs�	Q���%�ֻ��C;s�j�*X}�R��|R�L�[ h�{����U���N_���|�����W�KΩ�szxw~qz���[/_�r��_���ZO	__]�GN������W�������s��b�T��|Th��ƶ꫻����_s�k����
����(4"��::o.kC E6�/�8������GK����O�!�#7f"rHm�%�EK��`8dD3�DS|#2|�M��㴙q�9UoZ�*� �j7Z�1�>�
5��28�L��F���f��|��Wc���߷�S]]�Ѥ`�j�w*&�J��&���I��"ȝ�%J���  #Cp�SV%���kR�}��
l��O	���EV�uP�5�n�0��=z�����g����������sJ�Chv��E������*Bswu�ꫛ�����w�w�o}���]�p=�z����_]]������B>+�U>jv��?����3���8R�;�.>)d��hpS�DQ״BKq;ILӬ�ޭ�9#�M��?�y�>!��O��)C��� ]Z�	���ޕ}���Q0���qU���޹�¦VeGՖa�o�$��pY�PcNj%"�1��I�1���s��jM���ç��ɩ��a2˴(k��?�375��R�6yw��ʩR?r�q�s��jE��r���� 8K�iJ�n�I��0�
��/���,��rM�$FH�/Z�M��M���lbk ��uzر��{0�)�+�F�����B8� �٩I��|Ϣ���O?�T�L;���`��������Մ���5�?_VHEL)�t�A:DJ� dz3�>Mdcb$"�TT:5���
[�B�V��\��Z��p4�����G4r:j�Y�NN���W�\`����`ɩz���K��y82!L"F����B�6"�m+j��(�%��8q�g�<�3��q�:O(8�����ҡt�p҄��drMᎂ+5�8R�,��=7|�%Jl� �qAp���tF��#���hs��sx��mH'�8��TT�gN]����J-�Є��*]?�w��!]���U�J5@G{��pU(��D�Z^/|V'4�����'Q-Ⲉ��s �'b�hg��J�� )�����EfB���(\T{t�w-�O�6Lm�l'�aʢv������%&(��E˭.��#3[Y�"�\��8d�!��h|��>k~^be�DV%��8dM2~�L���4��ɩ�h�[��U���h�.e
�GzN%(�ԕt�"f��	�t����]�I��*�>���ي<,�rE[��4��!sHpZT.0~ˡ@��aEK����s>��O֝5YvW��9#$��	�`i*M�2�Q���fz����KY?���T2�E�"D�$�sd�����9h���/_�{�sODܓ�^SL8�`�4G�#
A��ϗ5�CH�b�odڥaƩ��	��ϯ(A�%��� M|�&��tYN�Aj��ԕXK��f��)��1+!�/ګ�/�23��@+%��Fs�c�id	rX�F��Ч&��/*�	oZ]��-0}�8��S8~#G�zU�Mc�Tm� �7�����d%�]�
9:d�h#��H͛���F�e1�9d��P	�r8�|?��r�	q �'��T���:��W�XV���c������B~R��|=;���d�Z5�c8�%�Oc�J7br�3�g�^h�S4�R��^'�&h"Z���SSzY8� ��� w�
I�ϪRi���	4�QhM+].��Y!���[#�D#��i"�����6��R���F`g|j�FS4S|f�'kd���{e��,$䱢0���VQ �V��Nu����B("�S�77e��(�U�M��]E��R�U4�WW:3%�M�4�bd+�ɯ�,8��q�Y�B��4�D9�C�1�e����LɊ���1p˻�9|�8����_b4 �2���iU������F��/:�7R@�*��٥��z7f��^����`B��H		4�^K�:Y��B��d�@�Z�T�L'�@�&j��"p,9��i����J@*m��2��q��+��)7�Ѯ�?�Nk�@'Ov�����@�4�I�Suc��!#�>�*��l@�a
3>e���K)Zn˄ ��45&>U&wN��嶓F)I���a�I!NLR���9L�2�2��/*�M���`��,���,C`p-�0�&��a�+a���;}!5CPJ6`nzSh�߽�h*�?��~�Lԋ�%H�]�J�)�e�[N������W	��A���vT׆�-(���.	߉�덒��`��
ў��>{և��9�)�uQ�L�z*��q�нI�m\OOZ��s-�*�DZY�3b���R�!p�P����J�ڻ��������U��үg��nIX����[��II��vw��ק�.D���UHp�`;���tW���^�T���;tK�ڝW��{x�z�D=}����ɋ'_^������͍O�zzv��L�x������c��v�����z`so=����o߶�cm��9M?&��������m�����w(;���N�����_yWǴ��|�_�������������=~��;GǗ/���_���|�����:s}�����NO�<y�Y�j���9C�8^<}��ً���>�s�{S��ͨ�u��^h��4�.�o��f|��̔`8?���)ˎA���}b����!#4�tR�P�,'��4ME+�g��`�4%�m�D�h��a5 I_"�V7��;�Bdq��DC���������6��Ak-���:!`F�7e�RKR�N�g�:��ȇ��䆸�!���PS4N�PEk��sե��Ω'��r�Ĝ��$:xѦRvG���.�HM?���~8R��_�z�}��j�Fy������]n�n��Ϟ�Z������˽����;qt��O<��w���Tg���$��w6]'?������������S�P|prx���W��.�[�n����A��9s��?���L�+S�ykN�3���6�>P�b��1Mg���c��~?���o���|���s��{Va-�������>1��+~�V%�뚾�W��i��!WX#��m_8B��2֊J�`,�)�KU�NQ#A ���M9�i��x�8R裙�E!v�3e��Bt�2Bb_��뮀�IM.�L�,&��
�2n��E���7-:Ǹh,�9S~%JG(��Tի5L�ȵTnQ!��W���&e��mT��9�ǡ�k�
���2ng~���yu
��c'�n��q(�2�K�}u�D�������I�2g �^Zz�]9u�N�L�������>q[���=A��dnQ�����%�NKRN0�H    IDAT�ґ�핒Id�:�0q��W�!�eqb6U��e��.���2�N�~4�)%�X��|:!�$�G�cR6���2�pVim�94���/�[�&D6eӪh�m���l{� 5���U�)d��U~3RN�~Ȳ�`�*QEG�,�'�qp�+D��
�8��t���H���J����ݯm!��� �I�N�����^�������h�'��+�(P�]j�?�l������r�R�4:-U�@����g(:qA���EV-S=+��
��XW�bBl&<��d8p�~� 9!�D�L㏓�����
D��!\���ٖw[���О���؍F[g���%��,��F�4��ۖd1�G���Vs�?Uh�ˑ��4�� �G���4mu��
����HA'��TM"�ndUOJ(S+��;��8�|~��ΖԬ�D���3�r�g>Ac�R�`|W����)\.P�n�h�d����ʲv~��)�~��"ೢF�
|̤8�J�S
�S��534Ѥ�k{�g0��N�ơ6m��0K���c���_�3�����3F�($B��]r�j��,��&��%��]�VA9�~�D<Y�pSfjM���ʊ9QS`�Btbv�(�+�ƨ��eD	�d�3=�%%�YjM!C��[�9F/QHm�;MƑX:��>|�X��9 ����p�v�m�[89�[�$��B)�S�P�dfjLg����֦�bR�ԭ��C��d��o�db�V��!p�M9&Nxd�)Bj�5S�@ʳ9�*�§����Y��FՅ8⨕hJ���9��i�h�55Je[��W�;�f-��p*����i���1���R�H�*�-�Ⱦ&NG�V-�h5÷	Br��#�Rx��z �!���o�)��x�������j����9�_�R]xR
!$^oBq�	�� f|Sx &�X�g��R4ZY�	r�hdY�
������X'�͜B8Y����V�ԆC��z��A��JY8>_�:��e	1|�zd:��J�N	!�i�O�~�Ĳjc*N�-J�*���C�f!��L!g�o�X��i���H�%�<�����m�����3�o�mN�Q�/�[�t��hL�㮳��oE�I�ϔC���M����'��tw4�%�r���ڥ��I�=��Sn��鳖�y!%����m!HY���G�Z��s Ma�M�l:~Ȍ9�bȥ�BY:FQ֋4�uu��@
���V�P��0D���c�1�	L���c��Q������3D�1!r��KY��|�眇����Z�Y���Y�P:��׺i>��vLi%�H;�Z���I�%�À��R�Ӓ��x�����m���8\�}2�ʢ��9�uK�� ѬmGÝA��x��%��>o��}�G']�W�7W�A�@k=��r�6��E��Ӂ��t�n�G�z,����]z`����8�	n9��[ypa������={���x��ѽ����Co����%�X<���!�뮧�QJ�G�Z����e��Nk�7��o�8�+��z��5O~�[���1'Ѓ�{��/c������{�y�Τ�8<��ֻ�{x��ޫ�����c�>J���O�=ֻ[��AI?�G��__\�f����O��9Fn?l����x�S}��������v�����/!vX����zw����l�'����/���w����~u�������ruyv�������oX۴�Sp�d|����ػQ���o�������V�w���|+�S��ض��1�a#�h-�+a3� q,A�|)�@X��N������1��sr��qL�N����	:|�66��Ѐр)l��lY+B�J��S��eD��0��@���@sd'�D!��BF�^��BX�ݔz�d��F�Z-�qc-%?�Ґ��(��pNu[��f�w�t��W���	gr�ғ�]QH���wD��S�)�\?�k�Z���eQ(+G"�~�X/�-1���]�C�/
᫨.��\�)#�Б��/&!4o�AHy�ح;S���}e�٫˷�aO�K���s�{~~�c�|��_����>�֭M��l�=e��{G������ή�����'�_�<��郣g��鑙�
Y��{��m����:\ϭ�T{�o���2�c'1��痲�����c�@�jǒ*S�p7���1g�ڥO�C���?��-t���=����+$��Ubmn��PM+֛��,5\1�b:�g|H�|��~>�����@� 
�~k�@$r����J����`M�f��4$�h�Owt����`o��8�F�N��B�F6xS�ğ�Gh,�L���(�9��	os�Ji*4�� �#���r�1j��«��*�U��W��n�`�CS�۫�M�Bv��0����O��O֡3������tP�o�&�b{ұ��_{]	��9@�L�y��nPg�>�%�%�!Ȓ���>`Jt�z�p���1��McE���2�-V��:DJ
pk-r9�ш3!|N�1�A*�P
5��	d�!9�1Z������U}~)S���`��\�J6_Zm���c�y��z�A�@�,٘��� ��3�	�w�tVp4P?8t�kC�Í�CL�hE9�
�5�U���}y�׈��^((ыH�ZB�֘&A�l�1+��i	A�i�H�NHW|�4��p4�y�h�Ԉlg8��������Rd�J�K�)�tF&���pb�2S��r��
M�,��p�
��[�h������3��U�vd�N�c:M�	��nS`|�FS"B���#E%&�c��h�L�TH]���(Aǝ�
! oy�[-]���Ԃ�b�v� �K���"ht��Y�~�{9�1XW�p���TVu%��#+�|�#�?����yk��h�H{�S��H'p�Y��h��Y9S_N6挬�\��(�| A�t����5�Ʒ��hq��6���⌟���>�)}*˸
l���a闈�7>}�t���1;1ve��h���|�� �e49x|�
�>����)��Yb!S���\"�"6"�݊᭥*-�BR����Y��J�)�����0���/=����v��L3>}
�;k�֘H��*�-����1K�/�+k��Ml'y����L3L�)6�ၢ]�9�h�9F`�C���j�n�䦃&ר7Y��EM��8+�5Isw��]r�Յ�h��F)9��i~-i �L�����r�g~RES��;:�b�m�h*Ć���?��l�t"�_n��h��@$2GS3M�2��qF�cӀ���mc��U;��L5P�1v���(��h[������K*A�(��Z�&�`
7�%΀��8!F`R��BH�����)g��:��n�ӈ͈9�1��ٮ��ئ�&g�Em��I�2��*ZK2��?��	q��1ՏQ-��7�\#�,!�o�C
5PQ��B��<��j5��(�jIM3�4��Hu(M�YY-���V"?YHS`-�C������/2-�N=M�ҧ�Z8LT��2����%@�����Ҷ�D�巓�R��������d	�V�_-�U�I�\�8�B~�U=r $���U�pX�"��-D�q���J˂�ْV�p�i
���C�ί��QFk�p֞@h
ɍ�g��h���aS�,g�0�����p"1����B��;���7K���?R|�dq�\&ן<������X�Zާ��_9z]�0:m��-jZ����A��Rd-�g�@r��o�0!��ƖS�B�z���s�E��[=��6��W�u"lOUn/:��i�F���R��#[+�Μn�|��G)�A��Z��zp|yqy�q��L��zI���6�'���=��s^} �/�t7�}Fo����\�{����-k}���i���(BsO���S]��;� ־��{�N��l�o=���ua_�5�G"7�Z���@�d�NDܦ<:�?��њ�㇧����O}��������d�YO5yg�]������{	������9Y�_��{�����ʯ�v��\oN]x<4u�vs��r��b�r�����kϕn�뀠{|j�W���6�ۢ�Z	�<�f����#�]�:�|e��z�?����'�|�����O>zxp�����w~���O/_=�����������=9������ŗ�����3_��ɧO�=���/�����������/�Q����:%��Кs���y;��Zҡq�	��qƗ>H�2����1+'Ds�m̶c}W�)��][�m�
'2�����a1�ESs�U�����q��?Q|�5c�lZV���ΆUN��M>��1JمnL�#?�PK��C
�!_���cW�\{�Ǉ��s�@��Y{Cn�ZB�*�k�1J�6�����ۙ8Ս���ZU�3�J���ƇcүO��B��:�c�M��~. ���m=?��1�V���>��coО��r�{��w�y��o?x����������/�Ξm����g\#���\�Nߣ�Ѝ�˛�S-}��;�������Y���W�|�o��|-���������h�W!m]����.�lɁ|`8Z�oOvG!S�6�c�q�gz�;|��}l��F�Zh.V:'�'��v�������1�B uK���*��g�ٍ(L�P�4JdZ�3M�H����ф��Aۀ58	"�q�EU7�oĄLA	~̐D�1S3�(�P%i+e����>#��\]���|"iV�}4��v�� P���J_Xz��Jd�F����(��,�>��B���#���Z8M�:�}�ۤӣB�+w����� 8ݼ�V�%3ۛH������?��Sӆ���u�z\3���qV8]���է���)�q>�2!�M�@>M�4�qǈr�	d�Kl�F�R$2��&�L�R�y�힮��-]R�MɊ�6YrQNQ BK�蓂hj�`��$�����#�Bf����,�_�(��$��(,JP����S0ŧn$"�QhQ8�4�r�B���9BL"��Z�]���d��E��ȡ��h�"QoM�Wr%Y�w%�t�q(��u"�������������=�����^,}�qw�����aM��-����^h^YB��'�eb\�5�ԵL�Bz�n�CF�
�+�1f����"�a!c�|��8mu�!m�/K
�PQS6�Bs���L��1�W���)�(G�EY,��
v��@d������g|8����	A���m���XB���`��`�����[�� �XJN�8JD�3
�i:�Q5 �0Eu�> �h��(,���;�w_��-�&sR9��{nwyO�Uڅ���mo������3�"��9����`Z��%�;����#�W.G��kH\{1'Z�sP |H��5����P��_W8��RS�'Q�[B�Ƒ�5x>�X��B���X{F���Bjc�x�Ms�G!�Z����!�¤��5"o�3}-\��;��|"��>R��GH��P+2>'�4M�Q��Eh�C�6*�/_�pH`=�M�.~����� ��nV]-��#
�5�_	H�,N�M�ሲz�R�'����fQe�U8�j�2S&�f�n*�����s�D�)૳;Gȸ
߭��O_��$X��7���*�O%�r�m�DQ����,�t�������3q�6��K1%h�`��1��2S�(N}��@
��V���T8�F��Ek�X3u8E���'�i��h���>�G��дƤ�HgU�O�ᐦ�z��d��M�A#d��:	L�N�@��Gg�Ĕ�h,7�fYz���3���(�����%j��Zl)*�O?AT����ݫx��r�E&.j�_	�@�
��YݢJ�
��@�
��9�Bڜ����)}�,�BF�t!ǗH���U?��Ѫh�o�0#��X:��|������-��h�f �|��A��Ķ(Z)��Ҷ��)׸+n��r�[?F�B��DP"���Tb-M�Ѫ.Ti����|�Z]mZ����J�ml7G�8��8D�>5���0�1�Zm�^��7���a)Q�@�6���'�t־�ӱ����K�U���5�bDK����@�����Jt�OA�aG��i���	n+%��nWKhEK��+�Pc5��H��RH����E�Fh�Кv�M���-�A���Cf����α��1�?���qX��M��2m�C�,���	�F:j��4ӏ��E�Xc�tL%����$�/�B;��G|�|�fBn+j_�m��b��+wps�$���ӵ�{'W�r��ދ����#}���|_*���o��_����"M���>��҅���CE�����;��z���䱗��O�=q��7i�]��z�z&yzt|��������_��\x�^��xsy��O��-�ۉ-W�����͜�=w}������������ë��W�u���cu}a�ͱ�����g���ٺm�;�뎯���'ۓ�7�����7�y~�톋W�g���G�^�����H���u�s�sv�u���`?EW��dZ�}=C�~������%B���}s�5Ĵ�4���7�1�����)��G�uz��t�4`'�/y}|�C'��c��;�����O�`K���z�����dm�����<�w�ҪdrW��p{9Z{����V�_nSN�����n4)c�4{q��b�>�N`c��TȔI4Bf�T�8���� )�y GJ�|"�Wn��/$�+�&+����8�ܜ��b�ij]: ��8C棵@�pc�A�U��oʄ�r|�[`�q��d�n��6Z���4�8������&ŇT�8B�"R��Ƒ*���fD5����(��Ȗ8uӔY�����4b�9'2�k���W��_ޭvѺw�1���|u�c�]�����LW��a����/�/����,\_�>y��7C~�՗O^������+�_�ZO��ۿ��s������w���]o�i�{}��n�'x�ϛ�9kE�Dh39�w�i���f�	v��!�	�:1�v�(�����*����xC��4�[�땆]��gC�*w�����kOr7�*�	�
h��!�B~��m�\��	�)�4��|jD�h�c�El�&��f�-U�E)�F0�E�-��g�|d�1��z(�\☌�mE�k���B��5R2�:��V�l�8��i+�r�@~�i�����:rLN���Gٴ�k�k
F3�3!j���:È8����^:��l�� �k�q�H��IG�S�"��G��Z���J���C K���mt��B�#��~Z��|����@gWg���V��+�\RS3J,�	o?�H�b�CYh5f�,V��JG����k���@� �r4��G0B�iAE#0?��:ASc�7�Q4$�#[:�&9��X�N0�:�o�����v�(�r��gg�M�>�c�7��>q�G����>?����ɅS#R!
���NEW9>�!�R��j��qz�QA��E�Uc��5�f�}�����>�UX�N<�S�k��e���>wO���Y�^��e�.���pu�7��x�5�
r;ßMS�4�F ��[/�%�2��F~��~�߮W*�m���
EK�Tn����~��P���~~�ad�j�/��/�����udY�&�.����.j���--�SK|%Z~k��V�@c�h�3��(�J��:�ĉ�x:�η�Bh�/�4!�F�i�W����A��"r�J+!E:�R��v�2}!��ҍ�4������'S��QbMr��fd�9��E��'���|w��CK\4
1V"����B-��`֏h��s���4?��9F�ƌ)�e��M�4gu��^�Ȁ����":��7*��lZ(��*��&=>$��w	��-G	c'������|
9��lS#)��9����J s�sp r�m��ݫ��A3�]�~ ���ߴB#Ȫ�B�V��#kƴ*�hU�]}M!N%����+x"��W�r�UlZ����C0� $eAh�9�q�Ф��93��#s��s�R�wr�A�_B�|�Xx����h�D��p�H�T(q��I��e��V9S����:m�Q�9q�B���v��c��ѬcV��p�T��K�h�P��e����tcN )-I���?=�Y�ӪL��o���BY��U4Jq\�#�J��E�C�Q��E1E�pX�#��5d��b�\*��s�DL�1m�P���    IDAT�>k,�9�,\:�O!%��PSmDC�d����YR��mv/�U~k�,���]�G�3�|�T1E�h�B�˅sK�P��]��T�hm�Q�U
�cC:LC��4NuNY���)k�)�gXI�@���-n:L>[��&�TĴr�NZ`:����l]�F4 ��m:FS�DD�N�I�$R��vY-���S�W(ZYh,q��ĎE�(���%�tR��D��o�n+)q��,den=�,1��e�,�D-A�ɶv")�B���x
�%�Y%����˂�d�\8B��B*�a�S���B�4�D8�!BF�cmsj�?�i�r)4��v��h��ZM�H������i'Z�����"��4� @V��	P�	E�:K]|��?~����v�3�LiS�Q!
h�������'�ŗ(Ř�&-
�XtB��1�X�x�	�M�)Kk����l��j�G����[�����S`�XS����f�ݬC�����طO�����Z�t��ʭ7G���K�Wmn?X��4�/C����ۉ��^u�>�֕���-�=9�&����������__�i=�h�������s7!�,rCԗ�~�\ݒt&�|]�ONݾ�r}֬�;����pG�m�Uq�IW+wX�vx�si׍=�z�S��C+����B̋��������￼�Ք���Qp��������W�y��'˺=�k5�_z�-M�������<�{vuy�汛�V}�A�F>�>9�麇n����7�ί�,�V��q4Z����8���1:���o��75�����{n��x�j����w��������'�{������B� q���˳ާ���8���%��ʇԭ=�s�j��؁��V�������Ac��!�Ndc��r��OD"��1S.˹-��4J1�	����|њ��m���eG�����g�qd��mg��E��Y�)���[.!zse)g���gZ2B2~�C�[�%`�8���uRS�S�إo��ߘȴ�����Om���W�6Y(�K�Sf)3�dۍ|4S�����Q�i�,wdEmz���I8 g���bL�i�� �c1GB�\j��un�!�B�F?2n�{߸(Ķ��$��{g�X�*�+3]��\��O���<|yy������9���7�%��+W
K�9��Q��������?������o���������g�}���o���{t���Ǐ������o}����mm�(��yS�{U{�q�0�Y]{eQ�U�W5g|�옵���rDu�����V)v��Ў���ު՞�B5&Ż��ԅ�X�v�]LY�K���B���˿��uK�[M��v�Og/0o�3+��ʐC��[�n�t)@|�"H�&�1*ϑN��X[c�cL�SKñH�~j	M!u)T�d8��1U����D͸`�u��z�C�@�J�?Q�,s�*��i"L{Ȧc�z#[c
�Y
��(� 2��,~���G��� ���GܔaԵc��lqD|��[^'�?OJ���ч~���d3����z������B�w�竐ו��~ui��C0M�hd������G����&j���dZ,�Ӳ�g��B)8���eg��JG�7��)��K1����%K���ў�t�מ���b���p�E��M�o��%X q`E9�c$eJ��U�FC��D��6
�k��YIM�t|˜B8�O�h��!x���dnU�k��hR��Zk�)��Vۍ[��8�s�h -Y�$�Mш�m_]��
��S��׭D��:�e��'�7�}Mj�!�W�Ӫg��p>Y|/7/�"$z)Q�FRD�Ĝ�'�H�0]�]��2j� �~�Y�l��τ��C4��סi9��+!��'���F)����o�χw��ԧ��/eS]��n����,�s����M!WWu{e�l��奣q�1�
��|c������	�#3E�����hF�-Hd���ˉp$V��/s����SH�#�(=p)n�zg�(�$�	�H:FQ����裏\�#���Cpֹ��@;��Ӑ��V3B��2��:�c�c�0!��KG���|>3exk��L����9���B$� �49�0��f��u��l��t(�G"\E�p��"*�^�H�5��"ue��J��X
0�t��u��Y��7�J��o1MC��5%(2�Ĕ^W�M�$�S3����2�A���O��F�NLьb�V�N�Q�OKZ��M���i)�.��օäO��(��V��n�#7��H��k^Դ���t���p�6���D�D�ϩ=��N"��!C�	2���36�ҷ�z�B]�i�AЄLNR)���J7�2ZI͈7�p|~)S��-w�
�9�6��N-x��Em�EE����Ez��n�z�DPtV������"����8;	�׌�ݍ
�P�!�P�ӟ����-�\L&�4��B����C�8tXS�ix�BvC��Fx)+s;!q8BFU:����&�NR@N0\��r��F�Cp2>}�!b���R�C�� :@ſ ,>Gn�td���!�0���z[>�����Eܔ�n��� �*A�Á3~]m�zɣ�G�#�̏�g���(D��2Ei&B����p�R��7�'Nu[�)���/Z��'n:'-�B"e��W_�G4�:ԕCi��RR��{BB���_�p���Q�/��N�|UDqRqN&Z��������I�r�h��v����tH�4��&d�o!���gw���� �.>ĴQ:�1�� �9
���Js�0�iL���@!~���*P��d��B�8�0Ia����|�+�Y��T�2"�p�A��ow�HS�"FLY,G�*��&v��g��DH-d��	&��q4�Ӻ �� ~-�3�b�*}����9rwK�����E�\���������h��#s�(��Q��3�\.r+2��Bj��8r�1Z�����|Q��ugs��[�H/}��$=��=���'���?4���Q/����#7�|����r�����_������my���]})&ڡ{z�7n���y��ϕ�N6����N ���h��R�Ļ���Q���ux쬥y���o3]n_�6�_V�k�y�r;����۹�jr��_��X�g_=��֣Û���#ߚ�N�z������ޓ߾8>�:{�ȫ�W|]�ӳ�n�Z��0�s7�N±竮�Owvy��z}��뽫�מW]�ܺ�ps�c����]�� u����/v`m�v��
�7'�7��~]Gу���_z�����/��p����=���{Io�C����xk}��/^|�N�Ճ�S/��_?��7�/�ó>�멷jѴ�V�����i-9�|�`E1�(?��q��h,Y[�β�
N�B���MT.?0�4͐��EM{5	�$e,E:)�Ԫ"W���%�h��-��'�� �RPވ��986�T�6� �KAoE@!�,#pi�G �Qu!N�&1e|8$�|�ڈi+j�^!|!KG��q��m?�5#hD��O��Y���Ch��*S���I~mFK��nᜑE~!QV	�(}�}Ʒ�^tޒ�|>�{����;o'��S����������ɣ�gG7�|�Wj��}q��}�|���r}p�|q�������ދ�O���o�����W%7_��M_����F����-eWџ9���oA��I?X[�)Ǟ8����:�@?�L��l��@�BhL
��(4Y3QK?���|-�ub�٤o�{��'?����p����?���|��yR%Iԍ����e��R��]I8����%x;u��P��qZ��"T�TH-R�S"��<d�z �<��^���Zn[�0f*|��G��%���խyⲨi��1Ǉ�b��BFH~=��j�F|���?%�JLSY�(#������o����/� $G�ҍ%��-�
!0�ݣ�����?��O�<옃��o~��:��D9G�>"�駟v;���=�z��]^��s�OǛ銶�8��C#���4ocq�;�HW�r�h�s�#�I)��**adU4�>��7E�
#<�~�U�iRH��Hn��7me!M.M`mLc�[��Ñ���W�#�AV��Hg16�g��t8��X!���S�B�V����M]S&KQ���FH��ç����x�?�!s?Fz��[�[!5�ٔ!X��G���m�&t���Rk�1`�1���rj�ژ�"�PC����~�3�C������j��V�~��:�{x����[tJ;�)HW��_�Ә,MkԳ�|/����R��V�:�ƌBȺm��M9N��2eR��7��O e
4K��/�_�(fk���U�F�pf*�X�B���ΚF6�'��:�o}�}Mw�l �W��lH��F):Ƙ9��,�~贽�����B�8��y'U��bNi�Uc�%���hF�@>�M���cu�*�zX9ے�?r�j[cq�Щh�DqZ�\!S���M)�:��ҵ�A+TE �(��p�,�X�3d���"@���׆�����5!�r�ҍ���h�R3Vd��F��)�/��*�ѕ�i��Ɩ G6�cl	��IA'Bhe�n���KAC��JJ4ń�W1���
����1+J�	6RBR~�T˨Cf#��NY�0���tb�Zu/F�V�߷NeI� ��P	E劚�#3 ��i��l���k�1��;�-J���Vo�
]�dA$f8���v�ç�p�Y��|4x#05!)�q���4`� �B]�eRXuӬa~:�
>��X���BS�4Z:�!��j�+��RʕE��(h�+�\�F�*F)�E�E��m��g��`u8���I<�g!�z3
Տr���0E��I!S�e8�Á����h��B�~rM-�)���m���+�6GH�#�=Y�����F�F&R��k:�)ZȀ�(G*B��eդr�~dcm�>�9�V��iZ�ìHԴ���p�CD��r�R�ۜUl�"B��cl*�S?8��K�N�i�h�!M�����B����&4:S��*��L.'�P��l4�M�UT�Z%���J7�"ǡ���:	�`�+�T
@ӐjA"�7&�� ڔ��B�DK7�4�kJ
�)愙(�uq�Ԃ�N��ąZrQ���
��y��`͗bL$~�DR0-Z�F��4�i�>Ĉi���T8�V�G��2`8$P'��F�}aF����e���3D�*T	H|�R��R�Ww�"�)����-o�,�_��v�i_��6�0sR����sW8d��W7���� eSVc~��%&4
!S�QF�!N`c�,�U`
2���B�t���}���|<�^?-U�͏���~L���[�)g��5ή~j����a�p�� 0m�G�\4}b�Ҝ�t�l�!�m��eN6�_�T����`�9�~�������W붦>�O�<��/F�j��4R�7숨触��+t閡���q������b���핥%?�/������ ������ҹtKn��ZR�')=��;)o��+�%�>(u���8twt�΂�{(�{�Q��=jxx,�!�Z��Z�� Y���tkv���M�7��,o?xHp���n�_��y��>������|yqpqpr�����#_zv~qsx����˗��<{����w侨��\�c_�|�K==�������µQ�����W���Mwɻ��v�η[����� ���s\��f����H�}���z��؋�W��姯���ɗ_�?}�S����s��Ӫ�C���7N�?|��O�.��l�w��\�>5�ſ��O����7�<����zqo@)�1�X�J7�k��acxBb�iNS�-0���9���vXb�iY8YՍ��uCz�%^ۦȁ�$+��	Y���R��m+%�I�t|
|g�PW�Q�S0������nÛr��J���c�.Qu�t\	o{�N�*6�sbw�IOM���[�h�3FF���f��]�p)9�v+��F���pU"���LfSN��H�ū�S�q �?S4f
�&���P>ZN�М�Q�!�C0u���t�p ����Ե��jO����ӗO~sxtϿ�8�Y�v������������_��ܿ���}��[o��//�\<;���O��_���_��x�������g���/~�󟻻������Ξ7�TR�&���Z�0'P{pm���i�DZ f`���������w���# 	�W<��㍌�C�,!�{;���yS�O�����>��#���P��NBf}3���
kE�2j uK�a�D˪E����H���]�u
i�Ȍ���,�T�.%�b$���M�7jI�vX�w�1�p(1S7�B�fd��42~S��|8edj�p��1~��0)�i+�|�R�I� L.N4#�1�5�	��4&B�)Z�@
�!���X��!��I��3S
�񼔻�׌�7���[5G����G}�q,����#�(�k��c�0ռ�&AZc[dZ�U�w��H���� �YpNk�qj�Y���82���l��N˯4�:��I��w�D��1����hjD����2�lF0�����T��X��Ɋ2j���� ��Ȫ�(��MƇ3<_	|�l�Z
�tZW)�!��*��b!�\ጠr�jY���m�����=����i4e{5"C�`���.��;�s�:���e�5׫������ٟ�ٟ�ɟ���?�؋���u�=߲�����OʿAq5�Ѳ^h���|'��7>���Qkzp#���+m�|K
�C��i���%Zo����[b)FSQ�6��	��0�,#ƏVT.��3���D��蘆?�i[���.���N��NR����%BJ[���صT�u�US�D&�k�7�D�84!MU21��Bt0>�Q��UI���NQ#��Tj�8����Hav��]S�h*u趥tg��%�r�ܙV��a�m�O�_c�j5�RzS4S����و�+U�r�ɤ"�q�#��7�bmNucN	L��(�bJ�o���h�#]�t������S�eApNH#Nէ+xg�;(��R�����*��7J$�W��yX!�u"����;1�g"��npLUguG�$2����ª� L��ŖX���Q��pS8��#w���^bV15�"W���d�,m�Bp�
�W�% ��L����ρ0Ӛ̯zuklr��2M$fG�B!tL�ŷ�Ui{S�gdVȔ����(���4���E�ml	��iV�P)Se��SgZj��XN颉ӬCSfʪ���r�P0�!��w��E9F�D~#��є勲����I�a��@�V]Y��a"�1�vC�-��4�cJG6�8@�v)��#D3Jd�R*m��(�Iߴ�L:�t�>�����no��)�N�Mᅌ��j,$��-��=ъBXd�Ħ��M{]Z�c��󢦢�S6!R�I�O��]4�ÈLR�뭳9������n�t���(T-)���)�X��"Y8m,��[�)S6��$0>�F0�T�ǡ��8u�#9GEV�4>�E��L�d����3#�:�nMB�C���I"�*�Nu � D���XԔf�qL�K��R ��r�L#�k0D��K�i�������j�,��;LY��%�ol���)�������7����-�!�g
pS��5iQ�� �L�1�7M"�,�u���L�ȏ#�ܑ�WG�9T�(����*&,��^Y�L��0�Q�C6��S'�c�[�d��5
U��ZQcL C�7�Ʃ�L�V�(e#B��L
G�_�}�ѿ�˿@�c�Dh��UbN=�i`��V����D�+Z�8
4JQ�*��+*�ѩI>��D�Kl��!qYA���'��p�YM
A������E���rw}"+a�<����$Z��Y=X���Sj!'��Ԅ���g�:�<Q�n3��Peka��Fm�ׇG>��)b�/=�x�=�xu�	KV�=��Φ#u�>�����ۅ*������g�n�p��+t�f��E��Úw�3)�����Iw�X��8mn�g�k�7\�.NO.�=�z�]��<����+�+��>�����S��;Etzz��|�[��q��m��wz����zDuݎػ�͝��N<؉`tk���o;7ɯ(~�=�__�9&��m{YᴴN �����N{*}��Y�w��:������b��ަ��ƛ>�V�o~��w���S�e    IDAT���xrpqv�YU��J_S��Gs�^_<{~���ܾ�����ow��~��\��f�+3��K�mSј�@ܝ!�3�5�7J�:����t)��E��i�̎MJ͐��7�3#'ӳ\�h��67� OK��]�:@��K�h	�����������S	~�-m��w�`�WcRD�2�h=T����Y���J�=� �n�U��4���j������g��NSmȂ�jT����x�1�n���*�P�+]E!�4N:D�43e���y?\�шC�����1������/WwA\^��[��{��Ƚ���G�{v�������;�}ʴ��ٯ���z������o��K���/�z���ջ��?������e��O�^����_���_���;�����wJU���a!�4"X\������\�V� ��-<��J�����C�v��y��n�4솑�v=��u�.������Q4���ٺbz�����$L�������1�Ma�P[79TՇ�o4o��I��1C8@#�<[���D�,~�����"�!|� U���v0Bj�,�����H�ՒĜR��q*D�X�2��jPo������2�)��)dv,�(�&�4�.����� J'k�X'����_�b�As{߿���i������d�8^��t:gH��7�{��y�4u\�@�b�����+�\4#D�_σH��_Q�UѪQo����(ݵ��a�@d��5��l�F9_|�8FΩ=���?�(P����E�ͥ\�խ��x��)��d�RP�a�h��LK��m�J�i�U��
��˵�SK�NcQN-��]'��(YX�C�)ם?�ƭ��W%�s��|��\S~j�����(
��F�~�jةk*d*Q���dʄ����gd����F��������?t�u�R?����Lz��I녣�V��ez�聯�Zj�e�:��W��=U�D�~�p�������� n���R����W%!8[ɛ5��� �����>4Q��!C�^+��7{�j���d+��6�Co3?���J����H�UpƔ�N��Հ>k���� f~1� p��`T�@����j�e�T-RF4c#S1��P�؊�ꐓ��G���VK�델3�9㈴!aN*�SW�i�mjz��%�� R�]�������>Z�%�Y|��1�d���U鎩f�h#�3S��,_������L���A�/W��������#�G0�CJ
#A!N�|�t!#7q�)+EnE����7S����Jd#(��X{qFG"��������P:H&h����D��Ç�3S�y5�3\.��*��v�\�Ȝ������E��,@�#k`��~p+!7�r9E�5%%���dh��l'�i�p>#eblQjBr9Ɗ.��5a�@;it"�evF�E.K	��p�B�*�~�$٭�u T�4�_	j�Ԩ�^KS���G'�#RW��Es e1B:j��C򫞦[T'ꦙ���B+*+}>&5����M#�2!Sd+�d�B�(N�3�d��_���?�!B���n[�Q�|dc�(�gV�0S4&T�X.���qRL�C�@��ߴc���$�q�I�"m�D���4B~��@f�M'+�:�q�4̡c�e���	A�ղ�Y��"�G@⭥\��~)��� 4L
8�`t^!WZ%F�W��S���4��B8�%T3�h�R��E�#�&�RL�lk�+
�h"�VʱRL�Q��62L�։U�aӲ��e�~��.B�KoZp&W�ǔoD3m����1�1"��`��O�8�m?e�[���6L�6_zM�$���jQ �3#aq -��|L����ٖ�vC�R��ǸK�I�[S�Ϝ)T3D I!�1k,\���� ����;�t�ρ�&�fj�����tآҩJ�$��K|!�uLY�NR���a��S�����*(?B�HI�$o�C��z�(*DA��@�����85oԧNH���&E�sv+�S�B�* bj�xՆ��@�G2�B���SŔ������IR�8m�7�X��BA�o��UnxEWgw�,r�-�?�iJ���2����Pz�m������õ6D�|���Ķ!&N����V��8����ʫۛC��3bm�Z��.���Y�Z���k7���<�y}��.��kἒ\�������S�����{Ǟ���mE��{'���5=\�Z��<�_����~�#+K��t ��Y-����c�:�����hܔ��G��{���s���S7:������<�z�쫧j��RQzsn֮�^���_�y���z�j�~��>�f\'�!]��-j�9k��t]{��gs:u�`�tr�.��+�������ɑ/ڼ8{���������i���>xt���w��[��|��������g�~��ӓ��j�s��n:�S�qZo���s;a��p{��e����m`u���|���t��K\��`I%��6br��8��5)Z�/�h��|7
1E���YE�,���ubD�a8�x��x`NWR�M1�� 9�yQCֱ�~O(�Ȫ(=e4�1}>A���,�|��!|��W��/6!u8ʦɶE��ؒ��By8_kB0��������t�� q�5��Z8�H�!�ZM��j��(f��V"�-B�J7����9�!1ed�VR�t���돬�L`�s�������~��o�����ë�^���~r�����������?����ã㷟�x��WON�8��w�������g�Κ$��+�WU�֍��E"%��Ŵ�$��dc&Ӄ��g^��8&�6��� @��� �k_�w�_�́���{��q�7"#�3:2�Ս��gǿ}�ԯ�s~����SM�����8}����ޞ���[ɺ8{���8���h�j˜�9�
KcJ��k#�aJǰ^4LY�BuiR�w�t��»<�=&�ǁ�t~򓟸��;i��1�R������w�I �$��b���[[
[�p��QӔÖ'�զ�{ۖ[����t$�wZ�q�R����=�����&=��22Z����&K �&��X�>�1ut�-P������1"�r	��M9d��BZ����B,�ƚ
�ΑH!���xM�"�')rY �fR{V״�9�E��1Y�@~"U4uf�7L�s6�];�cߜs/s�_W>��DKAE7��f�+��u�N���*䔥��A��m��Q� �n@� �zV"׈�tw��O� ��|L4Y�N:�:�p�����jbQ�,_�O͔��(a'���ZE�1���(k�R��씨����|��r�S�����@0�D�w�C�)��]�6U4N�Y���Vc���ȉ,d��/Tbǈ��:�M���Ux9�@� ���(谳K3VMM:�%�	�O�
M���'%�<���Կp�{�jl���u6��dt��N*J�<I�o��o�I�:��p��:��^����k=&�S�:�h�҃}�0;ǋrc��6D��C�^Ͱ�B|����7b�D.�B�G�cj���r�I�o���B���U!"Lo|��6͒�w;�����gX�ҥ�Kd)���� �V�2oF_Y�h�Hϑ��iۢHL��.�f �7�q�t��4AdH���A�����g�,��Z.��B	�!\e�BDL������+���ؿb�0?eL~+��9)�g �U$>��R�����1��ʦ0��1��l"�i�!Z�S+��K�2V���#a,D��F=�&%=�~��5�V�1ъ������j��7>P�˒B!S��M1�6N�N�54#ZE�o��hxdL�Nj ^�M)�%RP]��=!8Τ������Ч���3S�1�����BH�3\Q�,�9\!.�5lR�Hc��`�s
I�',]q�8�pc�y|��I��ǌ^���G&����'%R.;u�_'-�Z�Zb1gS*��l)�hӖ �$U��H=W���D9u�|Ӝ
I1/�����Y�D��X�a�1-Z�%B���le�)FH]ɪ������NK+M�D��$�z+g
4� �#�BLK��y4��oO���!&�h|j��L)@�Ѭ.�5UbV���􀖯.a�I�HGj�KL�����@E�Ɂ8�9!����a��M#gwӀ������)6�l�ZE�L$�f4�J[_�(�b+���w�*��!��&K4�k�����_4�p,?e�/�v\��\��[͐j1���dM ��UӐt�J���+��RK�)D.+�oj4��>�S�hV��Jd!>G
�����vp�4MY��%�U?@0CH(�V`;�7��l��K�W��Y����jJ"ݨ��%+�r�x!��9��|xhL
���@�|>4�P� q�
�8lS!:|��������i|�p�J��t,V���,mw6�ґ!�v�>��.&�|���-��I-?Z��t(@��)W#�S>k����z�r��� 5#�2g�F���'D0��#�4<���{�O��]�_���:U-��J'�\k2��W��Tz����l�K�+��h��is�C�y�z�`�+>52�id�B��Ҝ��oZ��� 4�K4u�MI7���~�r=���c�A�f�������W�x�f���';��Z?|	�n~��w����}\2��xtRo�ַ��G�!�g��˱ڻ�d������zJ�c�.8���g'�n�y����Jxr��h�#zp�s�/��yxy����'ۧ|��Z��ȵWNLMZ�/��*R�-��:]���X�GQ�����S�|��Z�GF-������v��	Ի��_�A���\��}��/�]�mn��z}�'\ײ���37b���c�V�}ɓ�Qo���(݆e���J?�;|�(�#wdM�aݤ���:99:}��o����z���雇G��^��?9��?���������_��R�F�0�.;T��o���ϟ��'��F�ul����k�tC֔����s��S�c��+"�r[uʤ:Ë�mQ�t؜R�R�ߩK-�)_J��Y��!R?Ï3M&D���%�LWM�E�	L�� ��!�Zy��_�6�Չ�DNvV�C�,DgMg9|%(��a�����U-���q��J�f�C6G	�m�>�Hd��u�h�[����y�#�BoO�D�a��E%,k�8��i&�k@�K)k���{x#��~���1	w�������׮/o�_]�go����������S�V��������ߺ��ӚO�x��'�~����7�?��{/>����G������)�|y��?8� �ԧ�Scv��gL-A{@��3�pW	��N[�i/1�ρgK�V��͘:C|>	Q��c[Y�p�^}����W���u����aj]?����@~9����*������Ic6࢝y��k�h�[�2�\�Z����h�K�BMT��X��0Wa�[�t�8��H�#�h^n�!�*R:f�~����ڗ�� ����?�%�3B3��48�Be��qXS#R�@VE�G���h����a4Y9�՚NL��iCh��6�tvj9drθ�BǞ�C��n툺�,�q��!� ��D!�tS�uM5���8�g�����*����,Ǵ%��k�G������@R�TJ�tTD�d���-S��3�Q ��B,�u��9Ȣ)sL��35Lђ%����к��B�e�΀���f�}�^��-yp�B(1>�Z��,a��͙&�f��2��YW�D�W�׸(R?|N�*�A�o��
�ԧ�F�U�	�Hm$���S�
�t&Ӈ9�L�����&0M%�tRq��
9�N�/�;
M o�u�r���2�*��g��s��U�Z������U�}�J{M@�5VQ��X��璉��}E��c��%K?*��J�Z�:kjp賘�e�1�E�d��9)Ą�r�U��	c���"�A�_��&:����:�l��"�]�&YB�Q������U����3���%�zY
�5S�)��`J�_V%򳅲��UdRu�P��[дfR�K4\���S�:�-YC�uP�	f�&��\���S����Nr�@���T���h��M���4�t�=:p#N�,YxU"L��k��:�����X&\�j�𘪌�?�*���������J٘@N~v�!��h�^!W{�I�R��M�n��s���l��C�ؔ~sPD�^�^�ʭ��ƌV�ɢqD9p���JpT�ܴ20��L
h���'+a��l��ǹ͖;��5 4UB��k�E+Z3���	q�|V��t���ӊL�i+L�qL%���ڤ�bV�-
�`�MJ%8��nY̦h��A6��D�Rl�(q ������4&N3�t>���_�]E&�X���)k�"��Si��o��6��,��eEMsX��l��N�y"�Y�YK�pj|�#R����E��D�(�����8��hY��B𥵩�@��i�9�q0��@��D
l�����S�S��($+�x��Jj5���PI!�X�4r�i���:��VZhR�|>��!��G$�TV)uk
Lg�>��W�:����lN�E���� ��L���� 1��B��F(h@:vD���r�y����;:9r����aVH�0�	Q7}ߨ�9D��� ��,k@�&:"��A��@T�n^4C�K^�0�mB(B�T���15LSfM+ԫL��Ӯ�Q��H8��]DȀ���'0��/�~"��d��P�)�s	��pL�Ŝ��'ȧYEV"�7�
��B���p��0�C0��1!�|`1!Z��lS!|�1F6���hM��VT���c�aMS��p)#�� e��Rx�9Ƭ%|���p�C$v�k5Z)d+�(fRS���i�DLq8�
7��**�+M&"�P��S�v�*5�2�cT�S�D�`-Ӵ�*DL�R���M��k[]Nuq��H����c�F�H
5���a��8��-V���X>e�ญy�N{�yݏ��]�C��Ֆ�lvGϽ�u���+2u�ޭ_�\YÒ�%����Ubmv��y��w ��O��%�>�;\�z�p�w��Z���%�l�uGq�u�o �����ro�&����e�����v�����v�(��*ۣ�#w^5�����{���۽�u���7����6�[_~����j��h=���,����;�^nG������G��j���ڏ���P��}? �;u��iAq�K}=|꾩o����_߲���Z�'[���k{iز���%�5�98w�6���r�Dw~.t�ZuX˧'�����ן����cw�/n�o}���#/?zy�1��^���W�[!��������7������z�!�OL�����Ϲ�zmk/���e=�J]�<i�0KJJY9p��>��O	!�)$R:¤�}�hH)��'��5e�Fy�4Z	�_��l�`"�CL�7U��·t��+v����'A�[�)�*�K�$�1t(�����1��xU�NϢ|W�h�Yj#�#HgB�z�Qbl)B�Ʀ���[����L���w9-��d�ڛVU��B��gw9�3VW���(��
oK��!���C��y�����ͭ�κ�yq~����O>ڿ~qwy~u��?QX�I����'��^�읫w~��Oο���9��罏��ů^]���Η��M�o|�-��|4�=����5}R����:\���A�(��!K�m�� p���zd�?��8�զ�bN����-ͣ�����'�8p�J��M�V�����|���� ]K� � �_�2姈I��(�2>CH��Yh�BZs ���&dʷ ��	��2��Vؚ}�*jt��հ�vP�|ҡ`T(d��Ȋ������c%��4�s^�D)�MS���D�ǟt8����B�����*�i3CTA�g�R�K�Єs����Z�AJtw�eM!���[6nc����
'�2�i��~��|�m�6Jqz����6��5���������.��CY]�ӝ�N?���C(W�a����_V'��0�uZ�ט!�����'�F��˒.�Ӊg�T������G�����;��!X~��F�V�5:u1�r�-$�*F�RH%^V%p4�O�E�e��C�+%֎�[��6w�dI    IDAT( ��[?��T� '۔f�!"�_Th�e�(����7l��,A`N�qjO"�z�BRF�
�`K��eun �B���+J!�B�uh+X4|�P�N���kÅ��v|�^)h�/J�f��\�]����������k��T]d��z�^}�u�n�iƛ��Z�}��U��ɶ�9E�m���	/�vLE5�h"��RD-<D�)<;`;	���b��N�e&%��+���+o�����W��Qp�=�9s�^4[�t;F�}�T�Ư�P��t���c�d�:��톐AD�XU�O_(&���e�D�m��j��o9�)Q���������
|x�rE���"S��(�Z��Y?"�V:b��F��r��jo�%��Y�ġ�4Z�Zŗ�tzH�����^�㔒�4S���	�Ϧ *�Nd���L�����i��cjDc�F*0�����&�F���"PH�Ω���W�Y)���K�PRr�P3�S4�UM�"=�t�[WRS�����RϜj-��@F3��\�����+�(��.Y[Z�j�FE�:��:�	r��W7�:�p ��9|U�!d�B��f ��VDp��&%�Ӕ#ѫ>&�o�D�i�
�!˔��>�ޔo��w{�աZ���V�|
@��|���'A�H�/T��L7�z+��]ԝ�5B�HS��=TtK]ʢ%�B�q�@��;}�׏h>2N��������S61�H4�L���1�Q�1;���Qh�ZQ��%��g)>��\�T���eUD�0f���T���D�C��D!)��R�D;��� p#_"�����	�njDG����eƑ��7pҴ�N*�,!�j�[TY5�H��c����:�Yk�ZѤ�S~Wz
���6Z8�L�&0>+�Z���E��#NX�V*j�F����4$f>G] 5SNV	C����L~ʕC�Y�����9)T4�t���r=��y��kcrS�,E��x��U�C�7"s�Ki	���SH�nc�V��a�!9���V�B�L9�Z#H�HMo�s:�Y��yR��_u�Es�I
ʹ�Kik�w{F �=���D+j�)�Ud-�q���G6�p8��!�Eh����@�2�-!�C� q�L�ƚ�mZ�r���D�R�ՇV:GJ:��kjt�-�5mQ��֕Rn��M>3$���W+A�j���Ȫ7f[��E&&�3�S^�rm㼠L���З�1d��%��`/�*b�fk�\��ҁ!cӇSk�!E9@�z�����+��iYh�|����Q@�c���G أ������Sw��#����g���norl�����~��ۙ�/��v��]�=��n@n�̺�蒢����ۣ�'�G'�%��,<?h���W�:d/�O<��iJ�x��ҧ�u�pϟ��=��/}u���U:R�ܺ�h7V۞�\?�����Ko��]B�;�['����^���Y�J>���ʓ�'����������]_^�;���ݗ//�髳���g�/�^�ܛږ�t����۴��_�mὛ��2�ǹ�>�g������Cy����b����靕��Z����u�Y[��l4�2,ǴC����n�z��o�:_�+{s}y}��7���_ܮ�����t|���������g�<�����?���gUm�`�������|�d'�:ջ�Qp���}t4��550��s����+�tR�q�jB�M���8|�jb���4�������˪t!��lHd7�B��ᷖ&Qt��ۨ�)�S8��hR�Sh�׉��b�J�S���n{![�	"S���Gp�*��%h��J.��.g�k����)�i7��XSjE˝�R@H�!��ar�Y��')��'>���rL6'�DR�W��5E��xY����O�+g?}ث:p]������W�7�I�����٥/�ܻ8;<�����d�����Ӄ���?x�G�t�ɋ��o=��ן�&��/�n�\���^}���7���O�+�>��/�+�� ������]�|p���.J�ٮrg��V�O��H�wV̹�B�Z�au|�fQ�F�S��`� ��Y7\-�[d"n$�NP������������|�i9^��5Pt�]SZ�w��Q�_
H���!:d`�b6%�m;8�fM[0NY�!d(�7�,�`U����,�VY���*�����L�z�X�#�,�pL'����sFAԔ��,4��ب"j����w� �;�B��b����h�����]��И��p�����j �U׊d'�����czG4���C![�OD�BN*75ݏr��;;�����C�#� ��0A��,~��h��B�B�eV�)D����諘��Z��h8�D�)Īe�%�\ �W�f�Ji`BD�Gl�E�p�l�Ƣ)W�R���s�rqB8��a� ��h�9�5o��?!*F�i�"�&�J�	M+]oq)�:��n��B�F4Mr�� ~U�B���;!�.,)� �Ҍ4�бLS ��|�/�c��;�L�"��t��G0�ME�9���b���D)���Mw�,� 3@̿)]�)�'dxa]���t%Kz[qM�����KA��`*1Y�	t��[����SY���BMirLQ���3�B,�+jr�@9u\������g�n��Z�Yy[jD�02�,!�x����e�����z��b�F%��i��iӶ�k	�Z}�Daq�X���b
/kQ7Nk��HU��!1G���vS~:Ô�2w�H��tu�u�8�X���e1����p���t���GPHT����S+M�F��'��ac6�Kp���Ȥj�5b
�Ӂ}B�+s�z����!;GDzY�|%K(�U��c��AF3eY��q75L�~�*��D�ɲ�-�(~)���)|����,�P���Ͷh��9U�������U�Zh�:d��I�8!����lj�8�*���P.~�K�Zp���6e!¡ƉL�P|v���R���^Y�t8�܆��g�M�68�6pZ�i:�/p�4�1�$�Ҕ��2�#tz��E�	��.q�o
��O��m�Y�:LMiC.����ZZ>N!8�����\�h�t��j�Y�r���*2\�`���ʂp�Es(M���0P�Ԩ���[ N8q
.�5�G��)���:��F��U�8X])D(�DF�~�e�8V�����tR��)�ggLq�uU��{�LS�(�t����톺:,e���)L)F�VD'�,0�����L�8Y��
�5���^��_ݎo�*���C���"�k@�
�ሲBI��R Y;�ix��P�B=�T"r�*���i����Uo��B��Y�\c�Y><0�t�ì.�Z{�!d�,	=n�D�Z�o�\�=�:�4�X�e�������B8�t����(�B���I�ހ��9;�<M 2fV]~�H���N��B|��5�i��6Z�Z��.��V:��|��g�%Q"�F�)��t��U����||�(�V?U5�Q Z�
mJ�yk�&1kU��lj�S�$���@Ri�b�!?�DS� �,��)ʟ���O���b��>Ь\�5G�t�BJc�w���\VL�eq [c����2| kD� ���]��|��M��Gj���U�e���uŒ��T�E��T�����J�R{cs
�7� =q�D=�EшW2 ~%X�/}�P�R"�MIa�9�������>=>Zm���O�]_xzѣ��m'�s�ÔL�l���k���n�I�~#|{br})����dp ��n����wٞ�ݸ���z�=�K�G�{{�	uR9�7��z�֛oN|���� �Jэ���N�w��͕�+�g����ƍR�ѭ��[?��~�M>�t�"X[$��ڗ̺ǹ~~S��6�V\]����Nvo����l�����7���o�]�~��������߾�;�O/_�|����7=~��w��ՙ;���o{�Ȩ�� �_�s�X�[�U�����9>y�6�ށ��t/�������z��O���n\��9׃��W�ZHM��݆������ֺݶ]{r������NN?�����/Μ`����o��廿�����_~����>���ӓ�_�yy����o��̝絙��f,_]�a���j��-��vp���q������p'�#�f`Y�k�ڮ#E�zN�v���n#��%GW!�8��� MU1R�UfZtjq�ψ\?�ʪDm!��tL�"!��[�2Bh	�&2�A���`Rq�7�J�)��,��ǇǬ�D �)4�����X���JjՍ��Ǒ�DLN`�	���2�b� �~*���XdK���Ȗ������V��!�ïJw(|Jizt���cW@���������Bv�?�8��'���?���<N�_�u�������W����ݛGo�k�7{�������wϯ^:���|�|y~�@��e�>��,k�ۥ'd|�������5�����n�h��8�E�[�m��=g�[$B{b7 ���6߈ ��F�ISL����{N?����@O��|�'�V$K��Vۇ���'��5����QN�)<���f[v����J��7fU[Ė��-���ՀD�k�cY|���D��XEM��
��|H�r�XW(T���n����c9��l�,+lCj�x;��fs�RL|���7�Ah��,1$>2~��2xۂ�%jΉƇL���:��'�-�5Jw&y�[�N�n�xA��_�%.��m'+W��4����Y����qt��H
`G�ˬ#�@S��Њ�W��u���S)N`g<�Z���M�`�+�MVi#����e덭79ܺL�-6�h�R��8���Vc����r����r�B�𵑯��q���ᚑǯ�tLq��䤄jC���h�]7T1դ!
G�[���!�x��9D���`��g��쪨AVT����R�DL9i:�EE!h���� �IM�ۃ[��Y��s����@�vؔg�-R����&���Kh�]|��(����4��wJ���?wG�,A�}�%������;ﴫĥ#��4��΁�Vmum��Z8���8B���80>2<0����o�z�[Fbms�P�c|M�J�q9b�-�f$n�.8.Gv�6:���.o�J���O?H=G`QM��I '5�@�Q&��OQd���8������|��S�%�?j	U7ASY���\>YG�]^=���Z��Y�!�cph�BЪ(d4e�`�� ��QK�)��il
�E#W���Dj)+��n���8��#c�CY� �(D^�nR�HIG*����M�cǁ'aW����J�,K
9��D�8-A(���-�D����U�j .+ȧ��In
4�)��v"sc=��I��iRZ��ъ*5u���g�[�mY��[�~��8��B"P�g�҆,!#2����zr(��ˏi���R�{�,|aR*M�N
��c�^�U�nR%�1���B��	OVKS�D|~W8�N�5�m7X⁕�@G�8_!V9��"ǔ5)���|������L�UQ���LU�JG�k��,�B!������ch�@3�b��BM!L��I���)�B��pBL���n�U�x�P˴�k@�J7�����UQ>�i"���Ư$��Eˊa�S�j��n	YFkW��Eb��"S�+�A���,��~��ɇ���Vm���du����*fLH�i:��*=��Y:
�h*dP�K���ʝ&E��?[iQ|�*YH`8�i�N�@|~4~_�#��$e��Qk$(e8������ ��M�a�hKĬ����OQ�S"�2�T7��Çs:�l8�ч�j�q��8���'���^�-�Vj���$Z�i�imq��OA���*�e?\��ȭ��QKD:~jB�L�e�����s�N'���S�k��~)ȘFN��J���L�p�]�r���V4��J��Bv�pS"���pY��P�i����hV]"�):�mE�,~�h�éĬ�Z�V���7ꭶ�8��.y��+��b7����vf��8f���4�ɪ6AQ;�/��o!B@N�&]G(�ᵍ�j��8��Ys�`�-a��)T��0��w4M�#>Y8����(���*V�)�!��L�O 8ח��o����8y[;��Q�Z��f��)�*��m{Ⳑ�}Sn+�}�*)Ojz��P�����C����ټo�=�U���=��s�Ww'�M�݉���h�=rg����_��E�����x��]ݼ��#���s�[�Ψu=�����Nw}����o1[h����-�~�s��P߿{ws����݅{����������y~���>M^?�����ۋ��g������+w�]����3"����{������
}y��d��t���MMG��a����٥����\��^[����v�:1:X�A���e����znD/��]������7���g~K������N������B3��g�~��O��ռ�����o�=}�-�{;���S;���3j�rB�u�a�Vu�/j���a�tv�DD�Bv�Ctt[{���,��#�a�
��o�o�B��E+M���tA�@4 ��#��ge���'��6�M���#���	hUω����V�p�?�FK�~ڨ�F3|v�/*Q{�iYI!s0�J̎尻ʘ�m2���ɯ:;`�,�,��9Ӑk �e� �4�:�5��B�Z;�g���φ�^�K�ӕ9A��w(Nǫ��T��>��^��������ə;�)��˃�s_<}s�����ߜ�G'�}퍯}������;?�?�|q���]�����������4��7���C�?��?p7Gi�v�������r�M]��k�խ-{�D c��5e�jpt�����q�[��S�YG�w7tS�?�+	�=V��m���N��yMb��-�b�\`�U�
~M��Nd!���4C@���E�h����H٠C�#���Yb�f�h;���G�>�|�Д#np�9q*YSW���oA��*���h)_��mK]���
�98E�OŦ�'h� ��p�An�W��">߰�8b:��qq޳���!8����$/!/:p�A�T�;��4��Z��h�*'d
��×X�~%����UuUtV�8�l�����1Չ��D��� �#RݚA+��7�H	I�OG?5�,�>EkIe��*�
'����� OQm!^����'�Z@��a���*���x��M�\n�����Jx�$吵��t�5�&A�qN~N�p���@�ȇ�>[:��t���@����X����K��݆#��5S'�r�U�@��8�rm2���\b��h,���Mu�t�R
P	4��M�$���{:���d8�l��J���|oNޫ��T���*m�M�l������h��1j8�mW�.���hm�r�%?��I*�i��X�)�1���G�5`umK�Q���?����?��O����?��(��g?�k	Y��1Y�V�aO�%%�(��CLM]��!�Cp��Y�DY8�r�:�pDU�ࣱz�.���1ٺ�+=YY�F9)����a���UY|N�q����C�Ч	�a�XN�(��(1�5< �:/��@�VK�@����˪:ۊ��w���FXr�� �S�	���Ւ˷v�_�-Zܔ�.&gwu��`��h
J�?Uu��UhLV%��T:N)��k�T���f8�e�Zp4 �ۍ(_:K�&�Kw;�!��d�����#Љ�R��h����CY�R�,�(s�i��X�,!��8Y�xy�3?�I�g!�h��J�P�s��DF3����*JQ7�p��єN�40Vl���@��u=�MzKm���&D`e�M��0ŏ9k�p�8��`��.4Q �H|�P|>B����A9�SEӆh:����ʱR�2��v���z��F���������Ue�#�w�U4)��dq���opQ�ܖ3|��=[Z��>���E �T���j�V|U��l`��n�i�5��9�.сT"A�W�*���Igz���,>�4P.��Z%Rݐ8���>�ED"��1��N����B!�ΥZ
L�U�X%ۭ2�
aJ���&������9u4$��vn����8��ԕ�\���%�B�A    IDAT�˦Yu>j����*�a�VsJ�-DAzd���ώTL:��?Ҵ��R��u�L�Ѧ�V��/eU�)�I�_�:��f�ꦭ�N�i����Y3F�ZԪmQxէ��I��� $�7F$M�@�s)I�s�M|%<��8A��42B��J�<QC������i\nY�zS�4�JO:����n���LJ����U�5#dj9�hD�I-^W��q�	\��W�8r�ea���B 8���B���8DQW'_ȴ������C�$�5>�1�!��ME�BR��!����@V	��f�m������}�]`�n�4d�l��Є��Y��h��p���p ���^���!��5�iojI��5@��)wQ�d[���UQ���>:��	~�у}T=^I�'�6��z�l�9��X�<k��#\���ܛ����CA���i�n߭}1����ŭ�+!y;oW��\Z��=9|�����O=6tu�@ܺ���M�޹�K'软U|�I��׎�<��ʽ;a�ۓ��խ������<Z/�u����Lǽ:a�Id���:����\w��=V��;��7����>������מ��x�Vߩ���OO�|z��'�>q~v��tm��Z%��:��iO��]x���޹���]���g9���/�v�n�z��U�j�|�o��}pw�����;c;l���mk9�}�h~��W�ao1�ke���ӧo��o�����<�쓋W�����7�~���޺���>=�p��O?�ŧ�����GO��������N�~����W����Q[�X�[?|�C��b�#�Y��#[�#k���	EX�vM�Q(�t����/D05~%X�P�Ԉ�3��SW8���t*���|�@��Ser�B��3~U�O�*E���!���,����^k[�a�F��4�&K��b:��e��1p�@��SѪg��5�.�� ����D���$}L�09�r����e����Qe��"TÔ�,�;"�z'r�mO���c9�J�?�MQ�bV����V��t����}~��{<{������/\|����{H������ϗ_���������~��<�.>[�����7���h�GZ���B��{��g�g�:�����������������$���R=�PW@���Y5p����w�M�ِRЀm�w+|M�@XSj=)�	�3�c�>��P���G�C>~js�h}��`�� V��'TS���w��.��Ye4ׄ��H�R�AV��O�p"T�7�ZB�^�/�H��3"�=W�2��1�8h5'�Д��D�E9�T����Д�B0q�N��a[����r��7R�������%&eZ:k`��R�`d��QU"Y��ajQ��s�������+^3�݆�Sm��ѭ'�!Q�v���0N>�ُ~����q��itb��
ѷ{��%C]��C�U���ꪠ�v�霈���:�UI6�f�,�R���0+A
�舣���Պ-�H츰��m)b-�<Hߔ�鬆�KAT�)?p6�%ʵ$��I�����q�lN��F;P
k�Ր��D���Bj !�f,�xE�#D'+N����sY�KI�,�G�G�M����rDl,fH�lJ�i�)�C��t~��p�
n.z]б]�9�@��u
����W��p�������������B8-G?^G��^>�Ԁ���8�%�+G\��.��ӁӘҁȔ1���dۈ�VQ�>ã�o �W,h BG:��-��Ǡ�\4���*1�NE��+%�Ē����&�(p�����mξČ,A��Pi)�A�� ��#;-E�D�sj�,���"�'���?QmD�i�~�ݢ�R�B5����oj� 6�+�n�5C���t*EV M}��	��|��5#�hC��V�%I|ח/]�B,> GEYCT�S���QzSQ�tCVNY�,2�rl� �� �OVR���CK�)��mZ��b�?�U��^	��i�O3��8h��6D-�_'e�lS�*hI�ҢB��i:iF.��1f�|:#�lh>��d7�Z/�~>PE�D!S�Ę���4u>G�ט(�h��F��h��4Q/�����2N;�"(g�G��3�(����B!G�*�"!5�!b�)'��Ӂ������(��H{:�SVb��U�q�[/ܶ�J�'�Ju9�,$k�8g49@ug9!��AV��F"�Ѵ�&��S���!�DFh	U��k�%&n��t���	CV��L���C�'e"6�1��0U���,���5�p8�LU�%~�"���5Ŵ,f�88BR8t8��r���s�q$���VEn�SE4��SB4}Q�*�l�_�m�SE'�ȊV"�D����M��Z�Һ��;vE�}����US?�&|`j�!9��W(9�L��!�h�BF>�)ѕ0q!�(������oUꦬaY��9z�	�
)��o����g�(�,~�ᬩt
��C��E!hOz)@�Q.��,�B�j�f�=j7⳦I�Edz�(D'屩�sj�ݖ�rɶ���+����Rԅ�V���Y?����H��i^
��tEM��Y��1Yr��U4�Σ�G�i�'�@\���H?��Jn�k��Q�i��*$�\6�ȜX9���rq�m~�ukj8	;�|�{8	����r[RV^�R�)��dt�||߀��t7�?�arZuN��+�&����5��$Ċ*����"�Z%.�P��B�ګ�!�ȗh�E�R��η������Ϡ�%����頻��S�u�&��n��=d��#�(kH�)���(gE�bo8믍�=���ڃ�l�d�g4S�8�@A�����!��J�M�ãu*�E��0tg�zs���nm�_�\�@.w������<�:\+��?��2���vJ8������MH�OO�O�<yy~E�G��!��b=��{f�����r#����7��.}�r��h����չ�ۻ����c'G�7w�~쇭�n}!#c��zv�KÃ���5���s��ܹ*���5�_�;�;y������˳���)����O�nϟ�<}��o�}��ŧw�� �����鳣������Zt)m��~<=9RΛ��#� |z������7,ד��L|�[�+|���Ih?}�.ڇ>��������Ж� �c�����O|�����_\��ї�gg�g���G�%�kO��]����//���?^�ܼ��7����[{O��^~y�F��{w/�����>����z�@=��0~���k6|��_��'��~\N|ScW�T� ��϶!l���4X��.l-��rU�6=�ּ���Y)S�.���@X��WDͰq��,&P!�iN�q��B
MY�рh���(sr�9�J�y�D�Vuc&�ߝ�1�j� g�z���Ld*��/������g��c �"�1��F̐rTEc���4�xR�~%A3�B�w���|�ڜK�ΜVZ���JW�=9y���Q�/n}y��ѩ+�������w��O�=?�ڻ;?�zq���W������u�㋏}`_^��9����{��-�� >�5�n����/��/!Jw�кt�Ї�:7u|��{7��%Z�UH7�Ү���m�i;��_�j�@
��1op�s�¡��z�w���0���/;�@��n���>������jW�P�Ю�!S8��)�3[+E���9=��l.1��,>���Bu�����Bl
�����#*�aR1�V�@��R�?$�Q��?u��*��~�TdՒ�6F�5!l+��I�#K�'�m�>2+�"�Bb�!^�VTTz%L�����y~Y��������
��m��tW�Y��+���N!/�����s�NB,J�*�$ZH����I��,�e�""݀h	�g���Dd�w絛�^�����(�����I7�98�!Gͫkp ���y)�C��+'�O�/�Z�ɇM��h
g�f�N-n����Dk P��1k5e�Ҙ�*�������Q�b���4�'��[�r�g˗�J��E��`��z�R#�Jl�9!D�j)h��
�����V�P�h� �򩩒,�*j�8�6R��ag���m�\Q�@�p�ԥ�u$�4\��[�����ɟ��d�pA��^YhnFWTu�� �.4S�.W3^S�cl_8D�YB�z�Ji�u�����Ū�y�88��
�'��h6U����)@�i*�Đ|=�!N����f����w]�c�-B�'j�m��R�BA�OPK�h�Dk,�����Z��*��f�����v�%��h+�g!�����	�����XMo_�_���8t|A��Q�}tw�c$��o�l&D�%��l��Sі�J�Յ���"`��+QW�R��8�)��w�e3e8d|���-��!k ��
�����X�|��fJF��I��:��8��X/��t^)a:l��bj�n{H�i3��*�$�~CbY8eU�8��-�Q`mN���j�S�D!�(kБ���W��+,��C8�rYg����r�8�H�(����^zpS8��^\�O'>dN�Y�t)�A��@p�ʅ���δu-e�i��u��b��Mn⦉�RL��Ǭ�tJ�I [i
B��ҵB�f��
�S�Z�[u�,D�&����-�	l��n����-A4eu��T�������U�bJ488�)*�#4�I�2BN6?N��@�=�"�hO	R��Y� 2��YV%��&������@��o+D�#+�1J� ��lc���#��pU ^,�uX����/�r8V"�5F!?�B!�ZI�X�uG6���I��%�(
)�~=�Y`{¶!���Av �z� I�_�(��i#Y�a��bH�'�N��pJ�fp���5�T��B���˕hZ!�6d��n��)�D�0���m��r��L��t�4{;��K�mI��!�B��R_
�,��xg4���j>�uq���VA3�t.M3ā�5o�a�L�0m�� `J�D h�	�W�P�%���|6|�~j�UR��89�%f�Se�4M�R�����)K���ʉ��G�ˑ��c��c��'�tƏ�=�V.�\Q!� N�i(Toh�FxlKjN��5�@4����hį�Ze�"t 8hL�MI1�!�n��t�������&[�i�?\-c�ꍆ`�J7Dn��[��.�=�������w�˵j��ԲD1w;���	�P����N-LG�)Y����.]�5$VB�i�����,�g�r��2_W|jF�d�G
�]��O4������~��s�^�^�7WRY�v��w��<+�[ߣ�F}�{Y��tߒ��[�[����gr�]����^�p{�����+���������{��;�ƽ]ώ�7wr�#{�����+����ӣ�'�������y�R�~��]��_^]�d�Z�6�Ñ�3�}������Uv��_=;�`��y�@>;<>9<�?��W�x]�Qm��ѱ{�O�n.<�s��˫#�#��l{�g��9�M�.�z�99𳚫+_J��;�7������L�s���������Z��f��C�m��y�7�� ���������������_�g���9>8u�����ӏ�m���b��Ͽ������32������>�[�חg��$�կ��o��gN���������v@;���!w���1�)��7����Qdִ�4ن��P��q���{U�+Q|CA���o5Y���Lkɔ����S�Մp��I�b��O-~)��J@��:4��ѯ���(����W.2YS䦜e:||��`��s�n�0�z�7�,dJp�ȉPS-R�|c��TwlL>�z�p����9�I%B�������pU�T�@��g�0ҩ�gII��8&e�!>Z"���J`�h��"�]�c��O�ػ�_Խ�<:�{�u�$}D�����G/~�����>yq���Uk���}WWg��{���w��IiCQk����y�����CB�q���LH>�s�����u�R38��C��	'����ԡ8�")�(�Տ�����*�Pp
�O��O�ҥt����-9b��ڞR��iF�����̼�֫%	��5*��b�F�K��e����i�eG�#(-�ID�h����#K��uk&q�D6e>B��wHl�ϑ������ig1�Q�~���[�T������M6���R:��
�|x��@�C�19����ۺ�泶���a�q&8��[N&7f<��~����i�\��;��������TA����Y1]�(�`E8m���WŢ ��O=�l�T�h��\cj�2�C��l!	"p����ϧ�"�Qq@W���X��X�kL�>@���
Y~�|��D����i���h�SWp���Ek�SE�@��_(q���$>�}eEv�Y�A�R����xEY�JU���+Tu�:T�a �������N�)��B��ƪq#P9�!��TB�p̦�C��,ˊ(CTV���e[B{4��ɲ^-��y��w�?�����n&��KFT��\/��}�{���+��w#���U^����������}�nu�Q����E��z��VǶRA�����.˔��(�͉i*:;��8���FjlD��.HG���t��"G��6���ź� SC��>N�����gz�`�Ei�*"˂��v��|gU���l��E��"]�B��D���� @���ֶ�eN���M�����?]���o��Y���d-���)��8K]�D�B,>k��0%�h��lL���]q���-�h�a
�U�4谦��/=���5 
�)c�܎�#�NC��4�iT�����p��2-�i���I��$�c�z�@�.�P��g-@�	�#��.Y�R��j�LX�Qn�N�:t^E�'U
Ѐ8�Y Y�E�ȉ�	�@�h� �@㔢VR����&(W�B��;V-xͳ�7uR��X4LS~�B@��Y�F�q*��J�Q�� �@ck�SH:�8���Dc����2q����,��	rX�e-�&�j��҈���&�`)�ө>N-���jLԘm��/�YVQS:�8��H���5	/�S���9�ҋJ1��@4��9'_�t�;L1+�Z�P�
%�J�(����EA��*r ��m�Ư��]��J�B�VKD&E�]"X���p�pj�i����c[]�&�,eH"�k#?)L����5�¥����[EL�S�c*�V�5��pL[5ĨCN��do��+�"L���R:ʦ�R�hqX�*@�R�MR8�@>�1x�U�^b}�7Z�c�C�p
����*�5��\	�a�F� �n�کb�C��%
,qk��ɺ�&K����u�nI�=�B{l�����w��pC���`"� @�ݶd��-uwu�ֿ*�i��S��|��\�=���ޕ8����Y�4?���ʱ|��]�� '���*���/�T`),G�P��#�'�C(Zz�����4��SY�Y����rj;))�(=}�f'�Ӏ+Q�Ԅ�?��[�L�	a,�5fgߤ@�HA9����D��'$�v"��z�@���A0��c�[?�h�pL:UA�4-�Q��L�(>?'e�"��8U�a*=�D-5e1+���zD��r�G�\!8'>�2���Ⱥ�׆D�v���U�7��\�`j.��ϟ�5���cI�غ�R���ޯ]]�CN��d��@V"_.<^"~�p��:j,5!>��az��/��Ct�����7
l-&�f�����>�F�'k0�k���t��K��(��88v}�8�נ?����T��{�*J�g���g+=�<����W�z�����z��������V_��N*d���C�}���٦��7OG���3k�9��c���!�|����g������=��Ώ8��멬��>}�Y���ȤVoO���i�c��'w�g�_���{���ϟ�ݬ��9�;Փ���;Ǟp��ٵW��v�MDOαs�����Q�)M;��7>/N�= ^��T���O|�RYQ��V�{wo��w��s��b��~��]t{A7|u-MȢ,mI�_a�B^���է�������?��+�_|����'G�����z�������k=��9>9�@�޼��:=y����|�ӳ�[\q�r�8    IDAT��u�V�k���WuVk��k��)��� ;c[y%?V)�Tn�E�eߺEL�R9�_�j"}p��L+m���-.k5����
�MǊ��q���B���ڿ����2��k)2�B��� B��R-N+
WHJ��	t �ʲ�,�(���5F��r�W��SȗX�i��L���h���ȭmޘ��Nz+���/;ȭ��iY�|+��X:Ǩ�d��G\"Ĵ��� ��G�>Y!`"��Kx����x�'��������ʛ���˧��?��7��[Ｚ�'�O���������śW��j}�އ�~���OU��7m�����Sq����^M��j�>� �ЧP�dYl�Hp��i YEY4j
��R�~ZC ��Дh(w�6���NE��T��t|��ަ��?��co�z�t�m65��x�S���IB���$Xc5uw� ��F��K��+!�2���^tqti1�W�{�ҁ�1�u-̐HD"4%b�>A4Y�dD�h����R�[>)S�8��.�c*����%�O��$�|�n���/��Y��8:a�I������B)kn�e��*e���vm�*Ί_����	���ut<������H���+Ob?n����c��R��U�Y���,�n�r[5D
C(���� K����\�� ���PU��Xc����'Y�\{/dj���"�آ�ytpt�I�f�B� G� fSn+�:��rqL]Vt4)�M�����&��dqH�:!^��ɟ�*��� ��d��BZ�I�V`x�||=�)��+�.��i��� ��1unxm �BD9�P���B�B��Ԍ���r�
qpM�D0�@4��Pu��h����������>��"rc��R���i�7g���:q����D�^�$���̱RE�K'|
#H��~L)�"Kc����Ϫ���r�(L��@�0ۥȢR�� ���pH:Ua�z�))�,\����?/���4mud��[u;"|Y��>�j��-rqI�+g%jb�YL!N���Ri���ETH�J�dYHg�t�U'n9|���B�|���Xs<�����5� ��	Q1M��vz �l��\'5U"�h�����R�iJ����Lg*
A����r�9چ�n���G�!j�I�0eMK� ��5rⳢR8��S#�,��X��C$:ʔu[�{h�L�ŧ��q��A!~%:��X~����hC:$}N�cg�[EL4�����ڋɊBt���1e	mi|82G��>p��Ň�X
���Q��TTH'��Zќ��S���1L������@ґX'U2��Zr��@N�}0%E�>KD;,�c:�D�e%�Zw��y��8MKL��I$\3����p���P"2�׌r�Ui�����`Fc�"������)C�9�"�'�4��hǴCY�hBQ�d��3p0H�JDH�5�lQ�FS�֕�%h�Du'��=�\L��ȗ+�H%p����� ';�8JH�Ȑp�������e#�G�g�i`���嚎_4�,�B�p6�(�mN>[b)���5�"@��ON�b	��z����a#8�;L~ä��]�,����8!��ZRN�l�h����ɩR|cB�P�DxR�j񳜺�HL�%�&�BY�K��Yi>��PK�
B�cP�#T�D��W85Fs
��d�9ӌ����!�ϊ�UOg�� ���	�S��ժ���h!)�����,�mR��98��c�Cvd ;{�`m�S�����M�d	� ��K�ş����@��fX8��&%k�>.�r!U��L'pC"NߵF�,�~éO�~��L�z��~���Y3�c� 1�k�MgQM�ߞ�a \)@
���$��[��4#}`���P�i!S>��\ �PR�O�/��	7�T�5 oٲb�Ⰺn���cΘh��h ��D|��F�C�)�ϻL�N�&T�}�����@R~�bs0��@f�R:�
�>}֛�p)�J�8�!
��0pJp��UHId�EM��h�YS����/��������!��cߋ��KӾ��B���r�6ן�\��y��x=�t[C�7��ժ��>�#�fG�*�O:.��S�x���/�����)��͓gg�y_���v�sHͯ��&�~߭Cs}r�Kf_�yvw�{#uƬI��{�G4WK�Q�^�:��]OÁk�HZ�:�}���}WY��g7}�ӝ��J�|P�b�E������ճ��������3��.oU\�f��^^{����g;}�=r�2�X'ם��zRz�?>��q���=[���*v��O�$w���z{��#�~��S�������h%.�}���������&����Ͼ�?��������gwo�_�\����D��w���{���ٽ������`�^�_�^�h�o~��W?��okW�Z�ҟ���D.e���5�6�/nЩ&���!"d��a�%���ڍ4���1LQ���K�S"[�R�A���Ԫ"ASC��O�ӪP�Ej���B���M��(�������x;ȻyU_��}���2g�|]�h9l�&F��Y��QIq��^�ʭIN~��ƟZ�\�Q�� 1@οB|YuR:'_z��q�h [n���,���t��I8g:�U"�!�,�q&T��X
���Z��C��U/@p�~_ �(�Gt�WB�K����û�ח�����<ռ��z����]��ts�%�7WG�Qő�9b��|^o�Q(M�����oӛk��<��x5��a�z|�I���)�Rh��R�Y�8����:>�,m�5�,��
�}HKvz:Q32\?�{:ѡw������� ݎy/�����O${L�	��۪j����Xy!�䘊qD�]���%��Y<���}ݫ�dϟ?�W�A4S��M�DQZ+D�6���gp�M�/��Jl���NY�/]Ȕ��7��)��Fˑ�G@�P���r��M��ÏOS)6�P
�C��W��6�)`�m�9iG��N��-�������_��_<���������&ש����A���7�D�y���g?l�^����WB!m%���]j])S�k  �աz��\~{&��\4Y�| d"�!�D6e��8��IS

���D�/kZ���C=�LLkg��m>\o��,G9"���b
l��@"��O�HД��U�J�$8���Oy
K��>�@ "ȶ|LULu5�
H��Bu��i�7�!4��8��q�# �8��p4ƒ���[�ۥ5&� J�m�!�3�8�|t��u��|��Uԫ� ��\-���qM�r�����qk�ߔ����r|d�?���+�����`�ՉA͍��+?@#@Xd'���Z�뷝ዪα.��(�6j��MF�Mh|d#eL�rJT�/j(��#���4é�$�`!.|>��sS�|�6��|4��i��m�r[Zu�R�S|��uhj�E�G�|�@ZȀG�N�MT�;R:!���tdY����RK�J�L�7T�Ê%�%�n'�4!��Pvi�)����<��ibv���D�0f�%�����a��E-δ�gm�+�i����#�4;4!Y�7wE�2Y5,���h��p ��i3�)$�4$>G����!5��*։�e�T�O�*���.��zA����YR!�Z�n:њ�����d*��hՇ ]��@��1V�hH�CXQ��@)vlVGn�Y�!:[w��`RR���Ň�k)|N%��Z/�ZY�iI^]QN�V�tNK����,`L�*9q
�1S�P3:4�h���ᷮl�Z� �+��Z�:��"S@�ԤۂP�R;�W+{��8uX��&�Em�fJ�?�B�lN{H�OhjT��� ���P�,���I�C�(%�">_��$�t����z�<�@$JOg�%ZkZm�pd~�b&�V��-]�%�9�9l8&'?>�
�(fvhC�c�R������@`Uj�C"���E6��J�hBD�䨫�8���`u�xuә��jm� +G$�h[u���j!�_�����u�(�ހ8���2���0#���pU����Ԙ�N����f��JW�0e�Z������M��?ͦ|e���)�#�� e�L!�!qj�.��C��ٺ-�7o�m� j��蔠PK8NY5����#�#�g�i�*4�@�hHQ���Dq�N���[�h�v,FY:�t�O"�F�B� �q�gk�8����<=s�D#4��u��SclQxHKp]@���
%��O�T)SH]�Bin���X��~"�4��81q�|�p�X[rS�>q$I�1��h x'"@Lc'-$'2!6|rKdqڇ���#{(�_���`���;���h�o����kQ!�1�j[8��߈1��r�O�5�֡�o*�E�փ,�_pR&Ro�k���dE�HO�*�����S�R����+dL��:��6��T�%�M�/���ה�#eJ����9�������{��7���YAo���6��*���%a�?ZI�����3�1�>�xtu��cW�W>mtr��
�ٻ_�������o��������z�5��Z�:=:��x4����ϖz���>/)�j����_ݝY�ÛBj�xd{��S�©yV�O���S�t��ԓ��קO|��z��=�|s|����/ͷO.���F;�>��+q=�F8;:�����a�!�[?���s?��
\����5��Yό=K�/�׾y��Y�g��� �y~Ŷ�ڎh��	������8	�<�T���؉ww���^߾��ӓ��'W����_\�=y�a��͹��d}��/���z}}���^^�Α���n}��'����s2��'��]������i�1r椚i�t8А;Vb:	F�^���e�}+dQ��9�%����IES��c�Rt�-�EH��c���Ǘ�,)'�D�@�-Yn4�WQ�8Z��IM�T(~�|���E����qܩTI.�d��U��,��Lb*�g�FSN�B�t�8)#�f5��5Z��CnjDΑ��s�h:��!����78R�6G4N/�Ҧ�^�;��H�D���yk��0ݚ��eΎ?}�ˏ�����''�<{ߟμ|����X�ֿ�p���6��Hާ$�Q?ڠ�-A�;+�+!�}�>�kÛ�r����W�ۦ�W�y��kX4r�U�cM��|E�p��l���*v	no?Ji9@QO�YM��~����Գ�c���o��>Q�F���?�P@��rPs��-���K�v죹Ρʧ �А���F������!�}DK��JSL=�	�D��t� h�i�u�U����F�OEvm�%"�������^G�(>Ĕ�V?�N�:�Ǚxk�/�f��r��2�2��&D��\S��ɲ|���7��O~���E�Q���~��=�����%;�=�q��&);��Lo7��d�
qd�]G���" ��
J=���B�7��Ŕ�~JW�8ܑUW�.�p;+j�Rf!��Dv�%HD�I��Q�&���Y ���2)��T���fi�F�|Y��OИN�4Q>��ڍZ�9��R+�&-������'�C�1�`�㞫4��h�6Y=�"a�g��*������ԉ����;��Z��D$Md��^9�RCPn8GD3\J�������*R�ZBxm��J��ju��:�L�U��,�e)���+J�1��E��@�됫�?2@n���d��jO��:}�Q�]��	:%ષL��Κ��j�4� �CD�!*%�E`)k�eZ�8���H׭���09�	�Ӟ�9��7쌕��BKp�H�ғ�k����F�v+B#�����E]hrm�4_:��#'e6��`�YC�C��8��r��фXS�ශEYS�t�S{�L8ۈ��3UnԜ 856��@����ajD�j(8�����#Z�ai˩.'�M��,UZE�L����ڟ���ر+�T��s��� l�X)ґu��%���9D���pΤ���#d`v�A�U��̊}΢FV
�8�"Cp�^�f��4�\C-��1�h!,_�p�IBf���P�f���)jT�5�d�:����ZUp�
DਕC<�*�AY����7-h'k��;
��Gn;�I�B�m,����'�!t5!�\8K�Z�Vb�3uu��m F-�Wu�lTH
N8Ĩ����X���s��Vz%�M�%L��!�B4Y�My8��ڇ�����&j	�k�+�r��p���ֿD��_]���rB:��κ� H�ںDƦ3�����ZC�V��&E���9���fZ�8��4�������;
SN"4�ҵݑJp�)��5p��R�K��VV?�d!)$b��?:�µ]�h�.�h+29���3�D�r��a�g^s�7Q��tz�N��P�/�=H��NW%� \�hkN���"CJ)��Ќ��h+�B������{�eWV���ӴR`EY`U���ܴr��AV[{��H7G�~.�c�h��x�P��a�����7�q8�����^))HQR'�,A�tx�B��ˊ@
a��L���C(�KGor��3H�t8�M�WK.����kW������B��	�,�u2�s���h���0��V4~m�O�C��2�:N!Y�ɮwՋ�1gJ�\Qi-1[i>&�hR��a�Y��"U9�,=��ZW=@��95v*Ƅ�����J��E䋲��
�瘖ˊ:��_U��.�Z�ѵֆ����s�m�\SC���J���x�"Ru�f:8J(ǩOx���+�w)�~����=���M�p"!|�Q��zS8�w� jAZK��A��� �ۣ�UK�C�}�?]�{���m�-��^�<���H�����'g�E������u�y��oi���yw}s���&�_{H����>�x�䝗��|��E~"z�#���2����׮�sߧ��.�_�W�#�
{�:m\�#��oC��_�a{w|���%��¥�ן�ܿ�x���@ףG��Ҏ}BԊ|��!X'���מn�z���w˾�����^���:�=}rl<y}��wמ��~���/}�v��q���q�;����r��>��[vf}{�����>�yꏀy���=x����/�]����n�}o� ֝�_�Z��o��t�p���Z��s�)�� w&�k��w/�����}{��{/��x�鬹��؛��x}�ô�P�/E;�;;]o�Y����U�,}�v���s���G���
N�)�-i�]FHʦ����ϊ���N��g�c$�"�1!��rbN���΁4�(�59������ZN|�HuC�L���'�f ��?�|!:*z��O��CQdQ��bi���V�.��^�1�����40i
k Y�85�iY-��¡�*� ������gP.�?�����^�'�igD9)�����J�VΔ���9C�as��|Y�]�$�>�,���p���J�.�)���;�^�*-�g����?�է�ك�Ͼ�5��W��~'55hjf7�v�t���������?��я~�����z��OK��:�C��%��|!�6��
AT鵌��C&Z�|�O͒�Y"���ַ}�!�B^F)k��)}z��E�Nݒ=�*5Qu&��5gJ�L��D��jZ��Z|�P�V�PNQ>5�g��j�c �M�����Jp5�4�֤�s����V��מ��!��hi�!�5Tw�H!k7]I���2w:Q �BJ4�9�rLe�Q�|���,�*�?S�9����t�\���:LJn����9��E�sc����q��]����gr�L����C�i*j߼i�(���LI�8ڰ�C?l-m`��i�:M���Z4�x��I�(��g8�a��1�����D%d��pY�4�Qi�H��d���Ü�Pp�,G4qVuCi!瘨���'�a�S]Ġ�aR�L�B5BV-#�Ć\d���;�>�NT�n]n|ǅ�,"�V�G�5Ƒbo�"�P碲D�K�?�Y1��!�\�A�pT��V�_��t:�B���>s ��T.��eV"5��3e5N�z��i�Z>�n�,kd1=��裏,�?����qzsz%���ٟym���W��˒�_P��?�q� �7�U���[��୥JlE%�BZx�h,LQ>k�M�Qhp��h9�'M��$x�k�    IDAT�)�XB{��j�҈�;Cl�5҄�;��l+$Rn�8�n%�?!5C3Z�R�4&���%����&��7�N����. �c�Ik!td�ˡyj��3�f�����ɿf����#E��|�;���N���z��~8�~|֢pBD9���A��J��2Ǻ:��p�㛆7Ň���<�D�ڔ��Yq���F;ID�4�)�"�<�f!62A��b���z0�2��8l{�F-�4Y�H"���jYWx�5��B(�UQ�(S>�}�c��>�C���;V�c�M����1k��	�,(W9C:;!���ȅBLRlk�����R�������6�����O����2k7T1��zS�x:pY�[�P���1�L�D��)��@&�fJ���ѩ�p0��Z4��058!6�lH"|�5��_4�E���9�3�+7�Ȧf��ͣ��CH�	�n� G
��)���ж1Y�C� �S5 ~�����|�>�8�������4S]�r���!��<V.�Q�nS�����q�#�n��I4>Z�nCZl
8B�L�֫=#q�NjnD�gk�e`�r�Y�;:��pjC�8�B@�I�UH�&+�L9���mt�qZ��E��| DXZ�~����atQ�@�!bT�B��R3��C��։� I9�,ґ���.�!?�o`�b�҅L���_nU��cem�B���ۜ95C�c-)`VW��o	�F#��&�'U���ۨ�آ�4����4B-��Ԭ�����Nsj�Bw0S4��9��|Y�%Sk��?��ϙS�f�)T!}��MT�_S����i�h-���1�.����%��o��YZR�o%JG�/�Fq(�@[nH��ߡ��V۬���L��Bf�]8�R?5���*�O�)[{�l��:��P�s��@�[2?�@�z�^��Ւ(���I�[�c���i	����.�?�rl��t�8p��9�l|�=AVQ���>�o+~q�=�z r�S0�S��"AS��)���z�J�z|H�h%hJ7B(8	���0-]E�E��{���rp�,��"d�Պ�����O���U7�Ŋ�M��r)x����"(q�!�f�ǋ�_]�!�[ߠ�$�� ���x9>pA'�jr=��S�3�{��L>��"�۫������N��d���W͒��ͷ�Z�/���zR�i�&=�t�םg�>��A�����Ү'��T�W1��E�^�hg�'!׶��ܔ����s��ROk�u��n���������W���������x|ŭ�u��d��On�~��y$���������v}ˮ�K�n}j�BD��ݮ���s��f�٭�]Gǟ�\;��؎yZ{z����_���{8�������$�:��6��t�qgE��	|�����p����Ȟ�x���~�w�'�o>���O�Z�]�v�B������Fu�NjC��*t�5�6v��Û�BM��)AH�����l8$ܴ�*�� ��qơ��Ց�#�4�rI�9@k��U��=�r�F���r�|���v�h]��lP��B*Q�t�N��ȦBR�A&+�*�����%�J
_�,V�uC�5���M�tQC�X4
�E��مfZ?�9�A��	��_3�Q��9?\	�D
��D�:) 2��J�H3��sp�Dr�
2RD�i@�|L�aZ9H�uŊ���>o����I�m7�#��'�|�7�+�w���$��wzE=�Y7�����(�(���ܠ�8�~Wu�{:���WR)V�
A+��Y1 p�Z`��Z�'�*����r��B�"@=�X�wQS�S�����o��'������ַ�[O%Ȥۦdը�; �E����(P�u���S�B����k��8���)#4�t���rMb��/z�+��U�d1!)[�獆�����2՝^�G�EH�(\iL͐���z��(\"ߨg�5v�?��p8+Qu`)l�J��)��Z�IU�����K�3
��s˹�Zr�h��+��w��]��S�롦���l��/B��vA��fL;�]��]�t:�j!��E�vkL�:�� bR�"h9)-D��G�,���� ��I�	�V%R��Y�q���J�1 ��e@��A
��z@3��Α��Uk����,��6�/�����Uı(����]�pL��X�%4�� M�M ��A�hR:��(pZ ��&EcB�u�1��ͧ&W�=�����֢(G�#Š�0-U]xd��ķ(��pSUƧ)��Y��H:��X;��kc��/�h�u�c�iʭ�"�+��݀t�.�'��e;�nY�ܝ|�ٗx�w�u:�Yu�˧̪��.��;~G�5C9���V�����]88�B@K���p ^Hz��4�*M8�*�o:��4m�f�)���h9�Ji�ӳ-B��8ubs�˕���V�ԨÜ"Ѵm5d��O�=�FB�@#�B�� S���B�ԧ��)��:f�t��Π���|[�LS(!R�k�)�wʵ{h66˄�S�M j�Y'�cJ��nqYxQ�t�\-V
�q:�Zth�4)��J��6Y�#[4k!�V��l��Q��^����T�	�oLn)�%�K!���2���Լ��+*7�ܱ�2��*�	�UWh P&�gk f�:QnZb�HY%����15�EK�)M�-2L��V1M�U�4��b�
��F�bT�2N��@��Ȣ��S�~b�[=�6���1Kaӄ4�>�K��+�\:@m���|xH4~)��M��8�N|��v�b���E�����*����%�fN
l΀5�.�Y�>��hd
��L'�T7DM�Ɣ�NG�c�O*2��M���RD�J��ȦB���!�aH��!>A4霘�\��`��);�H|��@j�%r�Z�7���%)T�9�Z��<�+d�֧��5Ȋ�`�RQG�ܔ�ȥ�M.�����"1�F+q8�=ǁȪ�hM[#��6�����ƅ��PU���b�\K4P!C��NMHV�:|%؜��1ZZ�	뜡O�š9��6�9ƈ�  �b{��2��� ��G'�p �)�ϩ%�F�pS髛��^��8��C�=���ܚ}Y����|G:V�I�Ӑ�|���B�"����u�\ݐD���@$>B�tLEM��i��㔅�a�|us�j�|L����k�M����l���#K>�|̦%�j�!�>���pk��`B�%�������i��C*
���v	��]T�
�&�Wpۘ�����7�:�V@����oq h��3~�ȶ|��gZ"[i��-?��љ/��dqlB�5L9�ʦ�Fj��O-����ղ^6���1#+�Z�K���tj���CAM����K*�N �z��!���&M�B��}�h5�z��=��BN>� Q�rR�F ������ovh�I*��=�h�Z?�H�'����g�W�-�'����t]��爘�=�m`J�g'A>�y�>�y��3Z�����.��YƋ�j�{c��ȟ��I��+:�y�����Ҿm]�yr�i�wK��=#<=9�l�W��������ٹ���U�J�Rk$���9N}Y���H*h�n����⾱�r����}����?>�wk^�]y*ptqr���.��M_����o~s��_�\u��wON|����螟��ݽǷ��qm����O���L�����B��c�;��b�}�+�_�z���9���}��/�>���������qD�x�!��-r􁖌c�K����z=%�~��c�w�����GW��|}�����zy���N��"+�vo�o��<A�DΉ1:8�[)�6q��V�_.k�++f�@�D+��Xg��tfZ�*M�����3&���i��_�S(�4ZUL��NEE�>�nC��©a:g��ӷ	��8��~�
�@� ����|)�V+e�f�u��D�嚊�EY���7e�2"�7UE��*E�rp dR*�$��������2� �
�P���)���δ(���Dˍ?kj�Z"��F�n�"����Z�t���.yQ�}u��tK)�N"�ct�'hO0%��]׆7E�u����}&eLx������&0�H�E��g>�(A�Ԥ Y���&jh"*׊l�T[jJ����=������Dӻ�3u�������gt)A��BH&�~�����Ӗ��+��9�Du&�l�|�ʒ��%U��\HD��ΚD�|�)�iJ�4eeՕ&-�Ӻ��HI�cxr 7,�	Q
�D��z0���'$*Ī��hM�Y�i!ր�U�s�R�
UԊL	%�̯�R����Z!�9�SL��Skw��~��G��Z<&�~����m�_bs9)��qFz������,
��ַ ~�sm���m�|է1�!���r�cFgBg�����S��H'�XQ"n�:�?�JгE����tZ�z(�zm��8rk�u�T�]�r�L=d;�#Cl)"�V��팩a*J��Z)׏ZÙ
8�T�cC�TGW�Ab���SVB�
��p���dU�����TT.&Mg�g۶��#"��kq�C�#X�t�V�;5�_���Y ���a��R�c�/JS3��e9�Bʪ�(r|8��=p���|8MR
���|�]�-�fd�W������)X�s�U�|��>��󧖠(M�-ے}ZڣJ�|������JR�B���?���U��M9v�)��n�N�����sLH��h@Q�g� �QHdȜ���)�a��N!:��k��"*�)�����G�	֙���L��ɘ��t��_���g-|ӢheA(Md���Z��V��B���N��	D��&���p�L��A�C����k��T$(�����7���tD5S���~��@v^��z�֠&�����
��l���j5LD�#(ʁ�֔Ut��e�Ķ��~!>���}��ߴ�W�2����9�������rf��h��bX���ZV�D�)���]2Ec���&�Tʕho!)�$������,:)�?�-����R]�F%�F��P��H�o9|!Y��㋦fu�c�+�|���Y)fm�a�ir ƴ1N��ĉ��HՁ�X����N�9�zhE����_ݦq�D��8�qL�B�M�c��V	S~�C�-�O�T��)N)���u;�i�Gh�.1>���H5�ϔ��V(��D���u�����p)��S��J�C��p��$�''��T,4�p�Q��ΆP0b�D3��|Y�-$�����X�t8�R��;c���B�!����|G�kY���#�� ���6h�� �k�h�t��!"T�� �c�V|�d�e��$ȎN
��RL� kZu|k�f�1�:��d���'��C��Rnu!�]�T� b�R��|`�YU N�-��@+�)��PA{�:���I?��L"��1��)�V�c�3���Ul]L1'��qB�BR�����֞()d`
��F����%	1�L��<�@K�5�R�ȅ�9!� -��6�C�ͯh��BN|N�Yp��!Mp�RbNz���+��.�~�C0D!BN�78�*��^~��d����6Y4>B;�Y��)���=t*M�rfEh��������A N'��w�~Q8�Q�/�u�J�I�߈<)��:<~��D�3)S8��U�)�r�_�e!��r:�f%��y�9DLӯz�Sv�ڤS3d�D��@�t[�� h,B)�h,q����aV�_��g豈�M(G�Oh Sn���B}F��"l��'B�H9^z�-�}kQȵW�ݍG��cu�aW|}�Ǌ���8�RV�w+䣒���p=�����Su[��x<�0o}.҇O/<�ta���K}�F���-
CSQ-�+��?��?=[������'��n�FW��..�>�䷢�Wo�y����g�VG�׆�����c�g�X��ru}{��ݣ�Ͼ��~�kߺ��ߠ�9�7'���sׇF��g��<���q�������׺�Ï�N}��B�������h���c��:Xx�S�w�}�?~��W������ӫ�{�����|���Mk��'G�B,�Z��a!}t*r�.�="o���e�m��{C���<���o�]��Y�"M+�;ex�㭤?�P�Sg�N_��3 g�=8��^�<!����u����t�~�,^�t���r�j���esF$�d�6�t٢Sh�B�,2ǘM����-0$�~Uj������"�G#	,��a�(^�r�E �.��1��8��Ǩ��J	���Q�4C(̔��\Q�l��Y�������Y�*&�V������Z��3��)�V:�@|#�Cg*�2t���GM�풔4k#��&ݷ׽k��}x�[����\ޤUA��tTa��[D� �Bd{��6�w�=�i�8�"��rMOR����]V��׉t[0�K�Yu���?5Q~�l�|x�M[N�����t���X�A'��1z��yK�i��M�V��F����%c@���!�4{�F�啩0g-�
l��Mᶃ�^GSR!~����q8Ԁ�EB ~�7 �t���ʅ�F�1k�hֈY��W��(�&��,%�*�|��"XK��!�&��)����̺(�L
b�W���r�
�������q6;�8���tb����5�㴓�T��N-Y=G�U9}�ؔ���g����B���a�B�Im+�,A�l��"N}�Ȭ7S|}��C��Ho����� ��5��*�1�8�E!�\�J��6*e[���#ΑX!Y�!�8�Y���gLuE���[Q8K��e��J�L-��ŔըtY���Ia�h@��)2�|V�V)t2�Y�i4֮�4hʲc�k��8�iF?��v�9[>)#�\��V��K�NN� Y!`-���
i3�"+dQ��M�_EYĩ�P's,,�2~"z}��Pz�!b?e!�OU�X���k@Kv�%&D�� �5EӘ���k��k�lkyk�Bf�R(2��5��Om�JX ��<�B���*��|�_!����&�I�n[8�%�h[���K)�Y�Ċ�E�>�Y��h�J��UI�	�&I\:�����ي"����@0������$�G��ϟ?WbӗQ�T�\4���Z�`|dQ:F倝KR0�Ѣr�A��o��".�G��"����CF�B��!�CM?[u>A���P�JH��l=�l:M�Av��4[�[��BK��H�|
8�N���p��1[/)��6�C���:^η)�Y.�+T�>��ɏÚvP�p�NcV���88��&d��i!�8BlͰ9�R��hj[du�+d��J�{�i$�a!cBdMY}��$������R7��i�k!m`�	F r$����@��7p���i)g����Mp�R�e�oM!1�M�v���y���asD���u��<$XW�GF0e�	v�)צ	m�U�@kӀ."S�iִ�oM�#e�k ���a�1k[E��fԧ(�WjNE)��+��!�Z�rl>�ꕐˁ�ҵ�7��O����U�r�L*�D����(�ώB���¥�9)5 �����w��h�ӡ�v[V�)?����{�P`_D��B:1L���ZS��N��*D��
hD��D���"���ˊ�a!D(�mD�D��5#�Y!�,rj�d����!��)NL�:�W�#D�fʑ#i��9lӀ�ԧ)�+�ꅦS=��Y'�a�6�h��Q�1�@�����ۊ��IDV|�J!��w�VK�'}��˩G�ȦC?���^4YRK��e*�W��L�@ND�7�a��DhďI�S��ʊ�J�7�soC ҫ5L�0$�eq�!�[���VQdK�Б�Z��2����MS�l�T�H���z��A��'qH�D�a���M"Y9�7�˹�X�{SP��u%%����겆�1
�t�����vI�z�k��G(1͢��"�1]M'xE�S��LR洍�)��{4Y
�_K�4�#�WS.�Ҟ�U�T"$~�#�1�SQ.AYhQ���	&%����@`c�r�����+$��i@V��2mIܔe�Z���z�J��#���W�\���r��',�˞��Os�\�׻��׈ʹn�_��������\�o곏Vo�����4}��'�G�x�C��cT�����    IDATjzT��S���������Vv�Ú��8�����_ʹ�[)2���^��Ӌs�����Ft�<��5����+���+�/���9���i��W�q�u|���{-�qr������ɓg'`ޟzh�����N9~rv�^v~|~�j����V��� �=_]��p����ҩo�=>��׿����/�������������՟���������_��z���߻7]eށ��q���ٰ|�f��v�C������ks�`�L�_��e����b��i��c��*��`+�,)�C�/���{�����mʊ�s����E'SN��Bzпi�N'*~"YS�Q.*�;�Pc�'D\�Χ_��Hb)#XESṈȉs����P0����?K!�����9���P�(���K�e�A��)g:I'M�pZB
�PV�R0�ARf#$5��3�:��AȡY.A�R��6B��E�8�Nr�Q�@)tJ\B����qh�2�
q��pLL��lH:;��T�r��J�y;���4A�,��3�IE��^��kW.q�hB.�rW���[��+��˲!*z&��ý_��}���9�G�����,��Կr4ۥ�Ⱥp��ϦP��,�H�mBSu�\��}wHS�A4�7{}RS���k� �Z/�V�j�~ p����@�9���|U���7hB�K�԰Z6\	)!鎐�,���jes�-f-*�������i���.%<�,�i��_E֑�|�)t\�3LN%$&�j�����Vc����B���!�6�/Q��/>��L-S͠i/M���,��in@��>Hq�@L{6NӅ$��('�ͩ��9<��.��?��e����8�D�˟-M�������U�O�ژ*��&�!+N�GK8�ᘆk�O�U��a˯V�1��|-U�3m�'�7!N=�[���=K.�����FM�h��=8Y�óF�f��ʷ� �Iч�2L#S �z�Eub@&=&�!㷍�����w@��m������"�cX2�݇85Q'(d
�Η�i���0��t��hu��o���
��������
q�:m�q�c���	Q��lɝ �f�r�����ē�<�YY��0&���h��M�[S}���{@�UO4��}�_�8"?���m�OH'�R�4��Q-/l��y�Z�]�¯yr~;���)1۾IAK���H,ڴrS���z�Lӑu؆U�R!{h���C�d��6�g�d���0�#�	��h4��Hm ��Z��)4p�w��)��7��@9~�M����R����MYS�R ���+����l1�+�bګ��w�F���jr֞ܪs�1��4>�E�FQY��j�p>G4eSPc�T��8��9iV�O�5La����ODT�)�j�(p4ё��
��5�zG9B��ɯD�;��mH~Yl
�ar�Dn�'[{|�h2�&2LS�^Wï�i�V+��:1�Ǵ1=LÊM�95 ~��Y��l`"��4�>���KD�A���o�a�CAb:BhbB�J���δ��d�s�60Sf�Zb��[�(0�А#�_��'m��%��)~��~|�j[p8�2:�i�S���әU�!�4?5g;!ZN���ܭb��HGkH��B��L�L���=\M<����{
��薘�E��B�*"�&�r��ڷ���5�Kd�Y�yq��f�9"O.rH�F:ν�B8LGMY�����	���~�9�{T��1
Ȧ��j�j���D0g1+���8E�e��	�1Z]�1S��(�!���uaC�ښB
�U4���Rn�Nr���oj��Ք�Sn:�-�4G�[u	��/�<�9,�,NmT�u �Ñމ�B�|���1 N~ഁٶl��m��/jtnH���m�� 5m	|%:��Cv��Z�P])A�����қJG�fJĨ�
Q�|��J$�f�2�i�_?�+�؏���ŊV�E�K_�M8���	�5 ���m!)�K��h�*
�'�P�ot´:�(kDj	�1j[��&�%ʒ��hIV:z�C$r��q�z��&rx;fZ"BN=𕨽j����f-�4��9F{%$9���ab�t���*r �ç\.�3H�F�(fQL>kڨ=�*�/��Gc���s�S`k&��D����X��08jьɟZpH�@�Bp���;d�RH-)Yh��S+|N��/�Z���D�8�"4����b�ő�����6�>CdIoO�����G���B��a�˅��N���ï�pv{��]=i��Mo���]1�뙞�;����4�)���zz�Kc��mG�j�z���;/<�[_	{�;P�Jg�������u��������uR1_3�>P*p{橪U�ur�5��ps� ׽���Z+7w׶�׿����f�[��_�!����O�^�3�g~���=ףO���_~��{��}y��:��ƽ����{��$���.}}}s}�K[z��w(-���3OGh=o�#R,�\ٵ���~8�+�[w�����W_|��^�������_����q�wpC�c��"��ʷG�����_�9����Q�Co.���2;I���RX�2/�[�'���?��Oo 5@ʿ9Xĥ�����I��O�q���'@�!m|��@���@L�*b�r�L�z���g�D�5cj�2B8�n��_"|��JmqF$fW�\�Y��Nj�M���J�� ��Z��j�-��(��ZUn�h>�i��MY�)B-��bj�鋶բ�d9E��05�C�V1_�1��JW��0E�!�����C����b
�*�g�É�AP���CV�{�E��� F4� ^]LS4��,e�9}�\i�l'U�+='���ň&�۹n�\��:��Ht���1�*�\'� f
h���HE!�D�=�.�*�����_�����a<ׄ�[��_�>��A�W��!X��:4-�,�'�A��,<��r�'�v	�r{��O��O��m�<����=Nɴ� �Uձ)�a�Tb�"�kh��a���RW��'>��J�&+Ҏp*N�-0E0(�Yk�?3D�~�����d�_���:�R����kL�Ν����i8�Rc�����	ͺ��يR>����B�B ����[��s"������3�#�i���h�g�Ŋ4�z����ǔE� �9��WZ�:Qz|0M;��\�.��Ƿ��)��rZr�*a���UD����8�B�$:��.��i^����j�r{.2���;�|�&�	��Q KJo���x��g� X�~���\
r�nU4 A�EF���r��O�)�6����a�z�ᔎ�m+� ��ⓢ��q��t"l[��pD
F[	)�΁:�i�-��`Q)G�I)�yx��4��JW�Q3@)DЪej(��K�?��b�:�U�)�~D۷�2�TH�^T�:3{"ޡ��L���!��"z�*�EQ��?#s���*`��9^�� e-��Xۋ�@"�c@6eh~L>g��N|�J!q"�Q|����%%Z��V}�뚆�-�����~��W8��vY�a!|��$�iE-3�*B�!*�'2D����2v�G�����B8I�kÞ�w����lMr*:L5Y�BR������@mtL�)��/T|���������)��?��?Ғ	UEjD��[`k�R	+���[;�N���hK�B�02m�0���B$K�����UZ.��e!sd�(���r���Af�e�FՅ� �7e�Дl����=�Livߨ��ϖ��Q4��(��S>M���c���8X⑥7� �C*m�O�o�*���Rز��U�ɓH|~�t����҄����uo=�\Ŷ�벪���$��l6�
��/�;o ��?����t����]�:����p�>'dM�1bD̙���2{�%%ZE�P��W�
A0�/Q
Y�ҍ��7Ō\Q��,c���,q����*��1&5�h�-\
Z�!��h|gK>�G�l*�G�S�'Ü&+����C��p�ފ�E�r�#��9��3MJ�������Q'�,*��AH�À�	v�+M����A͑�Zʕ�G��g�	V��ٱ��'������R�re=�]��o���G�X��IX��7x�ȃ�r��?��Z�'�О !�L9�q��b�^�$�E[H��|!V]N�"� �Y݉F0� �ԤB�i�9lr�R3�r��*�t�A��7Mc�÷��p���9�V�_�%H�� %�ρs��5�T���8��U���Qb)dMmi�8�!E��3Ym>��Y3����FHd��a�d�&E@�"(��+:>'��B*.��( ����~��~��s���L4�f�|L�B|6:��Xi��X�yQx�cl	�j	i�V� �?'N��S�� ��B�L
����QH��rʊ�ld~��$�ϏVJ�3ӔO?`:�I��Q!:�0%8��L�~�T�; #�A��M[r�:O���3��tc�]���L4�:@���W��C)��O�����T�����ە������K�,�M-g%l{��~������j5Z��XYK�����<eR,��w��%X�S{�YH4�����Dh�K�*�`p~��s�K!ȩfU ҅�"2S;���kd�ℤ�V:R��А9sr$��.�c�h�(KTLT
d����m=�3��p�c}s���W����~gXO?�ί���o+\��V����֓�����]���K_A�X�4����zt�1�O�=���wn�y���D����U�_����6�co�;�:�v�_|�����O��g�j��oOU������Ź�ښ�	:]˹v�y�xws�ו��띗w���.�z8�~�����>��������[����<�����z�w{r��|q���z��?{���Ƨ^�y����<����Mo]or]'��Kz��η�;o��租}��ח>n���AAvsF��B�>��ԝ�t�/��m����~Cv[����ґ"�ݙ/�{����e��4��Ա^_f�>C��r���:m���EF����<Y��.,�[Kیh�ة�xz9�����-��\ R�p����jx��xę�Vt�j��n= ����i8�1��u"+'e�)�I~��J<��l{�,>NL)�|֒g���G�T��
mI�Eq�L?�C'BY�
�4�J1)!�ȯs>N�ٖ�8��f�G�̗�)���m����)~)���U��2̌8#�����op�ˑ(dZc�hG�"�x�I-Rc1��L��:�B5��<q��+���p�{���S���
J�(�Y
�z$�}n��9�JȪ[�)�_`�
���K.Ŕ<����g����d�MHE�'>5C����
q��ี�u�A4e�����P���EIꖦ�4�cf��;��Uј��!P�u8���/d��J�~�ӟ��%����a2�J�BCB�]U1�4�Z��Y�F8��$���5�/j�R��i��j�q*Z�B�5P(�A�㣙N�� � ������0�������D)�Dc��h��h�1����S{�p&��@d�Y�۞H/'X��i=����t�^�DK�)��gjC�ߞx��}`F?S=isVy�恁S�z��X�;1�'��?�ث�[��}�]O��l+,�y��3���ꪟp��B�eY��:LG�!�C��Y��ʂp����8~�s4/��g�Bm�Z�8p��+gBLq����t�@fZS!���eY/[TQ3�5)��u劓~��4I���ȦJ(�_�d�����DfZ���$'eL��p��p"��YK���:7����(�3�Q"�r���o����8�B�����C�a�[ى�M�E6��s��2e#�r(�W�ne��4L� ��/�2&Ъ{��-��tk-^evO�\f]���	�-��O>�ĩ�Mu���?+��s���S:}�V���?/x���I����#��)W�q�te-9ƖV'��\�Z����9���=��p��g#8%���n�ǣ���I)VQ�,�+�+S{�er�*�r�Z�p���h84
�]�0�<媕�lN:�L��-)� �$K� r��[�i:�խ���\�\#)��	�,ܹ��_���D!���հ)��t����3�v�٥����Z�t�'1ŧ�Ъi�Fd!���L��-�h�τ� ��J�"fN�p�Mc��d9,e)B�ɩVRe*��d%�/
�^{����Z�k�n��L
)��5ak��2�Vd��^'��9d-�f*��6YBU���p������q�#5�aԌ�]�9
U1�H�hڨٚA��q�)7n��s����M�8�7�uV'�/EKx+��,�BF鳐t��gE��r�K�����|BZ;�~���0<����^]�d�
ɕ�od!I�&bZ'E���f��r�`;j����*�h��b�X׫R0!FY�a�R�ѤDc'�,�h8�L��@���A��U�V�3�3��t�0�5l������^)}R3E�#pjL4�����p|E�M;K����4SYɶ���B"p N
M��rF�p����	�G|ӥ�s0kHgV�����DJ�`�9��*�4��#ās���:dt�ΜK|�M+�1�X{���PY�q�j�}��Ǵ�Ȫ���`�1����������i*��tD�a$�N4~�\>r�J��pV��Ay�@��π3�� ��<�ҥ�xd�im�w������s��h�8F�%�U�B�^�՚��?	��ud�Ќs�	MY] ��Z��4�◅�w���m��oO�Ve��7RP�%V�PG��p��h�'>�������,g�� ��B	�b��>?�:�&��[cˑ�������:�)�fL�F&%G�o$R��1+aL��7dY�D�ņKg|�L�B��Z����7b�1�HdRD��_�~u�_TW�dS�u8�����1��τٖ8�����zcd!Wz�dmÓ-}�l���dC���� �V�&DjZ�+��eտ��R�N�p���@��/��S9���
��)Z]	EcJYBO7�8h�c�1�+)z�<���B�V{pS)Ee!�����p�M��?W_��	����@l]|����,K�ާ��~�]����U]⚾��$x�+O�O=8� ѓ?�a<.��I�sb{�]���Еk���ĳ=�{v��ܙk��n�4�G�z����?M��g�mH�p�pG��p��cXd�\�W_�_�_{)��������S=pe&�~��񱞏��#�e����~�_��p������A���_��>?���羍��4���[Ϯ����c��r�~}��o����ˇ[�j��0�R=�\_q�lN��=����S䣻�/���������=�ImCw'܌rOƭ��сӪ���r��t��#��ޑiC�s����R�t��n��:ܗ�W��OO7�s��Prߩ�?gM}"ES���@�pc�78)Pc���Eni�!rG�W>Ј�:^R��D�ҟ)C��8B
M7��/WJ4�*�s�"h���/%?�*�3��;�)!Ԍ84��@��sZ2¾�I��~��4>_38!F$���3���s��7"ԃP),��*ad�5ũ��D-�#�hC�5b�b�&BH�pLSXU��B^�F)L�Z�!�u�b�G�$˯��@�F�+��r��2jC�4�z9�k��X��8]�{ͺz����ܺ�mF
��rL-A��h���+A�G�\���]~���{��͚���^RR�Scɒb|�u��\ۧ���mf~�||>��H�v8<{�R˄��-D�@Y���o%z2��^����ɗiynss��[��T�l��k����h�~!0�)SOǦv�M�Q]S8���jډ�#=M��2|~��h�E�n:�L�p�***޺�<6�\?`�[Z�Zݧ�q(p�&��&.k��V!:/*��(}$�U���l�B�ȅ�1�!9�t*�( �RƢ�
�Z�g�}��S���S/'I�:%j�E9�lܣP8��u8��c���uL��nu�37�I:8D���Pd/i`���-f�s���Z�%���!��ɽ���K%"8�(eq�������XB�`��:�̈ ˭[�>��g�B�݈`TŮ��� *e�>��K�T.f�S	�U�J;�`���br�����y��l�#�%QK�-�XbK�S:�����V�p�~��    IDAT��5ʪC�h1%B�h�
�9�v�*�9����k�����}�:�8���|���XZE��;�R���B)�")>5!-�EP].�4���e3}�t�C��z1���9:�,e��r;p�x�ۇ���-߈O�9�U�]��i#�^�	�A����5�9j�}���p�]��v���M1�&1��i)qLm����҇k&N�$�c� �I/�Ȭז��'V�a�~�I���'b�.�P"�g
�5m��7��k��t�L�r%���ph�e�1R��1m-Fի(��E�b	�'e��"X�)�`LgN���!B!�`:��h������/~kqV8c	V׈��rR�I�����܎�UH�`J\�mPu�:���1�*B���dS~�����Rb��	M������=�l�-�`��Y)l��N�z3b�T�D��^4~�p�ӏ	d!�|RƘ�� ��m8_��N:N>GȈS{՚)e{�YQ�Q�1��q�KDG'���8�n�ϊL�E[_i#�B4��pX����c+ǯ��G���c���[/Ģ�R�������Z�ʍ �����4M��Ed�8��;ᅪ�<�砉֞�6F!pU���CQ~馢�����	����E�KX�6��8-�����(E	�旎�I�(g�·R���DV{�!�zE�UAV�qHq�tš���>��隔����e��v.�cT}:�h+�<}�d%���2)9�J��Rn��W�Ҙ��>�է�S�Z:��Om������SR��[��ಊ����PuSH�O�N 8�$�x�r�4B��hD�h�1=�����s	M�-s��3ky���P-YpL4��ƴ�,�M��B!�n%tI�c:='M�D�i!���3&%B!��	B�C0m�W"���1��t8�L�8B�"��u%���|cݶۢ���*�)�V4g�h8ᭂ#�g��>|��D�ʏBY������t���\�q��CYn��=M�TA�ӑ"ݘ2G�	ŏ0%�l`��AH-� @2
�v��o�؏eI� 7-ª6?�]�h=����L-e�h#�Z��v'g|Y�<��mN:1��"��@�i��p����g�!r!hr�`�P�&4����T"G^/]+��5����K�����4e�Y�m��e�	'����ÑR?��Y��!���+�\Y�pD[H����@�b	D����oQe�3Yn��h���OA�h���1"RpL�]N�M�X	�F&�� W%ex ��
�����JHˤ)T��E۫y�" U���z�̉�gh9�)A�yǤ�g=�tWu�j��b�������՛'>��������f=�K���3x�v⸝;+n/�=N�9�ɭ�'�G�����^����������;,�}����Ց�n��Y���~��{���9�2����$Q���縮�ߞ:�y�#:�<,�E�k�>���ԉ��j-��~Z�vV��	:������.<g�Ƴ�V�0�=�jOkO��]�����3w:���ϟ]�]�x���q^�.�nח�X����ݵ��ǷǷ�Ot�r����|=�=?�_�}�N_�ax+���ţ�___y��/֭E�tV��ڳ�h܁���3Yc�׳������2�Z�v��� �[��C���XX%qo��o�O�#�-P�*�ҏܔU�@�s�3�_`e�a�_]�H���41� j�:c+?�9�M1+gĔ�At�8l�O*Y!:1�����l���e� S��+��C��UϢ�G
�.�L��3c�D�(e�Q��m�*�8dt
�Y�t�)4E@�U#BǴULp��!��V�T(���>#[J�I�ψ��%�5�tFNmӑB¯�D�LC����?8�؛/��BZ�o$ކ�Ӕ^M�DH+�����S�~^0/�
��3%�ی@M���+�m^Y~@@��)t����z�+�~S��r���).��SF�V�U�l4U���j)��B%v4!��uG�̀ZB�$.w�ncv[Y��}�]"��J���	���=x��[��\[���{�i�FP�f*B��tw��怢j�A����Ec86A����89pN�������Y
� �TT�����	Z����T	������6��F�a)D3R���c��&�4_5�.IӀ�B�G0�R^z�����V�^]Q��ˊV��4g�3�t:� ���s���6���9<w�%��]ꡊ������o�3O�����Oܔ~+uF	A����B���*��#��GVBB��q�V�r+�i@觻������,��j�I��O6`���U�)�o3EM%��T�	�i�C.˴������'d��D�C�6"xE��KDs��0����KQ:)Z�*�Tn�d��y��v^.kiB�R�ԕ�ȧ �Q��Dh"��8|t�Z1M8C��ȡC�%�9�BjF:��
F�.�O_�����D��f,�D����pH��`~m�sp��`	-�s#5����ۿ�կ\���X��z`~�xx�y��k=�R�]�\�4C��O|!�ӭf+2�kFc-���;H[�#ď`����3��C�A�H�����L�P#��H�`r��5�	J�s��h9�)p�5��e������Bƚ�3�G���Օ��������4��Y-�Ñ`��!h ��AӤMu�#���8�� Q��.��ǗHW]�$d��rD���?I��+�B���h���<M!#ZWf`��i&D0�X�� �%+QVc�;"����(]�r�dk#͊�h)��Vb�h!j��קi�>�hN�^2����|#�9�ٺx<C M[ˬBn���M�,{e�D)8|
�Z/DK|gTiD�"�%�4�*8����K�qF�T�N����O�� 1���NF�TT"ߊbrdMS"�a�6��/Z��B�nI�5������L�E!�8�Z���X⧆÷���HM]�6
)W�:�E�6
��$���I4QS��k��\�P�$b��ͤ���7�4��o�5T!2�z6F����,>~��>�O�p�v��I�t!])�ֹ�r�u+����Z|�1%��J	�\����F�t#?��I4U�T��l� ��!�@L�Y?�'*�M0j�4MN%F!�����,��@| ���~sP������-�s��9@RZZ�� 3u��7"�����Ϣ�"k�M9�rpX��qD�@�I����rX���MC� �፦ٔ�C�iu�M�s�Zrd�\
���tw�z�*��% H�f���S-��FS&��ȁo���t��2��H΀r�包w�$�s��r��d�R:4��Pu�u���[��GV:�)������~b"�*r *���9��J���Bp�����%��DFc�X���˪�*�p�JȚfȦ,��G ����S�82��5 }L�&���k�tY���.�����j�!��V�8�#R58�1eξ4ͦ��l�����U(��ԂD+Z3	�'&N���WG4!�g�
!̕�>l�5������Ia��CR�D�0�Dj8Ur��C6�8�m�(D��#0BE�M48���XmT����.D��!|���X�KB�egQ{e�@��0�Q�������8���B�S��縪(g�B0��b��P���U�Ҁr���w�D
�����M� ��ܚ�/K�h��M!|��F��@!����T��X�{,�7CzD�n�=?>��"�o�\ʇ����7�w�w>s�Wi�z$�=�[_~y�}�ގy|vr����i�}@ۋ���g�^�����m��n$�0Zo�<�΢Ë��o}텺���?����up|�>������ĻG�%T���X�:H>�VkZ�w��i��|U,�3�E~�}vx��C����qs���ڇ��%�h���oz��w���|���X������y_鑧��'�z/�_$�ع8�يs���
��x�����5�é��:X�|8�����s��E9�������9I�p�M2��ǔg�l�P��s@�M���pL�X��Ł��`�R��4�����3�Z@ˬ\w�,q�s�`���!��� ����1��@jɔπ��R�9%��� ���
Lm~�٨�U"<��'8̚�;��f| Ub��ԃQ
�z��.JMJd�i�tB���1%v���&Д�c����ՂLK�Ԝ0@�,|>�)#�&���Rn��3�z�$>��HDS�E��b��`��BX˩ɢu"1�@̈́�r*!J�/KuN�F����\/Fgs�@��)H��߅�!w}����t�XV�$JA36�s$z��r�º_J�#�4�uQ �a	���ǐZN���"����rbR�('���`�M��Z�ܟ��o����UG��x��~֥D��?�9�ikbU��3Zn���^�����fj�Z4�R�� 0�q��L�hF�i~N��#:5�X�ȭ\� L��RPB�DE��j!��c�vͶ�Cp��2M�iR�!ΔTBo�ȅY�:��>%���L<��4a2~Ӥ���$r�ʩ�8r9�2��pW�HA�ѩ�á�C��l|O�-D�[<Me�1V��Vc���5>�H���hu(��d)�E�'^
2��#��*�|� +�H�V�%���Mq��,!�H�	��%r�����Y|��#��|)B���F���� ���R���N�rT�SuQ+�2�/$�/�EqT�%��p0���,�\����1�N��@�[;��>�L��fd�k���*#S�J�.A]��Y�(��w�[�P�
�9^�NZ)���Ň�e�a!&��F̤¥�Q�Z���Ș|��E�IT�H�����C�:�<�d@!�����QT7Ռ(��=U�b��l�N��y�J�Z��Č/�]�����Ü�^���9�&�"�L��	��F_�bd��*�1q��G�Z���4�>�o�Q�N%�ʍ���E1E�z�K����v�6�0�P�3�0�zN0����Wev��\SKsM2�Z҆i"��Bp ������ �L ��E�o!*z�0��DH�ȕn��C4������(���I�4�hH��s��f;B�d�)�*��?S���H���tji_3�4�>�L�E�CPt�������@�($H���	7Z�B��J�� d�;ͨ(��ǝ�<�I9f,Q�V'��H��%���0듏6�\xH}vȒ����o�T��Mz��jY�=�HS��H���~D�#d��^��-㫋���P��8�W1m-h�/�*ࢵ*J-<�il�h�'ǈodр��������de4m�d��a�r7�l��	7�Ň$U3�B��/ڒ������W"e#d�1�n�PS��22��\~�y<@�E��u�\�l:xY��BR3
A��,��-Ec�-��d#&�BM!���L��K��@S�pf ��Lxu�"���(\�f�� N�}�\ۥ� ��U?��7>Y�!�F+��Pd�t�T�C��pf܀�Bm�~	��R"��c���TB
C�*�L�L�[,_�ɵ~�)pJ�T:h��)��j8Әr����Jl�*�W�O�k8YF)U�_!�ٷ����p
�ڐ¤��9�m5N[�l����Z��h�i��DY���}-Y�D8�(�����i*T��p�qQu9�B�Z�YEM�E�:ϯ_�ѴB|&�#�P�Ԅ�P��eq*'�O?�h�Z*
����a�Հ)Ǳ�k�쬨Z[��.�?#|�	��j�с�]@
���"���| ks���l�1���}��˅��)��r�8�<�:�T� 4�t&���U�h�Mk#�f u��ZD�D�'ܔ��)�!�qЈ������vS:�*'���	a�XS�hjdd��l���pj��p�8t���&_HJR1!��l��V��cjD�gE��c������k�%a��>L�L��ԭ+#�5M�ض�q� ���֘��8��&�Z�k�q�^�B��$T'q��`DB��U�%C�g�O7]]��F��k)�Zqt�������ӳ�W�W.�g">x�gy��z�y�1=�\�*y���HO�|F�ɽ��a�3��/�����M"7޻�z�'Md}GǞ���N��Z?m<,��zs~,�`כ;��~���|;��:�:Q��dK[��'���������&���s�	�5W5_�����/���������_�~u����u��kwpn�.}���{�s�����Q��a�n�}���u��O˽=�ko������>�V۾;t�F��LQo��6�h1�i�?�9\K�^�É������������u���QRĥ(Z�t!�::�=1]�V�HJq#B
�1d&DӒ�o�U`
�uD')��F�*W(���Ub��_�Y����ɂH�U�M����h�"T��_��t��㴊@")�N�6A{R�F#fE�N�����Gc��*4�I>�����6��LK1�[�l?k �i������g+$
��C��X�V����c�0�UQ�P�Bda��id��"k@HȏYDJ�)4���OMű�s �*W!�~�G��\��dMsb����T-�F�@NӲ���F�E-��fOp��#�B���.�9�*J�JYVar�p\jڐ���
�096�O^���M;���[�ƥ�]��.�ބ��G�Q��\�7-�7v�o���n����(&S1�2+QL7F>ǆrZ �b:�C�LE!]��D9B�5#�͏3[DC0����"(��V�Yj8۰��e��3��( �n��`-҅0�"dQRh֛�XWh�p*g�%�Ȅ�j��3|B��\��q6�5�HM����oQN���-ʞ�,���8��w�;Łn����?��Oދ���N���>h|:vO3%rR&��r璊Nek�V�� �šD�X�V��9p�B4�LH��p��ZY���D!V'F`H���,�#$Q9Q���S�1:�t�p,�_�tjh��w�����h�`�ٔ,�t�t�jY���7
1���(���g��-'��hJ�X�
��REV!c��D�=:p
�q��p#p̔Y)���K5R6ZBB�3U+f���^A�7���*> 5���n�����/սX��(��P�b�J{�Q]�)��>���?��8}�35��������'?��ך���hֿ�C���C��k/@�(�M�#S��Jatځz��R&�c��ᇛr�j�ӫ#��%0�h���EuD(T�:��gAf��*�3�.Y=�u��pK��Q��~M����	?S�h4[]�1��i��0�jY�����������<�S�����zKt�(��Ux��s#�Ȫ�Bq%��:��u�¡��\E��%���a��"H+�H�#�a9�U�I�r�)|˜\�U���g�6�5�#�>����q��9,0A�:q8pu����0��.��2�hSc�)D�����7�3S�M rZW��4�>ј)q~�e"Ԅ�E�9��_�O��J1吚�T.�S4_�h3���tX F�J4Bf{˂0>��N!��F�z(J�>�E���B�&��dD*|����7�<��N��Y?�p������3����\f
�(�t(T��Z{hJA
�SY��L���4���r�P�4R�r�M9I5*'>����ub�4�\�Fӽ���@Rt$�Ǐ���!L��q**%�q����Q�&�xd'9�6a��'�X~
S�u!�ۘ\)��׃Z�Bc�����4�*FS�Ƣ@K�4�������3�(�$�.�i ��:5���T��Q�+��Z�Ӈm@��qN��)�6�щD�rh�M�񒞂,G�� j���dM��Z�h���l���jC #N��(p��3ki`~�[�L\u�m�~��8�]MI�1R�����X?5дQJ���PӲL��h�%�`dG���Rc!Y�*!�ҵm��h���l?�M98�&Sb/s��+�Q��O�ΐ]������~J08G fj�!�CƱ. �PN!4�D��T�Lq��f��M�:)�)�E�/})n��B��/�e|�u����O����E�`�R4}��r1��8e��R�r�r���t�Zj2���#˝)��d�x"�%>������*�e�/�<A��Z���+R�Y��M�ҍ��9�DC��I\
)�r9��lx��1`��~Ѻ��>�E32Rh���{Y)]�)�_U5fd�@#�i?%�ǩ�DMV��?�!�h���{eY�7U*��V) L��ѢX�pq�a    IDATb��
�~��lB���p��&5 �ĩU��98����e��x<g˵oanڭ/��.Ho{<9��˳g�^�����������>����ZO6��cRC'�.�n����M�rIo��������[_����8;:�ߟ�NJ������>���t=�t�'��-TC
��Y�L<A\4�V�j�|0���՝G�~{�C��[;�~��rг��|}}s�����n:.އ�w�o|?�'�'g���g�����-���7��wys��*z����+;I{���8�s��y�y�����������^��3c����"�-�=��u���Qs�<���� 4�Q'�%���g	��Sdơ�tr��ϑ��q[�:����I�h^��#t�̔`gf�*�C����/Ѩ��Ѥ��crF��������^t���A3fpF��Ud�<�H��J����8B厦i
��<͗"���r#��&n{ESk��2E9�m�>;��̙��+�D:���Jvu��R��N��R�K�(T��td�BȾQ)�BMbN	��y��܂k(�&��8����eE���1�)KG
-q��D��!���H�(��
l �i!c-�d���v�3�����o�儐U4�*@���56�������jb�R��]<L�F�>5>P4������_�%�S_.�̗�#��o��V�g��J�Lu�hsyd�{���'�Ȃ���v7-}���_���%v�ML1���B~}��Z��$2>G�F�R:�Ԁ�xY�|��@�0Mc �C��ȚZ[�hԀ �5� �D�@K�����L��ua��f:���p|4�l!1���B{�������i�Ȥ��-�t� ��1AT���LeA2��A����g��6�t�oÝ�-���{�����n���RW	��F��ߡ�aG�����5IP����b�K�"�NkD5�Zb�r��p
Y�B��9��:��c��"B:h��c���[�~*d�O<5}~��2Hm��n�"h@]Q�>Y��@�z�3L�4�`���4����Ñ����e�*Zu`{�aRR3�	ks�b�F���n����L�g3���������d�E�5��}��TM:'}����*og������R��L��%��B6�д�b�j�uH\�, G	)��ő�9��|���%c"���5@��O?�-@�����ɯO�=ރW��{�@�X�Q����fJ�B88����tK�3��R��-��0�*V"f`ǫ��UeF���c:v� �(�?���?��TQ�p����/�#k�&Heh5�l><ľ���"�̧߁F��rY���Mq��^��+Q���:�jh]�A�o/�be?�=����)�R	)-$�v�����������	)^���ק\4 #�ӈ_9�Z���PH:&�)D�����(��֡�fӴh
�'7&�L��}.��!�i*1qR5P��!5OV�Z�$��m�-�)����Ј�_uȄ�l��O��ՃD!��6RC���XP^�O<NEM�ZW"ƙ�l�k8�.d���iZndx�m���X����4�a~�J\�s�ҋ6N!��>��3hL'��rB���:W���N[&M��@h��4EhL3�|Eg���,S�l�KDc5�\��8���6�S�\S=�vV�U�M�h�!n�au��t���c*�e�_Nڷ�r��"��FG�g��5%8��s�hF�č\��hF���f�v)��)�)'��(>Τ�n�@���n��r�.=�i '�S�˪a�t�5�d��6��	1�ܲ �q\	H�
4�^]�p�7d
���I12��B�K:��*⓪Dd�Q�b�|�����t�1�q�_(A�>��Ĕف����Hm��vU�"�/$�N�|�8�ݎ_W�ԛΤW�5�_��4!�<H)���+�d���^u��j�ֶ�:I�P㦽h"�)��y�B-����?_"�>#�jc+m7��٩Xzʢ�#q5G���Y��Q��SK�ɂH��4�ȁqR.��HLf"�1)H�"l��'rHU���,��t�jx4���ֱ���iM��M��5);U�*�f����H�B\-��r��Zr�|6���E����D�����qX�,�jAj�?�,�D)�rLeqZ�\�V��|)5���Xo�ҬI4���,=�*eq�l�ZEHhCTo�������RW�Z��1�\�_4���߯D�e�+�H!QN�V-���-$_bLN���p��Ϙ������2K6&�Ŏ���$�a*� I�ڄ�8��:SdӶ���qp�)'�x�y�v��ur}�%�ǭ:�ވxx���������a�8}�샣��v��X���͇��x~���ñ�%�����ͭO���͘�K�oc�}��Ս'�b:�xly~�����[yw�s��-d�Or5��=�h�n_&-�+�ST�N��n�3P���v�Y�]X�sws�����7��m_�y���*�?�Ԇ����o~�w��n����籇�������>9���QO0])nO|b��o
u=�����ʧ Q<9wwɣU����p����,�������Ŝ��� 0@Ͽ���x!����ہ�����Y��v��y� jRΙ��Z�,L!&�)YU�8�zC�;8��s$2S>f�_0��I�:>�|�LQY���/
A0�q�`!�r�U�(Q"��rY��J�(m�B!K�~V�K���Pԝ�:Y�	�9�,#&��FS���qG�˥0�Jl9�S�7E����9�����R��r�'��d�Ʊ��P�:���{�Z�sRp�wdIo��)Cp�o8�ҵѪ�RQ`:p���!�Y
�B���r�@X�����hʭ�#�P7�%�����D!dQ��ojdM�
�QEi�q���)pDe��q�qO������Q��8�Xoi�ʍc�7�c��ǧ\c|�J�/D_�.t�p��T]����%�<��Vm�����)���g����O�t#޻8QeZ�4�p�vn���:6*ƀ��,�� >'�D�W|�(���Q
0G�h�Z�K�P(A�qD�|!�+y3��eI�k�+��qBO�l��
<~'�\�ְ� �� ���W���x ����+0��6��'��A 1��Y��b���[&�h�����#�|�1s�T�ӑ��{�㬰�t�7{��c~��g�}朣��DQ®"3כE1U��0Ѵ*Q�-
��D{RZ&�Br�!>f>>�`�S�#CڨR��7R�i`��y����/Z{��)�4EE+��R"%��B:R�j	����_	L�(�ٖ�hCE#Z&:��B�I�I)���÷""�V!##h���|f:�tf�@���Z�'ᰚ�ns$�J"��(!��P:�kz���� �M!�h-?}�V�U��f���Z8
9cUg�8���l^�eQ5
	"���SN��*�2�*L����-��L�rr��٫��)*d��^t^�o�����]E�3s��\J'5�j�X���Fi�暈&kAŢ@)}ʭ%N�VS"�c�H� C�&�o,Y?m{|x��1��t��9��L9S�@j�#�o�9v�8�!�`eR:1�zE��č�\c1!1��)�C�~����7�V3�l�#�P+�)��s�ORB�O��N	?��IIĜ~j	-��$>ˬ C+�#$��ۊzЧ���1����7¥ S�3�}
?qc�Y)&j�ȝ&��4+!�Iʘ�fY�&�,��O���&���Ԫi-q�̩GT?���>�!�i/q�QRz63f�Y�F`H�1�p�I�i�6�OQ���^o��4`)!}c[T�BF���iL'ؼ�1gWE1;s��M��+rV3	B�I�t�<�qؓ�:��,<_�t�SK��8)[ER3
�-�Ve�}Q"B�A�D%���=�7��������kZ�����)+ru�5[ME��7b���"TBW�K���)�D$AL�i��̆�aj�)ė�Af�+���,��p�Υ��Ĕ7��R�:�M��G��6U�G|�fN~cE7��З�&�
�L��Zf]�V�ܡ�**�������:`��k�8�^�i&�U����B,�O�^&�}�j�%"p��� �ȃ�Y%�������e��� ����ڜ�Kz�oKu��p��|"�@9�fZ�\�L+�!m0����^(5�i͏B�jY��K,+��D/%�������|��z6�'�
5 ��Ʀ�xY��x���%5#B`���V"���sҬ�ҍm��ֹ��~��0����q
�;Fa
�D�'�)�Ԍ�6��|`ˑ�l<5S~��Fy���[Wm��
���U�Fg�+�V��^hZn�aR��8�����[Ԓ�,��S���\�9��-��P��-�Ȁ�1r��8FH�#,-~j|8k�M�gv/�Ԑg�|`��@�H65�o��vd�$�U���į��r�%UL��a~y��I��Mn���u�1��Dkg B�̩U�r�B4�j
��vTzj��To�L�-�8U�GH�B��a�B]YE�esʲ���45�
�n� ��I��GD4<Nx��,z��j4Q���V�={vq89{~�����^ܾ��hݗ:���g�����~��ձ>9ֶ��W_9�a�zG�:ϟ}���?>������[OJ=]O+�^��"L��κ�+����v�������$y�Iz_�﫴Dh[���ǟ���k��l��S�ux�y�����É���}������=���?//_������9o�SI��������G>�D��������*�jz}������2Mo�Ѳz\�Y۷^�gW������䙷������>��w��x=���Լ���RvK����B�����)��8a:'W��Adu��������M��0u!;m�7�e^4�#H�*�-]]ב��gQ�}��p�ۀ��4U�O'��@8}#�ڮ'�)譖ځ�S�ӌN-0_�%F�_��F)��������R��7�ۙڋ`���ԛ�,�(��;U ��N���-6�8��ld�z���]�@H��bW�ȩ��jJ��h��ǀLV�,�/��~D9B�B"e��3Z)D+��S4� �EK�[:��hD.טS'S45LH!����a����>״6�$1M�k�N�@��9@Ȝi���ر��lJ��CDW�B�L�(���'}�Ը5�삃ߋ��29.D�Z��q�?u�d�b�1��qX����1�*�Bg��"��(]�\9�Z޻�g�gҺ~v����e@�2�<�m��I����8݋�3Y-RgLgF�LCRl����I�t�q�Ԍp}'%_9�|K�	GS>���Єp
�!��a�!(������;︫k��㗂#���tK����,P�&�c� �[��v��:MN�����?^Y�4�bRc�����H!x���r�;�<>qr1�P���@Џa�����rhz1�*U��L	䬓x�
�o	���~G�><��`ʪwj��:U�F_.C���	�ُ���GCh��1��� L!'�r!�YpS�lu���Ո`
7�s�����釃�B�U�r݊������_���Ƒ�&���
qZ�tE��TN:NH�|U�B!-_i�(7"�u�aUG� >Bp����[��ѡ�i�*��8��
����'�&�̵��; wt0����d"@j�6*}8G?��DS"p4�������7��*�T	���yg�,�����z��R� Y^}�֌ߏe	y��_�b��!��
����2Lj �1M�rL�^��V�#�����9��*}
�3mLa���1#�5��_�l߹aɦ��2���qp�����ѹt:9F���)@��I�k��n׀��z�1�hi
UHh�����{&?!��S!)�<bD6ڙ�m�T�i�UԈ��Zg2&��CS!���,�K���|�3�S�Z�g�f�9@ͨ�Ƒh,��ZuS�T�󤽤"p�|ƩҬO
��6E��Az��ȩ
�8������/��5���ύ��H�r����l�,j����Lq#��p�2!~Sc'F��9�:U,M�Z5/T-`���N�0�8MS��0}U&ć��;��%Fƙi~���x����@Y)Ԫ�Vj-*A�! K��R�s�����f"$غ��k�`=�-�?�SK����d�Mˢ�>���k�+R�DRCi�C��Y�q�TQ�����Z�q��*Ϊ�vM��.q��B�U���*8锈������U�lSc��cl9�ĩn�J��M-x)��S�j�c�b�4vb���n�r�4.E'��K���uN}��!FS�qLe��7J$������ڐb�KT��Q��zP�Q�#g|LY�(Dc� ��J5րQh��A	H�𫫖%H��ӧ��i ���o��F�e��BZ�h�#ėՊ�����A�4��O�Z��Zz�4�,�!+:>kQ���3���0�g7*7SH=o��8���J�ڋVb��,��d1�at0k 0N
�I��@JW�d`U(���ԏ1"��Z�=Ha�؄8lJ;��MI�War����F�	��Zٶ:BR���E�m��N��OS�B�i:�C�h~��X��?u.�,q��P��+-eR�*�>���#�U�15eSx���T�mTG����id�i~�\S���'�%>8
��R��m,��[{"�`NŲ����g�mR0��os�ȵݾ��B}��,]nH% �R:�*k�(q���B�(K1�v��'��8)H�W�SQg#��@~�� _4�����
�iK3�tL#�_���*M�+Q҅WE�u��c�z�p�񍕐X9��t�rj~{��!�;9^�\��jٖK���z ��T<}~rv���7f��O�z��W7ח�|����)�[Y�u�NN/N=��<���Ƈo]�>��������WW�_}q|�sc|����<�m��m��m����W��n����t=5���������Ϧ]߬�*{�j7t���@EU�.�m������Է\����/<�us��z{{}�;m,�����忿���|��? �����^u�j�|���j��9uvt�G���Zg��&��Oo���ώ}&�����w�[��:�W�{�P���Z����j���џ�NQG�T������H|���c�^T(Y�,�v��R�v��(F�Fp�s� ��G۸�����5҇0JM9
Q��81q�֢���9�D�YE�� ������9�56�%6寎��G�i���qc��P3�cr��E�I9�^�)D�bw�dVh��8L�P�"�s*Zz�I��ӥ�S�-*��0��E��4��������$��0N�Zb;���\cG-���`Ά��_��jM'���B��6s:��R!�DR+2;P3��	Q�g�յQ@R��9[�Q's>����-��"v�Ef�N?�U��S{ԴW�L[K�vU���}2a��Q��h�,
B�T����qj����V���6N�DԞ%�R&��|�_�p}���=o2��l�W7ev�G?��uq�gm��s��`w���v���i�1���6�j�ô�-���#�1���n�ւ�_v�J�4N�
��2JGS�m�J��
��B�>t����f��C�	��K��TH�u�lp���eL--��z��gp�F���q����$2�pL6�B8e�탟�����p��G!���s���+S�3��%[���_8B/�NS��Ԭ��'��3���j5H;'�
I"7UH:�8r=p��gQ`�|
Rʒ�&)��rk�1�N'ZxKRTX�u�
��B��'Ȉq����X�(2��F�(�,�ϩNKn*�h!h�[/k�2+]��hb2�)Ә`�BD�u�J]աh
�0�-8D:��b���@���� ��D��J�&�NZ�f�Epb�k��454c���u.�Գ+f�����H���M�{Q��">#��������k@����q>��p�}��Ҧ�����)�z$�+�D�h����ިGӊ��ڿ� ����H�qJk�s0{ϟ�^Y�ۓ�ӘĖ�>q�U8
t�����C�Bt��S.ж����4B0����    IDATI��ДN]A(��M+�M�8M����9I�#s��N4�p�ǽZB����I�('� "��bHU�^���r�N$|�G�99����{��*�8���;�� �(B��O7�Ęld0��3}�o�wy�+�\멧���������ݖ\�{v�87�N]�h���B��	rT��?�)��%[ݬ�TK��"�ӇL�Y�(��!'2&<>��-��O
B_���V�!`���~R��0�4j��Ӵ����C���.��"��U���p0q��!����M�n��nS�hY�f�����k_��S����Ԇ>ކ�&3ڜ~qd�� �n��H��M���"�LּQ3�Q!�i���r��A	Y)�U ���a�Q0�bRZצ,q~�-�N�6�S�z(�o W���ɪn��D� U��l"֨%����YQ3�v�RK���	�;���
��g|C�&���J$�2\.�(1�o���O�~�h-m⪈\���5��D�/=_3�|���F�('K���.�?SEH:Z{����9���1ҁ�D��g���*�7&1�tΜB%Z�r�Ԟj�P��UakRVBbCp�s�`FN�A���FQ�����G��LĴ��t�'�vtJ,+k� ht��)�E�W��H��G�J�MY�`"��d	�Xի¶�+]�3����iL��ij��15L��%B��H��s#�ᔮ"D��xx:,)�BE�֏�:)ȩz��8r�݇)��"���RvUA`�q������R
��Bn[ҌL���4'��[��\�(*��h,"j�Hkd�g��Po~����2Ψ��m�ri�rM���4�����k�c�S�B��!R��Z%(�;�������`�v�Ec;���A�I'�)��d�S6�S�_��0eKl����h+���~�(���S-~'G
�pi�pvtZiS�P���/�J�E�GclB��u!�6ZNS�XH"�C�-J��|������U� �E+��*�Д�i`ʲ{��U�@��밊l'U��8��Q�r�
Y Gn)~U����
�lsL+��'U�P=x>+�.D����
�U�x�����a]GtPݸ%z(�}_���{���������:?���(}��O,>z8y��;=��psu�.��n�ן�t���9��C�|t�oǏ��+��:2��D�ɱ'�>�x��J��zxz�E����߼:�6}��e�-<��;���|�ӃCӝk�O�v@y�\��|��ۇ{���h��=��o9��c������Z,�its�����j;O?�.߼�؟����_�7[�E����s�
���^�/�k�}���)�ѧ���{|�ݥ_{��tz�������{�6�\eV��C��up4o�B�({�ػ�B�|on��<���6ҿ\w�!8����_�$NH�3 ���ҝr��/�|VT:���T!�
$ǂ�c�9Q�PYB,d|�|���mDQ�����X�:I0�B闒l~��s��qu�5V9L �Sn��Gb��I2e��X��L˚V�f�bm��Xx�c�+�YW��f���Zj-��r!��q�PEˡg	�����)M*��T��t�I�ő8v����L�T��ќE�!`�KįN��SEѽ����2Znp
�#C8�����*-�u�y&��o~�tޕu��0�����Ĵ.������M]#Ro�@Q�ZQ"�h�[�޿U���d�'���hF�6���i!���3qjF��9�`��4~f���4c��kRȭ�+뉤\����z���W����Jq���/~Y�)�G��H���c��_O��Z�V%�u�Ο�㐪Q���v���ą�9�`VQ!})4���T�Bu?)~���:�2���Ң��؄�7�q�ŕM#�˛o��{�s��/z��R�&��y�z�D�s��`J
�U��7�1�ou!l�%���)e�aS�	�Tn�Em:YY5c�wN��8�.!���N�|z!�C�3̥���z�l�C�{���4�����2Ւ�������83Uq&rKQ�@0��(��Ϡ|��R:sb"pt"j�Q���Q�8z(E�� L.Y颤�<e���֏,L�i�n��j�R���Ԑ �t>+�ԃ�))"��O?X�GT�A�zЛ�����RK��a�pQ|
�����9G��=�Y����+V	!ʬ,h�!�X��F`���T|��p�5�.�kw��\����JG�wRP�cLݶ��*eq�����Fl��� ����#�[R�sVg���\�� "�#�����v�[�{:�U\�R�"�LT�o�(h�\����cS4"��N���1!���Me_M5�yY4�u M���I���l��͈\E�4:�Z�,Ác�������t%���s�@.�\�z`�	&P��AZ�(ddqh
��_5����M5ɯPQ��,S��%JJ�:�^W5��#��ф�aꐸ�*��$��\gu��2�C�IQu[������H�m-����E餽J�´�W�cH!"ڔŗh(�?��Ov�`}��gzذ�!ݨ.qP��C��BRА�PE4)X�X���K�,�>��!�J�P���\�B٘>�'+7~"�+]�%T�#.j�ι�����4���[H��I�
���u��E���z��U�.:Y)1i��0�d�>�S.*qh�)��_��r��R�@����S��"=pp�9��0��h�d��W�/Q�p)f/:"B�G���
�f��
1�¦�gQS��!���%�D�����t1�*�7i��z���&w�P3�s~4!
@�r�9����#8R
��������8���T��j�Pb-|�(GE��#��.�t�N_�STWԪ�&��DGu��8�ï���U��&�(��'�CJ����0��x�>�B��|�\��45�
�|8B��l"
�#�1�A�Ɵ�S�:���_�)g�w,8���&�5r��V!4���H���
9RR�i]M�NY8��E���#�a��ub�cZz{Rb>��� 1���٤X�>i�>d6��r[�����'e�] ����h���� ���P�6�,�P���Y�rl�k��4�j�c���p�R�f�UԬ�?|����m�:LD�)?�(��o��Ek��$�j&B��_"N>}���-Jh�G(�B�
o%ⴓ���
�j�,��'�N���F�/�݆s�M�(d(a�,Db�,DT
+D�݈Y'��p� �HY�*�$>ܨ���ʅ�p���,�������1цÙ�&.���uD�Q�U;�g��t%RK�/D�tY��1Z]��n!6�)��aJ���-��B�D����"��2w'�_[(�@"���g]M]��p� K
?}-��Oe]�uR�:OL	�{��M9����LW4����h|)�=��X!���lS���:���8��3�� ��C6�lڽ�3���ٹs�L1�I��3��}٬�<޽�}�w���/���ѵs����:W��)�\��v��c���7>���P��p����z����q};��ɿ���L���G����8����:��ŕ��o��HК��S�x~z�Oc�?��都]�,��e�b�-sE=ot�[�MXOO4�������擛��ݲ��?x��x{st|~����M��t=Q���/��z������7������g�'�����t�ϒzB�.����>���wvo]8�/ץ��馝{srts����!ď���ǝ�sp��v�*���WE���tm����i��^��#�SI'�7ꝱpj�M��Xg�)M.�s�� N�{��!�6�%�2�|�\4"�I�D3p"p�p$��I	�a��S�V�Z�8E�W��&��
�9)S����&�����)�plx�O��,Si!�z��1&�8��c-!�/�M r����JȂ �*�L�c@L�� �
��My◕���ǩz�J'eھ�C%b�۱I����I����hWM5S�R�@#�d�(́��"�sLydWɽ	b
��bF`+�Yt
�j����(�^cr9d���ѧ˜#����=��U|��A�çz�����]�.m�g��ɺ�S �A��5����L]��?��� ���w��w�}��Σn+%�3�R��6��PT9S)��#��z��B��)���J����%��BԺ_�H�	�~8�X[�ӻ���&����;�=$F��Y�O/��]Ͽ�k�vA	j�u��Z�q��
��)*��hH�B_�Bb-h���I 
@��M����$��X�G-֤w?&��DK�:~��y��?~�����_>p2��'6���c@*Y��P��ꭆi�Ƥ�%*�-?(���i���_J��Cm������R4 �a-����h��z���/}ɷ�:�����Cv�8�t�B����Y)�(�(�y,��uK�n1�h�SH]��Z����p��tRZ"%�H��[ZS�6N��N�5(PcE)�:��"��h@	V�JD�a�ZR���H�⳩�Y���7 D$9�4帰[�tC�����!|V�; �D�TBWR�i��P��V��V�,#A�!�5�(�T._n
���JC�����_3���[�)�Q-)�#�LQ�Bm�ᘤ$�Q�X]��E�D�<5�Cֲ����G(�����WH9�@mD++����"���k�����FO�-^Q��@�y���Y]��rqL�+=��^c�������v��Y}�XK�ѼQ�����b�j)�(�(�)��%X�(���M�e� �͗sZ�@'���BtU.�o�UH?@6e
�B_~��_4G�$��rm�ϊ���W���/e��_IM��:�Cj���N�#*�_!�4�C��l�|Sȭ��F�]ҫ��&H_kj����\������Ј����ß]��YJ�8������TN�Uħc��U��|����~��,�UH+��i�T�(W��rXG�:�E�t�&�@X��!��VMY���Ѧ\���L�h�S�ӰZ�P��Ԓ�㛆t8�@�� !
q��+
h�,Z'��tV�#�\�r�T�\�:c�{}Y�q�`p�&�r��+��+1$Mumf��(1�b���ʪ��)�X~)	�_O'&�n@�R}��*K�%�vS�YH��C�)����Z�!,�l )C��Bp�<N��m�_o�z.]"��s�G
�h�ӣE�1�hSn��;pd�єh�u�J�R:1��� /��E�V�9���9Tn��'�Z�I���i����+״B5�4�uq&7�,��צ�Cb�9�ŧ����j��E�3�L���-5"J�5*ʗ�~K�n{Y��}Ìc�o`�$%�ú�˭tQ��R��H���gCHM�||"���I	�I<Ptt��A���AZl�[cL����Zo;�^av����o�s� �����E��]��x��k���I>�D���r�c1qj �ơfB�Ǻ#�9�84֨���D�&�FkD�oz��|�i����9�t5��(���c���b��hN� ��Mߔ[:>�=G��ȅ��/+�a._-�nYdk`9���
BU���B}�UѴĦhѪ g]Bt�4ˊi*����T�'5@�4'�8��Z�qX#��р� p)�iB�����@L�B�����l
Dk��9|!�I%R��5��["Ũh�t4��:�`�5L�B@��N�`Y%V�B�,���E)2k��l�r��B�:֐B�����;X|�+B\"�������� ��k�ę�YIB�^C!!czF�70��Ҫ�i&�2夆�g��)s���Y�������Y�r�'�;��?�UzTy}rN���m�"�ã��g,-䈲�QO"=�;�8[����>��ur����í��i�և.ݴ�"ܬ�S铔�5�����zDyu~qr��_�u�K �V����g��OD�Z��o�N��d����ד��Sh���?�ݾ���-�^\��]�\�x�������x���OZp�X�":�.H_��M��������O����
��ǻ��WD�c[�õ�k��f�ݾ�����֟�\x��ܳ�[�3u�o��6��w��[�����4��w=� 9tk�s�H�	)/�"�"������_��KǛ !���sd�.��BXQR�L9JC��4�c�P'UH"@Ct�=�Ԁ,!�T����y.�@38@YUa�8B��%��tR.p.�%���
q�j�P>���+)֨��4�+�Ф˅�1e����MM%�&dZJ8+=�N}2�:d��%�b���DF_�A�"PcS�$�I�2�2&�ld�P:��F)6��!�R+SԈY� �F8D:&ǔ��4� |�!N�9��%�f�ǔ�ï�H��+x��/��Ȧ��D�w\��}o�z���w�$� ��Y�����r+��.+��(|��yF#j]�>��ӟ�Գ��V�C��}�{4!������7�����c���X�DM��Z�����S!�&�Ab�_d���JP'ҭ(h|���涷�=���kI����\�6P���.�����o}�[�]������YSC��� �*ƷNǸ�T� ����S�R:�E��>��!e�tbj��Z �fZT!)�ڣ��_�"2g�`{A^ߦp�ѿ<ｳq/ߺ���#"�uY<�)RVH�z�~�_ÁU��Ad~Y6�h�T3������~M�U�FI	Y����m�iB����s��oS)�]i.�v���/<�t�8�	�O'�k�%��s�� �,ѓ'�ff�u,�H�iՃװ�8����R�KG�@9��9 Xo�9�7G3e;{�-ܵ�l�j��7�Y��9��H,�tM�E-m��V]��s���('��Π�R!�����2��>�1r�k)x���'Ś�tf����`{�
|zHY�B,�g'D��P(E3tX�r��������PW��ݮ�����;n_l)�$J1��Q�Y4)��7�C�Ҟ���r�9�>e����,LE!���q�������*�8�vPz�E
�ߡ �����m���%J/��R0՘�QH�.�vۦ�$ѐ�� ]�A0�`��_���k�b)������0�Q�=	)�|!6&��dq [����CT/�r��ൄ�_�U�V�}�X���m}|]{BSE8�i^Ѷ]
��^'��t t�ȒM�.���h�� (d�r-�>�Ǆ����Ao	�JA������������R�ٕ>D�K��)V�DNk���D�C?���=I�54�"N�t��\��ڮ4����i-R�p�)����!H��S"F�,��,Դ�M_��Bq��8l'@~L~�bu��&g��lj������X�1�s��J����ű�!vL�h,���8�	6��I!'��p֔&�&�f��AN����ȇ�	���8���g�Vԏ���?�
1j�dK�D�t�
i�0�#��Oj@02�V�[iS�9m�v�h,&[c���H�_����ES��^_�?�,C�88��n�B�5��OR
�Og�8��J��b�+Wn8����|���q8�#��4�R��'�B������5�&k�H� ��K�c�� ,�MPV���G������9|x=;�)ŗ.ʚ
�8�w���$�5 l�;!C���/�j��:D	u�igdk�Z8j�/�ϊ��~>Y����^!QQ]�OV+����[�-$?��e�Yop"����)�k`���#�̪�l�R�t��|dmˍ�x�!F; ��>-&�h!�Ӳ��v�j�X?) G`u�N�u�Z��!�C<��hF 'fjt��T駵M�t{��������W�ߢ8�Eu����%9����F+�f���G0 �p EY�Q��G�F��*��B��E���
�C�(���l����)?����#8%��d!#�3|��VH�.�%"�,N�|鬨�^�8�ij|�Z�Q���&���CX�X�d�D0d�oH
D�@Y�*:?91[�Rid������#'�&?>!�s���>~��LS�t�h
�9q_ʡN铛���,Z�-�4M��ݬ�:S[1GG�S��3�9t����h����j�C�Z��چ�2��9p�o���)�ӑ'>�/�.��{��U��    IDAT�#�ϫ��	2�z@k���@ǊR���Zb�D��}_��]^����Ų�strw{��߱?����u�~����(�3��G����?ӿAu����c�>�y���Oެ�v��OF���ĈW����e����iz�����wbo<9�=��?��{�?����c�N�Nn^��|N�����®U��[�ZZq|c.���\����]����+??����W�z/w��p�����Ƕg��aw(���s_�{|������FY�J�л���V�}�}F�#��3ߺ�>-zw�f�!�u��7	��^+�h}����[�����5LǑ8>�p�C:y���G� ���F�����k�w��<�H�	)�O'}�49d�Դ�C�kg��D*�U,��V�)��/��2|:B�Ej�iô�AL�.+N">v�R3V��'2RS� ?��)60䖌\3�3�Kpz�:¬�f F%F�6��1����[�t�����o��p:qJ��нX�E��1!�a� �6��TW�&g��h��u�)���gk/�P�Qk���g�p�bu��L=�Y8ĨS���@SCz�A\,����7u]��p�EiH�^�!�2��\���z(�q�ך�^�ӟ�Dٕ�N��W�"�.�7=@��P!��*j��R�	i�JTH:Z!#p�ka{��HA�B��J�(1jͽKoh#����ַ7B-�&���(��L�-BC z7��l���ـ�n��a(LE�W�Sm�EC�u�
��qh�u2�iv��,C9)�Y�j�I%DG?�L
ǐ.T3��!Dj�Y��]T����ۻ���������_�����q��}x���{�}���{�OA��(�5�
ˇԭ~>-�8�p��	&4 R���)���)�[�ҁF"Ƚ�q��BKpV�{fi�m�3پ9�<kq�`z���9;=������&%�Jc�::�:�DQLS�:E���y��5:�M15� *W�$8K&e:Q>M ��p �)"�A��YB|�lj�hRm�2)D6���e�Q�&�`kA�Uz��B��#g��5/����
�eq��!��bJ�U��l�D�(K���i:��c'jӐ%��(kj����7��[V��tki���r 8R@�M0U�O�@s��@�lj|2B'�#[�)A���ew�LU�!�5 h5t^E�Q��V�l���:1}�ꕛ��ˋ�/�j'ԋ�����\q�Ӌ��z	�o�; �k9
���Xյ!Kc�m����e�a8i98�Z�������>����Y�)���\[ʷE-P'8��2o�|�d�eK�׌�	HPzVǨ.GV��p%�GH�҉{ Q�F�ȥ/�A줒�V����7$"k�,M�d�k�A_������mj�|�hdNj�5�y��{�̪q��$rt�CNEu�M.G��P~��8Y=�V���@8Fm�1ZNU�Ȳ�8@6gr;@�mN>rS�:�(Z��L��'���u�$����� ��859�� ���61m��&7�E`C��`J1��j���J�U��@6��/D
�T���9l�1YQ�F>N�� g�B���:���$Pnʭ"��)Y
\���u%����.���r��i���\J
�� ۜ��]Yu�:vB�8+$�H��F���
�i�\MT���|!�L��H��>�Z��V�bN��������X#}
|���sOE���ᐱB6"��d�GP�Śrj��d�i:|S~6~~u'W�ߴ���N
���5 i	F6-*GK
�@��!5��~
���a�4%�/bZ�h�a��"�qR��-�o����3��Vb>���/1���^��M�'�t �R%&H����J��e�B�(��)�rL>�.g)�O�!��&��1�!�f )
��ɖ�D���z��UX�,AQYY�J���*F(�Z�n;1k�h̢�R����H4��h!|c�ӹ�d��g���M�B�B��)p8�ȏ��&�Pk�I���X�FRe��â��b��k]�G��$�j�0;��$�-*ˈ?��V�s���c��Uk�];�&�tUz~]H�4Z��_����*5�T�Y�iT7�F�hڏpht�����#8ka�@6��R��8�t>�غ��B�N+�P]֔f�m�၃ A�1�ӡ6�W�f���� �����4)b�tQ�G
f1)�i���餝��i���A�D ߪ�@0���6'��N�!���4������;�ɈZ�&d*��)��8!��3m�@���S֤ (�14>��(��aJ���J�_�M%���s$փB�w:o=w�֐���A�\ή(C�S��|u�z[��Ϧ����(}��?���t�����CJ�a>������}���Eo��{j��M�>�߬���Dr�x�[��zz����#H\�
��d��j��>C�{h�>�S=_�v�kuz��+���NZ;o?y}{��������u��o,�B'G>?z������ԯ�G��i]�=�y*��	�Z)Kq�jO%ݯC����6�b��E}{��?�_���Et��V�ܠ�[�q���̡l�u�u�# CL�Z�w������.���k��S�1�V?E!d���5Ȫ�3S��5ɢ"� 5@ʿd!�\L�,�!�W�l��;��ˤD`��M�R��M���gW���N�0r�҇�K�O���G-�h
�R�!����(P4d��E[�QELÔE�ϒ�ɶF�&>1�ҟ~�_�&I�\9�BL�e!�������MVnE���B��8F}�Z���)'���"e�1�@Zi�mR���c '��*�imK7�*]V4��4�:�HqdI�f`�p��o�[4��~!Xn��09��:�=v�7|.ש���r��'i�|�]�R:ϭH9�B�D���ϑ[c�e�#H��O�/��SC��j�usC�
�{��D��� �.AS>����!��Jw[[��	ӕ�ל��!'Dfd8u!x�@:����2X|�k%�0��o
�gtd!���Z�|���"Д壱F�|GКX^5T�&�/��I��?��o��y��^���}v�t�{#/�;w)Ԓ>��M�ӔcX��\�xV]b�4����p6�r)+�o�Fw�㘁���4峥�d�㳔��ƢN����G����T�I�~^�+��<�$�%���^�}O�X�����Z��m�"��L5f��bvr�5�I0�9?��Ua�8_ԡ)�c@�(Lc���>�^�@"|YJ�����@Y��k�K�Ӕ�$�i�Cχ��h�:7�X�1SHdY
ǀO-��p�:�AS{���aQ�B9p�he�+xRB��n���U�F�'"�i���x!R@���j�rd	��_�i�A�c�?RrjI���<5=����І�B��ʁ�#E��ɪa!W��Ҥ��<q7�I�زt���?�Y�k�*�Dŕ�7�S��]�d��\���^���fۅ�"�Y���ttb��F�9eQ-��^��P�*�!��1ń���Y��!"X.[;>'�,���
Չ��v[��bsl���8X�����7��BF�6��bj��0%U-"�zS��;"DhvV8"8�@L�,!|!�p���`A�pm�9+�9LU78@ߐ�:�:�hTnU�u����v��k��\%���*���J�(�Sf!�)D�n�u�h?�hF�p 8c��gSF�X�#�lV�Q-N{8
t�����4��d�K��(NuY�����9�ljD0`}�B������a���5EF�o�D��W�DX:9Ȧ�>��줈��\!��\~"�R:�X��D;���y/�k�3���Ѧ�ΊJ(݁�1��>�d�။��!��E�$��3�8ړRpS� ��JK45��9�|�B���zp^)D0������h�d;5 �RW��4�P'���0����,���X'	"���~�*�b�H����Z�d�-�f�d'�P:|N���Z�@���v��T�D���!ȝ� %
1��8XQ��[�=$�ch��Cg�$u�
~H��H�ZL�ZbCV�=�?>߈��>��&�G�D�*���7m]�����r��\�R³p�p��� ��D�.	��C�����@�r��u�y��*|���1S�C:Fl���;�M���B�3��l��t��i-Պ�>�~Jl��Gkʯ�i#ӴU@L������*��#W��[��Q���sL��`�:�e�Es�ҍ�[l�,�QHzY8|��F!�BF�S"ʶ^x⋺�%M~?�$k�Y1�-J:�m�2M!Y�br YNP�)A�i��.���T���&Uo����I�[K0&B�t�B�I>�M�X�,RB���v���:�hR�R���=�©"�o��]/=<�M�[>)S��8�FD�M�0��ⓥ �aG���,y���R 8��jL�Ó*�dY��A�$֔5*AJQ��喒5M�J���g�`�1���B��]�Z�bJ7�-ĊJ1���V�~�8�|ʘM��H$<K3GH���,��p�ge���l�CJH�t���YB�*I	YӖ3�����7�F��$��V7eM�֧�(�*M�9�)�kP�>+ŝNvB�q)|.�k\/�>+�X�����j�������˻���㳛u�=z��5�����K��J�KR��cOO��_Zq(|��7�׃��xf�����������gFώ�����I]!O8ן�\�q���g�{j��k�YM�n=�tD�|`'����=�|sv�����������������[W��|x���;��!����|�Յ��}X��M��ʭ��ky�������&��Kg}�Կ2�]�lD���O��l���8R�,$����M�n_;���O)B��їh-�������|�����7�\)�O~����ٴ,|Q)�p��f��iњ�Se_�	J7j���!�Ф#�
�)�!�J�R�YH��qL����N'|��,�U�Ǡ�`�\Q#����|��!A�C�8�`;vuXi��8� 7��0�n
4��Ï��2�o,����9��QV��t�Nz��J�B����S����� �4��;Y!�`Z���uY~�,���)'�N�|d!�A�Ԍ�Kld��,`বE9��5G"� �D���7-q�(|Z��T0]�>��m^dS���uQ���T:�\!4�ڴ1�h�M]֐��lt�c(JA�>���K"�@�-���D��s�І�r�B���ͻ��,�����w5Y|֝��i�v�˝y7�W�y���VPuf����TX�6Ef5jOU�����o��#$eDi
����m+k�5���i����(]3�)G���L��ӭc_7��K���}�;����������~����O��/?_>���/�ғj�-���BJ�����C��v%?_�������	������_	>�#�&�(��f�D�6��2#�Kt1�{�szx��O�{�q���^�z�#�=eqM:)��]��[9S���������h#BW]gEYvO���4kJǔ/���9�z1)'�`4:B��o�@�rE�"¢�����Z�|N핎�C�t!:8�K8��rz���iR�[���)J�}��[#�,��G"P
��V9��!.7��B��|�.
�����٢ ���d�R65��RZ�s�~�� 'e!CV:� �Nc�礵pGn�\8�8,�=Gh���m��5,��,�!��;�~��(�.q��N`��eϕ����eEV��CPZ����}��=�.ISׯ�3q��.�0k-�R�W��|�򕯐UŔU�U���X��C�H�d~�p��Δ�`h��d	�"�
�C��f��;��֒o'��*ڍ��{��-E�U%���!-�!RZ�,[D�N�6��9R(������_�hJ8p�B�;���^Q��\!Y��@��V!�_{�8�*��C����x+un��I�Q�d#$n��_��Z�l)�(Ĩ����E1Y;�� �kj����KJ�DhH4*ׁ&��(&<���)��8��B�n��G��`����DEY���d�
��"��I�a��j�?����dCȆ��B�$"�+�ƑH�'��V��9D���с��h�V�� MU/�7b�2(�ˏ�Q�5B��r!�aq�Ґn M��p�@j�+��إ/�����dW�].(kh�@:BYR#(��
u�I��J k5��f��*7����ѧ��)BS>#k�ʭ!��{E��1b���7=��C��M[Gc�[u4�R8�YNj��M��"r��L��yj�Jl*���4�a�Z?�j	Y
����S?����ÆU�4�E��� �S D���C0%� �~�1�F�X>�p4��l�z��nZJd���sFs+�e��
՘\[I��4(ۢX)����QW��bE��˭�,>&}�S]�,�D0~Y1�/$Ŕ�P��@S�T�תK�h��8�V����2�i~4>�1H��a��%�٥�H�3�)7��L�q��D�lk	�Ȇ�9�\Yր.?0Y�4�$%Ŕ_E�55�iǅB��"����Ҙ�(����SB"}Y��+�p��kf�B��KA:��Hl-U����D�W�cЉ�/�8�(�SuN˩V���Cr
�R-�
�hT��lf��k�
�U���;��#�VhB�s��+��4)E�P|S%XS|����e�C"�9,�/Zـ���4"���V���C�HG�ٟ�NW��]�b�f���éV�I��(��a��	�(vF;���D��j>Y8��#��6+%0r����3m�l��D;\Wj���l-��-"�%?�h�r �&YP�,���0�9R�������0E-SxQ�NU����v��+��'�>b�����X`��O�������������{�}�칏`z��I��<]���7�jO0�}r�a	�^���'=�<>9�:��3�6p!.Dy�#OZW���ۧǮ�^�S=Y�j�>����»�doW��ԟ�D�!J=�+����׏.�ή|�g�g�mz�j|�����/N�,�/d�8�\���G|A�ͩu�g��n�;���l�^N�_��Ǣ{{��H����j�m_h:o�Ms�����2�ٲ��+������K���=��G�~��r�'r���o������1'C:W�w��Ia
��l ntZ�U��
Łt}9FS�����T��Ӕ#�nS'��ݔ/w|�B

Q.W���h��Su�tW��j�R��h��T��fM�h�����>��Q�4G���(p��zY�Y�mJ�0��hpCV|)|��d"Ә)�i2��)�T��=\�ri�m��PoZ��aM�e��O*M)�9���.M�74�:��Å�B��6�r��a��	�S�O�fLS`�Kti�z��=X/.R4�.�w��ݮ�W�^����o}HÛ����Ȧ�Oj�ȡ�z���4(�5*���	i��q lK�T�$e��h�4	�GS�"���q� us���5������4���I���D�E�#Ŵ����gO�����T9���sM}(`%;�h/��*L�"�.xre�Gӊ��FnBh8�7JҀP _hJ��;r�`��tS�ьV�|x%ܫM�����s��B����������������G�����oe�~�>;��E�2a�-�=*Ѷ ��`Q�vl�VT�B��X�f-��Q�F�������&�N"el��ʹ��j8]~����٣�m��g�!.<��D������rQ4��r��e�;LJ�'Kg/t�VDn-u�l ��=��3{� ��N�0MɲmAS�8@YEM���� a'=pN�t���|j9p��� i��=�ȱ{h���J���&q:�[�D��.������"kj�9�1�@��0ʲ*�A3���2����b���dj�E�T�)_'�ǉi8�p|�CV��@��e����9��!�u�H$��$e4>K�v��b::|U�4UD�lt�(���ip��@7YUD+���b9�D�@�{7���.=��g5������D]�uKA]
1B뚪a	lغR��ׯ�w�yG.<�6D�h���"S�2_V��䰆�8||�Q:ؔ��
��:�i!�V�HAL��p7����W��)h��    IDAT��r�i� ��6���(��P+"hQB��Bj�� ���*���D��
Q2dIa�@ǝ߱�P!�r�l�&��BYg"����X'tt�Su!L)������55JF0����h��6�Y��(p�hR�B���(S>�P���D�X�G��jv��*h�e-SV��OsjIQ�M�>Nߨnm��R���՝����ǩ)�n�tLS8��'���A���,<��-jQ��9k�N!�q��;mB�ҹW�s5)Ȕ�ϱ�[=�Ϛ�$���t�RE�Ayh�CP� �IJ�V'򔼯MY�1�\(�%�&�p!TR	SqH��+Z��Q+�	�CH�W��D"L-��p%�_�	��ę#<H���k�ö%���,AY>2�a?pHuE�h�:Ѕ��!~jBr1������"��sC"?+iګ��sIT"|��x�!��D�]���a?2w!d
)�7LK$X'3͙�D�%dt}�V��i�>���cZ���/���_(�l�B���m;�Q�
��i՜)i?2�R��Z�8D
�GhW��S?�˒2�R�Blճ�U촁��]�I�˅�bO's!8M?x�K�t������ ��eG�h��B8p���[f�Db�Ɣ��7��I�(*$�X֔�Tq���%���)���l��~R�>Y���d�F���vGA�Tn�Ϟ���t(��B�6�mJ�guBt�tI�>�4��$B��vǂ����
�(J�T"d�SK��!�J�`jh�ᣆ`HAk9d W�ߴ�U�/e*"Ԓ��r������FDԈf:2M��AH��T�sR'���"T+��F�i=�� �=��jh�d:GA'�dG0DE|#<A���,߈��/�1���Z�}��>�pO0'��U�n:�B1Y��?|�|)��O�����z�xᢔG�����5D��
!������[
Ĩ� Z
�z4Mv�L��1KSW���LE;����@#Mֺf�lZ�_�(�*�9D�%��3�/��y�ɏ�A�cx�xd��(VK1K��+t�Wn����չ>��c�被�c�\������|x�<;���r���z���N�}�S!�mna���}Ucw"���G}���s�n�>\I���7}�����{n׃SW0}_r�Q�6�=�˼�Y!��w@<$յVW�뉦�.�eY�����xw{z�����_���i�?\�L�{�����������#���{��'<����ۗ��Q��l�r{z�G�5Yo��z������>��_y[����ص8m=���6}�Z��Z>;'N��y/k]Al:�)я"pj޳�ȏ��w�}��_�2ܩ��{����jֿ����"����&��~�JP^����B~X�a�(L�,�,ͭ��P�Y��r�V�6m�+�H��D#�a'�H�8@C�@S:�O\(<�����fj@n��U���@�Bj��E�1�̶!r#&?Q%�M�U{dR{�P<A�(Ԣ�)s�E%Zc%�?��F��ä��,&��4�)'PT�i|-�+��t���8Df�ؤ��c�i�����-_�v���d�Ō#��:�ND�w��
I�7j� e
��_1 B�`�?�я .U��}z��[��^���o~#�ԛ�Jt�R�n��h�������F���?_hu����U�����R����P0�4ʱ�5Cb��ެ��Bp�����#��Չǽ>��}N�&�"���򮸣i[�����z�ԙw�}��V� �R��O6�!wFc^JW��h�Z�3�4��78����*�ax�bH�B���0"85�ֈ����O�4?t��z��/}M��ĕbi��������>�]��__���>��?��&�!{��O~v��Bv����C �%�W�*BZ�N]f��2��:�q6�����E>t0-Pz:E�Ӝ��#k��3a'���G��c���L:�霓�:�<����|��g��@��<�C���Ƞ�ZD�����Ne���|[��'.�PV���b�O���@6_�Afs��-p�d1��!}Z��k��7�;ybā#l��fv����9�lxu!K��!@�-h ��l�݀L�A	4p ��k���âQ�1��vF�R0r�Z fYB8��$dՅX�z K�,x�(�͉��:=��4>�tgK�D��e��
�R��'�*8��T��1���׭�������ǯ(�P?�SG� �I��q_��a�<��������&ܽ�=ݍ������䗿��>	��������)���*�Hi��==-�i��5�A��	D3L�)1��5FA:��Y�R�5���h�* ����B8v�?�M���8��d9.�B�w�� Ǩt�U�&�RߣVE�Ԫ�d!��SV�QG�$r�b�Tb��#״ܖ �Q���+����.�]�ڬW�2Y�j�ɆĔ�Y	�BE!��Z"�!��Q�c �)�NB� �S�HI�,v�<�Kďc**�Q߀��`4x>+
�߮�>�P��,�o-9BFU |�[�П�J4�0?�EV�n��g�_o�6L9Sn��g���J�ҢU�P8Ut���@�-�Ca�K���h��R����C��G?�@�)c��,)���ޔk�\��Df!�ҍB�)�B����MT()#^-|N~��k	�0�k`N�*��*� ��\����,��U���R�uDҬ[�,G�ֆD%��b����B�f�I�Pz���b�k	��%�T�����Nh�V�2��g+�ZiV�0͗K!��#�)d�lh�ud*X�,Z�|Q����%v�qZH�t0�7Q��Q�;:��/*�a���A B�駣�B�UA�"d@�T�8�餏̡��ӶZ��*�H��@�/�% H�a��a�l Z�Ԡ�V�U�E&R9��Y�OVT�e�!�����*!��E:��&ה���Y!h��>:��k2�şC����dńs���p��Bҟ�J���зRL��ó��)�8P:�Dk"��~ҟ~�!bZ��Y�J��&%�d���;����HEMK�H�G�
��t�Y���2�� N�uhE��a�HDk�l��ф0�t�RK�W�= U��h�%��-kh�rXY8�ݐ�*8�!r�dk>�����(k�&�䑥6�5,4�d�����Z����Ղ���Λ��pJ)+Y3�eC��P0=L��!U�$Ŧ0�9X�=5��0F6�,�S�J=ԏ9�]�C����Ք��̖Y�����9�i���#jeA��THHV �f&�D �sm��Q�������ϐv��t�5Њ��� 7�E���&{g@�ߘЀR�m�`*+�|65 �Y�$&�Y(�VM���M�����A
@��8unZ3֛H}v��k���"1B��ppP��>��7�{?a~��[�'볓�*z��e�o|x��{b�D_(��^�֍���7P��#JB�>.�?��뼷\��?&]�ܿu����~�����|�����������'w��'>��kj��꣟�g���jT��:�;�ބ�ޮf�欳�a�����ýǥ�>G�Oy��ҎO����㫏_ߜ]��~����Û�$_W{}s{}��������;���3��?9?z�Orz����uݢ}�m�r�>���=v�����tr��?d��tgX;���۝/V�dN���|'Ǿ�@\G�>?����/��aMo�����d�3�w�zݤ�=.�.�N8��Z�G(�Y�}��[Ѐ��1u
��!�GçɁ���i�bҤ��D1�xӱ0�ZB�)�iiʢ!�a���j�-S"[!-�!��Yô\>�N
�k*
Q��ÓmR��T>��|+-����Pcs ��F��&R("�Se4I�K�j����W��#s��U*$���FǝC�����#�,0gĞ�>2��R@�]�i5���Ґ��@���V���R���KA���B��X�Nz3_�E��oۑ�����
��7����a�~�i�Hg��U�F%,���Q�z��M)sZQѪġ���DZ ͐�T����8Ǫ)XT�"�ꔁ^�9D ���z4L5�p��m��7�=��F��Sb��{�iBKNЁ!�.k�Vh�Iu9>Y�
�H���NMz
mD��������ɵ�a�OG����o����c�C�+������]/���������|ݭn�s�;ߋ������	���?����/^�����b����C�����NbCi]�D���f���֪4Yl>+��iH��W4�c�#� S0E3B������8���˼\'���߫��v~$��
H���CM��'�%����@�����,E"�������:�.Ki>)�Kѹ,�����>�1Cp��4����l�M�R(����)�~bB8�19-�/D!�|u!:�ܶ_�_ȴDN������G����x޳n4�3G́�B�4/#>:_`^f� <@74К3�]]���y~���FLW��|ٲe�="�bgD����٪iʅx�R�b`������FSH:>��ݸ�,DȦUgd~!� CX�S4rS��XSY�kh#��Q����5�V$�t9dB�1�h�f0+B0ş(܀P�	&�NZ!/<�R�7��#���h�|`L>�P�B䪻�:�@�P֌)MV�=��?5_����Ϊ���p�����>���O>!h�
A/~�Y:|�$�#jH4jL�VQ�Bk���!�˧3��=�dM��p4"���T'�����8y&1%bګ��B(��*�p�ir�pd!�E��%��㄰����(C	̎qC�r�rZ_V��ק�6��t�Z5�t��D0)d)�&�ٮI�1��)�8��� �r�E�ϕ�1S��:}LQ>�� ]
~+b�+�BD�JD68��*�h�8��i
D��=8N�2eK��W.�8�%ʟ���\T"2�#���>����V,��B���3�"�b�U��t�$�P��c��0)ũD
�E�t%+�&D(��ȁs�"Y�/�c
,4�9@���S�����'b�SQ��4�4iJ̀�H�e(W��%�9�EJ�O����P;Ɂ �F�JW��>w�!FR㘖��	�?uU����Wb�Hk�Ԁ��lN>Z���@�BDX�7�0�O0�q(�˭J0�v�&e>���)�SMܔB�Q��
��I���	l���k��$�W�%UWY�%��%JJ��R?Fk��bqJɯ��LC�(��K�kT�c���)�qT�&ʟ�4N��sȶ8U�Bt���9��&��^�Uw�EI���B-J�&P�0����>^w�Z*��lu�
C��HYuXҞ�[.��>�,]Ad��c�Ŗ��㛮�۞�b&�/
IR?j�CL�^_0�����|� �|�܊�rX�t��tYpY|��BZE:l�1����N�jIo���(�n���R��_����n�xά�Z�G�%����L._�@��U�1�R�L!�P�Ň4MB�~��EA��p��io�
�L���O�0����ó!Zmuᦲ )TQ.�!�ω �O����J]�q҄��[ru'��jIW%�,��U�/��4�4�/¶6+J�]�V	8Z�S�)���>ˢ 54ɖ�~B3����K�VS�VڔO<4A(��j��e��uR«������d�J��:���|C	Y�9�Si�N\wxo���3Yi�-:�p�)�2N��t��V�7�"Y�!đ�"�N����� D�#�5�sd�O�� K.��Y�0WCO/Lh�b��k���_�K7�N�s|�W �7F��Kߨ���Ӗn�}\qr!lb�֗�>��YU����i̫�뛻�,o��ǌwV�C��m���-J���&����7Ѻ�����ۻ�_oo�=�<��ǽ��n}K��r���o֝V�kX�Z�m\o��e}{�����[��es��k~r�ӗ���v7>sI�����7�=��M_�A��O������no�����^Y۳u���p揉��KwG�#|�u�`�w���s-��l~�ܽ>�������کZ�����3jg�&�*�ܬ����	��_��ht5��t�·�����޵Ϩ|����N��߀��C� d&��!�,ʙr�ԉ�{|���!�Ve�d��媳uV�!]
¡@_�Լ��o*����TE!Y���h�Cy�U� A���M�B��ƍ�z0 p�J+)
|C	C"r%�)s��2�/�W}J��F�\N����t���.����l�tRue*�_�Ij@!x)-�*p�JC�l|
�ڈl:E�ю	��F~�f�U���R88�j5���Ҁ�]Y�(�)'G��؎�9�Nc�qZ�*�3W�SiNS[�B���B�Bu"w���b��w'ϣ��ɺ�����-O}��>E&�;���M�T�N���������*Z'v���������G�=��[#�͈����c��]��v��� ���U�\M�B�
(��?�K��>u�-�������w���"���jkKa���(Ғi1�tf=�F��"�L��f�� ��@�
�EY�J�[m��p���[{��׾�;:^Y�Kw}+�Oj�_���.��n����nXno��ڸ�����͛���O/�~��۵'o��t���F.����"����h!Z���d���� �IA�M��G`G�D�QQ>��(����EM+�&����������·�����
j'I9m�����M������ٺ����FK��d=zk���J���!��C��`C8�5Su�8��YFғE#����X���G�� �+�����@ـ{@لv/DY�(�p��@���S{��p�9��F�r�rk��Ș�%���<��Q-֐N$P�K}���6�I'2��LmUݚ�2���퀉F�iA"�r��FOVz�O4M�{��C�n M��4#Y��Y���a�G����)P��j�4[h�Z�\-�!����*~���ϝw��L=};3>z��?��w�����[��<��SJ'�(_�o���7��駟"7��t4Ci�����@�K@[o����'�p���.��m��1^��B���C���擵��)��e�r,bJӾu�S�Ԍ[����i����Lk�"2V��O�L��8�,~�ܱD5F_]MC�UR#��(\�Z]S!4��8�ֆ\�R�5Ɗ��=��VM�#԰!`�2S����#N9pԀ�r�*aJ�	Ѷ���85F<0�J��|�)Mb�"�)+Q���J�RF0L����h&eZ3�6��*�Fph&BVV��D���R�Mt0%�]>�X�r��ӬC��H>7�\I7��օc�R��q��vq�MY8;fY���AL]%�v�Ь��j���q�� �%�3H?�Ґ���3F̦�4��!�NrDc.ƶ
P��<��>Q!=�9�{ܒ)�Zp��U`{*�l�09AWߴ4�,�\~���*�1�Ze����r��q�.
��V��M��qu����R�Fۥa����sRL��eZG4���N'p���Y��ǹ	�}������Ս��h�n�LDJ�Vm�)Q	䑂�5S�1n	
�Ԍj�r�-���4M?ǋN;0��z r�-?�QF0D�5/�>K��s �j5>�DҗgM�)�T�Z)�8���Kl������*H�/�r��	�a�6G�x�ӛ�&�!�D0��ZrS:4YCJ漓� 1�,�����b�Y����M�є�ɧࣚ��Dњ�C��劖��(5)Sn����1-M:R���rL��iǒ5�ǉ��2�4e��D��B%� O<\��)�-�Qz�S3*��V�JH�&=Y�Mjd�N!Y����1��%]Jm�q�����u�������Ш�� ��6D�`��Bh1���j@9��i̤XR���T���%����qTu���yL�tX̲B�ϐR55H��i��@~xY�=	H饰���x镐�.$�ȁr���D�R=��)��"!Y�:I��rhq�h�p����Ę�3�Fg�S2V�m$��XV|r���)���RZ�(��1�;8]������s蘆�#�ǋM�?)U(w�34�I��r�*��[)��E��nj�a^i���x[�T7�� �);|���Wȿ�p 1��Y!�NĐ��ڮ���ۭ��ۏս�Ar��� ���z�S�-    IDAT�鲺w��X�����އH�ٻ�n�J����Y]�d�߹�ށ��A����u<�;����֍ջ�����o���\-L��z�����W�-�M���m����}0���%��vi�_�1��!Γ3�w�vy������W_x���/]|]Ỹ�\~�׿�ݾ�����|��|]D�5��:��d����Z��W�<�~�#4��۪�X�`�q��{~�eK����=��
9vu-s��]�,rǣ�)GʶFyK�{���a�W ��l�SA�%U�C"ˑXK�~���nĭ���BVQAԟ�i(���4�Q�54�A�����8��g���h�J�U4d)�r,D4�����Ik��PY��4=pBL+�ԈO'%4)ś*�z��W�����I�U d�Dj���WK��r8BI�8�G��YomN���18:��B0���E�)T42�>�҉<�qZZCT�g[5�j�k�3r�C�9���>ʩ���KKV�{������˩�ކ�Lީs��{��%Ei��rGJb癬�b���Q!�WZ����b����Q�I�_��Si~m#�Gԉrd�TD���M+��2�vu���n��,��0��`*�����OQ8!ȩ7[�y��6P�uEh�a�V���RY}� Ǧ)�iǰ3n	���7��|�~��<��y��և�T%mj�]9��Q�+GQ�a�4e�D�EZI�Y@��9��DR��e�MY����t��[߁pz�K��z�ݺ��@|�p-ɓM�r���a��<��'W������7}����������zw8����^��o3)��gk�ֶC��֦ժ6�@��*k�!Y[?���FhE�u)� )��%��f�TD�˲�ES@�'�������y^:=D���);:�+ŽϮ2����a+��1j�Ť�.A�a��%�U�N�y��C�Q�1�BX�L�c��!��p���	�S������ZRZ2G����˂�X�'K��� (1��K:Z�7"���A��hUA3��^E�ކ�A#e���81g	hB�&�m�I�[3Ȧ|��q,Vn.}�"�EՂ�j�J��'X9�MVQJ;��~{k3�+Q8�+빎YLN?�a�RQ:@�ß�����B�1S5Uª�`J��5�hG�/�r�EI!�MO�t��Tl:�z~��7������
^}=ɛJ�o9+���gHmP3���(�a���G0�l��E�<Q[��#�I$eӪ��4�5oC�-��WZ	S[��Z)��W�xfk��0ug���oOj ��v��D�m"E.D?��64`�<&����(�*�QԕҘ�ʅH��EC`���4��QK����R(�qS�3`��[)�a�)����ch�T!��@84�-� kjT�5hnJ���N�A�tֈ�V�z�S���M!�g��&�VKb�Yl�K����MJ(��$«^V��EY�T��M�r�D
��(��"�fK�Ɯ(2_Q��o�?dM#�zG�/_��/]��$[SY��o:R��O�9Qc._-!�2�Q�,�@p$r��ve�ǵ���UH��tHIQ"��a
��/�m)�e&U����9��1�|��k�����D�sR�9��6��0$�)}x�l�Bؔ9U�TE.���,�nKO�EHm4�9V�ꁕ�O��g���
q�����8��D=ׅ��(�*��)��8��ueJR���c���Ya|��q4B�Azm�R�7�����*��1��#`Rf�B����
���Ȫh�R"�#q8�8����3������Շ`LN�:1հ��J�H�@�:d)��sR �����<˵�)W31)��BiXW�r"hNf�)a9"��|*j#?Gu��T�U�\x���e:�E �˚�MD��%b�q�D��s$"HQ���� �Mp�i��Z�Z����jZ'�0�L)w�$��G��
�A�	����~����Tn�8MY�U�S���ڥ���{tp���泃��W�O�r9�i�~�R4`@XW*��I_��	�Z`mW��Y���R����p�1%� �H��|��P�3&�F"1���#�S��~��oe��JS�Qb���!f>���h��ʩK��	����ka�YRഗl8�� ��"���h�U����ȓ�<�@~%�M���#�)G"����կ�Ȭ�,�R�+[mJJ���J�kb��	��t����4��}�K��ڋ��'
���LY�ԲDґ	��_���sUWV���)M)���i*��gח�R�����z�#"�l;d�|���T_�[W��g}�Ѷ����n��A���ԟ��qF��;�úRnlv>[�������u��a�
��[����r���7ޮ���<��QQw/�4<��z�X���ۙ��mi3<�wx�{l^{���w����{W�S���G\^o��l��	�����>wy�S����n���..��=���;~'g�n�^_]���[�'�����K�ӻnn�n�Y�ˇ�a��=c�P�{ ��|�t��ՖV�m���Ķ�
�� ��LLc�����ӕ��{ @\��/ד�7@\D~UR�'+�>�3��i������U�ФMcrъ���:��l��@�eqzM+$ţCEkԆCXV�Q8��49��lJ�l
�Q)5��F�w`�4S�cJ� 9@ƿa+��P���*BȪpz�Q��6Ko��ƚ S��X�,6P�*F��[-�:�#�Hvr�a�F_��c�ȲXR�ȥ�U��1�Ttd�m��R�`�s(4�[>�j��`r��U��׺���h]�tX�(�壹��[�����
!H�t{�7`{��I
��a��1=�XGE:G
��*8>	��u�����"��7�|���6�m�)h	G���W4}Rt��@F��_�4o� sRF�I"�i�N�Lǔ�C��NR�#��8��\�7� o�/D��5 *��h�>С�f@l���x#��J�G1)L"������?^��z�!�eæb���)�TH���.�Z/���R�'���JQ�����N&Y�8�uդ�hBj�9,M�J��Y^ur�"��������롸��3���zͼ���\�n__�x�swx}󥋗7��}�ΐץ�]oZ������6��4��R(�-�V���,��&�ӺN�c��B�����R��Volx����L��������=�D,J\J�l�Z��]u6>��S'��>(~����9Q���Uԡr�	���(ǋJ����V���hQ4�p����r0�Q�DS#��!Y��b-�8uΑU�������%vz�k*7k'�@G�!D
�g;i
�\�L1� �b]a�m�\_|ՁB�[2ǔ�)��C�d��V�%"�xN�%�}I��`�� *ѴW;jR�|!d�`�B�̩�,N��������/� ?�1�j@ԨN�#=��!�*�"
�(G�Z�*��1H�p�8�����!�I� ~��'?��4Y=
L=d��z!�����}�{?�я�F��NQ���E� \z���USH'��@<h���.�C��1E��a#�|��5��%�"&.�\z�p`)��
a��x�Y:��X�^wsJ�7S.��l�X�@�p���@�@���m� �'KJ5N�JChN��zu!jLb���>D3�4Yb�|���p�=�X��Rcq�8�r$|2أl�ŧ�����QJ��������B�E�2�.>G���'|�W�l衔㶅�C��oɢ��M��L�ř~Ъ�H�(�&��)��l�\S��E�r�D�4't�1H>��1KO��Ʃs���1gWCL�YY��jiE��5Fc�3"��JU�-�D��}��!3Rf%��Ԧ[S[ʦ,d��D$���k:��q�p�d��!��Q嶖
�rY�����u�S�8��@��*Jo���M��K�&7�24�Ҁ��A]�	��7-�eb�Y��8;�RJ����6E����Zb��*Ƕ��U4B)#>@��S�%�p�ކ@Lqj��C(WoZ�'�h��������,N��,2A�h�kjD�(����*��6Z���Țn5�y�$��t
�!4����GP9�'@L)�Q���@Q���7��:Δ�h�H���)��Rz�AY
5�j*�	��T�4����SKPJ����9�eU´DN)Bu�0H:�K�u�䲊F�NC4Ә�@�z�:�Q{�����V�Dd�9�A0����.D.G��Sc�B��:�*1����cLJ��H�$ב�:��!��Ij~fhK�I�6�V"��hK9�ÊV%}W��r��|d!���RyZ;D�c��t f��D�۴��~��c���q�r�E���R@8n asz��PK��M9~8�r5�!JJ{�VYL��p�@|�V!!N�� 1٦�)CL��4L���h
o*�X�Ԁ�tҔ#�&���YC�R��1�L6~dxEY���/�oJ�X����G��UD�JL4C��WW��Z��8�����Jߴŧ��1Y�����pj�������m�|���@D�j��@��YH��q��YH�l�&��ܤL!u�_'�:�n����>)��nZ�z�%S/Ǧ�@��CDT�B�H���r��f�X��e� �p4l
/��z�ǧ$�&����xh}��ڰ��u+��ħG4z}v郒�W>��ޒ^��N����5MO)>h���gC|��D\+o������>��g�����m���ӛ۝�m���ޮo��=� ���g��>߾r���CW��5lu�:���+��f�z����b��r��sxΩ�w���\>�����<w�r}����#��gWnΪ�>Pu���7��@��A�ۗn�:^���$��<�C�퇝<=��Z���A��r��趙�����w	8��@@S��_�G�qہ��*����l��Y|�����fT]���7c�L��a�?��ǩI~m;f�h���b}��GB�o���K�:�ޛ�y�������?Tδr��B�!�1QK`5-$(���aj��z�O�oyY/5��H���+��9�G��LUg������;ހ�Y-�m�!�lo)
��kR'���QV�@(hM�i@n|K.�1*�Ja[b�H���49�bZc�4P:gka	��)�kJg.���=!�{R�VߔZ�Hw�iz�JT|N�F�� ��p�c�I��Ɨ�ܐn�	�<�X�׿�5�M�㨂OY.�(���?�c�mIKc1矟>�X�鰦�4F���\N�,n��\)|"eqZ��	i�p��==�0�9EY�X��8	R�yg�p4�os���Ǆ���j�$��H�z��'��=L�0�"MQ4�Ͻ w�.���Lݳ�o
��b�|�(@��V�i��$:yJb�1�����VD��TSm`���)��3�d���������gkg/5��/}ٟ��-�^zϷ���s_{�ڷ	�'Y��ߗ�rwqz������p�r���__��|b���ŕ/#X���^��Z�:��r.���S�59�*��B���a�o��O�Xp�e{*d��IG b�T[m^h��Dk�#��ݑ��언c���V��M½\������9��D�;Xt�֕UȆH��!�B�5��*�։Lʴ��IR�8��UKg�*"�����δ=��ieK�1,��ɷFdu�hKhW��B�3�G�*p�c�j�&��\kji,~��re���ͯn~")#4e	J7�U+^Q�Y�l�?Й�@� ܨxu9RZ�pL�I�M�fU�H����X�8=-x��UM��L�����Q�j���U"� �=���&�����D��x�9]D������ ��W���'d�`ꄎ����V]o�MB0)`�����T��3K ��V;P��@��h�?q�[x8�@`���Η��)��)EE~�ê�&�rbV��.���?�c��Z�[�m¿����ߢ��B�S�-{��X%�P�_�&[�t"T-]I��Y;�In��d��4mV�m@$J��Q4��젢�hQ|�]k�i��E���E�9��VZ��S��ʚ5�۟p���I ��R8Z�>�DL��4Z�VTz��km.(���*���S�m�Kj8p��Qz��Q"+7B�(��1�e$in��g]���_�`�)���rYm�E����[��c�d�)�S%-�
ɍI֊��|N�1%*�ZY��]���@U�m8pNB�T��R�㰢���D�,[Z����FM��E�.ō�Z|"� ��%�s��K7��N>�+!)���@8@Q�6F�r4�u�G�m~�VQR�P�4p��v���OK�����o#! ��/=e6�r�H,��"B%ޱ���W������:�K��kɴN�ͧ3�W~N{Jo���f��E'���^'Es�,VI峦�sj��|��5�'�+�dA*/��(鹨*��m�rF�%�i(�ZQ�b�sTAh�*��mKZY5i�`u�E�B��@��,�ٙ��i���N�"���,���1�`S�5�J	� �,�#!��4��R��¯%�5 �KO��S� ���a:
Ä������R�M���d�b���V��,NS)d��95��dʵW=�Kak3�,�C�`
�i>r�C�� B\'�P��12Uʊ0
���EV��mɲ0��.� ������:��U�-�r�b	V(\.�@�pR��-A���t�|��J�+�?�i�p�@��g� U���s�R��i���Z*ｦN���į+L����ҁ�b�*�Ξ�u;W�L�Ia󁦆)�^=���(G(��JކD#��H�&�A����̧���кX�Q"Z�)�4�i�cH��oE�!�T��X���ǽ���WR�Y���p�gk����9�DԚ���׫���[�QK*})�*8t�+�|�=O��%Tz��S��H1�h�����US�Z�9���hˡ W(�B-���@Q��2��p8�AG�D|��m�7J��>�����w���h����K��`ݛ�Y�~�w<�~n���b�ܯo��+}#��t�Ї.}g+♏H�NW*�����d��v��7f�<����n�����joO|�ޕ����?���n?��I�{��t������v���3�H|zҝL;�Ki׳A���ڇT�;-����/�����oީ�<�>�������pu����܂���?�y����_�ȗ�z��o�>�P��>?�^�~����77�]W����'e��\_k��u_t]��ӫ�2~|z��"Rl>���+�-��8�-��XhC�J��y 8��öj?�&�e�Y"+�{J݄�aRk+�g3�t4��(�u�����% 5��\oЙ�Z���
��g?�W:U0�
���8�4)� )�����Z�P��w<��&�ޯv�Ã�;!�&kS���韼��rս��ע�yzQK!�-��AS-M��D>���JH1m	� ('M%���S4�D��Di"�%"�Y���Y
ͪ�I�ю�{�Rp"_늾ͱ�B����s4���r�\P����H��,��|S�iFo�1\e��(�5P?��p�.K�B�B��H�4���8J�K!,�Q:G�ETȢU�԰|L��v&R��Ӂc�(ZT��LqQ��8���9��c����2��ou
1r��}4!]Ub.M�M)Q�~��:�
��i*�f@���D+��_	���)M"YL��S"+����zx��W���w���[:z�X��!�Q���;�!�|���h�������)���$d1Zi�5*�,BjWImIo=��F������5pd�S�i���mHWNRj΁���''Ǿ@L�ov�����u&Vc�G��ׯ���|�g�(-����ķ���y����w���~�鯗����s���o��oV�󥨿$�^�=)I>q&��\�`��ajf�a����]�+m;�A�h�@�����RR��D(˙�ALA3ڋ��N�q1<��n�M���U��p��!����b�dq�ҭ��5�<ȩ��!
�"�M��J��4��Mu���,�NN���.AY8�>� ��Z�P">[�v�K,��%E��r�K���b�~%��|d#"7�$j����U{��L�g��`*���@�e>�DL~�AF"��c��4mE����l���JdEqh
���uP��    IDATq�*F����F8�\z��
z0U�>Y�EJ���R�[,f)��8ȪIg�ˁ��#-��a[u4Sk'��E�уG��@?~�Ԧ�u!�y���~\HM- �rq�*��{������/�"Yl=H��ز,�m�^S4�c���ʧ���b!��9l��-��CXB[��h�Ԥ6L�F!�)�<[�I��L����B�\ ~K7�T.�ZL���'��T:kZ��6��@�h����
Q�u�E���(�FMb�h�%��0YS/��=�k"��8d��r�I�P�/��FB�F
i�@�*����u	�8��L����(G�r��"?q�F�Ud��)�M롶��K����R��������dK�j�*W4K���B�рr%��@VT�_{��Rk�,�!R.$��r|!�T�4�l���jۨ�ԀA�¦��2[�d�
�!R
�P�!8�ԀE���s�[����)Hd������~d��@Ӫ����ґKG�x$��V�f���/���L���HgR�7��t����R��{�r��5��)���9���BC�A� �B�I߂�?��%Fk!��Y�B�`j�p�v�N�8p�DN�)'���ζ�ڇp�RؒOԈ���?��$BP�s���u�^L4#)���9
	U��|���K�O(7�o#B� ڔ��)ډ�����ӗ���EiF��_3٩�._�%K�	�c�3�C-	�V�DS�"�J�	o-	����3�j^.�ş,>��<S`�M�9D�㳦=�JO�O3&��v��������ۊI�Hmi8�!��"���M'� (��b!�R�lW),�͑H�Z1�bU$��\Ә��)ć�߉�bU1m!���^�8#8ˬ�jYZN��Y�D%���
�ѤD�b�5��=)�ET�C�$Ĵ��$�f�c�e���lQ5�4���o�iR�4��(��.K祄�$�Ʀ7NL�!:ô �ɡ9�ޚ���S�(�,�Q	Q��4)ç�@|��@0���'D4&+�T�P����h8���**W��4�q0{n���hR,+�>��R�M����X�n��&�wbcj���|��F�rڜ�r1��P���hYCn�˷���D���鐚�,��h`"0Mg{��?���PW���"8��L�*��c�S��gk��k�MP��x!�'�_�ޛm�W�O�ng��?�݃��>����c�tQ)>�a�ݳ�H_(�>������+e<8�}��b]V{�z��%�qq=۱��[X}	�[��/{|�������ӫ�Ë��N~J���{�]���M�SV̷�^^]�<��=�A�Q���zL��ו]Wٝ���u���[�9g���>��#�Ϯ�	y�����|���W�zss[�^G�Ϯ������N^������yqv��?�[�ۣ����r�π��Yw6��.�<h�����c�N�����ٵ��H=]�ճ��~����T8[ëc�mi�Q ]�xz���N�p 4�ɺQ�"�ҽs.��$)�;Eh�����f����-]�'��$u+�,D��ۇ}�5��f/��0��:�VgO����X|!��kƴ��B�8q� �6���.d��4��~�������>��D|"�'?���{I�md��@)d�#kL���B��v���z����Vod�8��U��dA�7L+�!b��y��(H����#W�ZQ�A���Y8:8,��
�8Y����|��I������o~c�4f���\zV3J�7�"XNq������,Hjd҉�8j�qhRNʆ��'j~��B���,5�RЬ+BS4��8��=0��#��,e�cJ��p�pF0��u�`�QVԐ��+T:ptDe��p��Q�eت7M���9����~�;�3t9"U��u1EMm����N7�?��C�{?��W-�3Θį}�k��>��������n��2��(!5L���(�$�vkH7�l�@�M���_��6�n��+!jTN��i��#48�Ѵ�^n|��%4[-���^�޼>ܯgUO�K�_��E�.�k��7��K�͟>������r��7n찋��}�J;:^�<����>���� n�����3,�)�d�+��7D-��M��H�N@j�����R�c�a�өI�^Ἴ���td>�<Dv	8��;ܘ��7���s<hB궺�J�8�.��=�@�HWHȓ�\�G������&��re�d[x���Djt�.5���dY`��"�����s�9:e4C���(����|�YlE����]*�P�QX��D0D)B,�oʊFo��B`[u��Cdx)�4�Vg���|L�6��biL9)!~�_��r-�Y���}�9?}m�44S?�484����$cJd�+s�@QU�u[!��KB�N�m�r����V*=V�-�O�e��|(S=  Kg{l�zB����\oz�	BȲ�uNM��m?n�"�e@�ڐK�����K$b��ՌA�%ᘶRM!|>&�%�����9�@� �9>}��;<8����d/�~R�ת�Jʴ�ɬ7�>q�ʹ"�����0q:pjl"����gYBp�Veh�W��3�Q�6ߴ��"����Hʀ�����-�a�C��z��QL���B��U���5��@\@�B@����aK��h%s��}���� ��[U�6�9����ܾ	q��I�VQ�>T���S��!�~RV�_�,�f�䗅f�m 'Y����Z���4��f +w�l7�ҙG3�E�X�@:���)'Z��eM�@��DC� ��s��Jd[GD�6��������"��A���:�s��<��M:;���!����~�Ƈ�A0SaM����o*1'e�d��/$�&�"i�!¯\)V-+�Y�|��i�A��N��c"
)d�mQR���7E��eM{�V�l���e©a��jq�H���hFuM�8g�Z�����d�)��� ��SM�	��i,��rc9U$Rb�@+�/�����@S"|��MN�����&��/�戶�����io�8��	�\�V�r�QjU\Ŷ���z%��==ĆS�������,�hB�a�����UdSㄛ6R�S�U�
�>j��T�)dK�pD�m
�-�(��eꡢ������E�yht�[�?�"�C��B���weS��k�*QbUb�5�p�Hhz\���"pp�F~)�4c����ו6�l]Y��&ZUǯN���J8~���O�#X��1�_��R ~ҫ�4����Ux��s��1�)h�r}f�8|d�XPu�\N���c ��`���&�r&G���~ \�j���V���C�RؤXSYvC(Xz�F�s�5|
:w���*��O��-��:r�Z�Su��7�ǧ�Yc=�P�*��z6m���i�D�y�����h@�D�,�*��Ii	���q p���SVQ���rKB������o�{A,A4�*�_b�z��1�D����JC��`
M���[|]/>+�TwJ�+;�@�BB����`����+������
wM�Z��-���������b������\���U�*G�ȹcwzᓗ&����!9ܯ����f�>���#�����W�J��2�g:}��}ϭ���Swo_^_^�<\]^�E�7���=\����~V�O�.>�ݝ�Ӹ},rۮ�/G��3�Q]�X}Ztu�s��u�r-��L���k����{_����^����ո���ʗ��_����W��xu~��q���[�>*s}�V����[���������۷np��i>���T�{�6w�Ʀ�����9��N�.d��׬]T�]�G�ӳ�ib�==�I�w�]��0�u���[qlw��a�=PHV
hΤ�{T>��$�������	��*�V���n�Û����w��x3�p&��֢=��c���H�h�c�Η��و���u^.eEY�ނ���zJ�����L�Bz��%
Yo�gwd�j���=q{�IJ3,�|���z����U�,� B��|N�c�b�fNQd�c��+�����^U�t~4�����7��S�"C����#��j��9�T
&e�~&��/~ᆓ�اf�M�&Y(+�&+��\�w�M�u"��Z�����XS'D������!qS)����(ڠ�%R��tf$R�!��/�,S�T��,��tGZ-�N�D��IK����#�����"+�j�jO���>�1b���"#���u51C8��ʥ�8�74�2�)��3�t�o��Цc*Q���i�m��sײ�u���O�S��Yh�-x����.��ߴ���:۵l_H�>�Y�����:Y�h�i֥&�hBX>�`Ѧ�Q��8v
���������w�K����GF�?;9���v����k��W��%��z�E�p����\���Z�oB��"'����7�gy}=�ﾩ%h\��䯫��p��i	���lc[�S��R�8�k��qg��7R�?�,�T�ct�\���8LZuɐS���S�$�u�� #Ht��vz��m�=��t��Tq��ǩ��B�M��׀��vO]m�E'M�]�6>���^�����ni�V�M_{�K�YԠf	�g�>�b��z��5"���J���'n�iJOS:�a�O'B��"k!|Q�P�)1�@j	n��j���ٮPt�6�*>�D��95R8��,B=tq��3L���,M�Y����t�ȩm�Qu�p��D[ʩU8����g8�G������!dE)t��m�_�D;!+*�����A0���.�&]=��q�ܿTя���ˡt?x��jS����׿��G�y�U��ʣ��}��>��MG�^<���q4�Wݔ�_�MYS�(G��S4~8��
�@n{E[cR��
A�4�!+Tz!{�*V���eO�O>�)A�G�K�ni���)Q��Q-Q>fY[dM�lq��\EYۺ�rґ�c��#�}��J�vj8@R@�.�~�>k���W?DmS���ګ�,�g���V�o��7YȦBvCȔ5n���L%��O>|LS��t.b����I�*VH���k��dFL�tjh���(�*!t<�/�����Hg��Ȣ82����dD ���hdE!zH���\�t��`Nb���l���Ɋ����ml����"#���2M��)ʡ��1�54�)��q��T��˭\uY)��J�����EA��n�hY�Yi�:����P.ݱ9�9r��iz���b\��1�z�)᢬�m�����)@��(|�9�����)�cծ��F��(�'�MqXxg�� �T�O�NL~����n �@C��/�/*Ѵ��U��%xkrp"W��I15�������J�Hd8�k����X>A�j9$���IC��g��ji�cp�B��b&R�L8Y��1J��m>�uU"�r�LͰ�&�Lģ�� �B:�B� 4�@!�^k��"Ǘ+�Z:F4Sӥ��:��Ș�b��O'���Ŷ(�PCV�T��&W� �l��B��72$�,<eQ��F�|��)7>�3
����s���N'�pR֛ZSEn+�(T-H�B�rgE�1{h  <&���S-X'�FG��0M�mᐹd���Z����DmhO��UdL:Y��O����)��;!h=Tٖ�9;P{5ϗ.� �X�n'J�,N�x�pʢ�aLHK����J�XR���i���e�Z��OE!���K?��ҍ8D��I����D��rLq��Y)&�C��r��h��(�OPt~4C8��-gp��yV3pmMb��3B�ps� �5��!1��p8�@3����rD9��pJ
�E��iT���T�g�:��i�ٞ�r\��lj-s�lǺ(��O� Dǁ��+�o(�Θ�#�
M�c9]>�R�F�"��p��l�^H�U�r�p>q�_V��(�������;����{�t����~�Q3��z�Y�n����g�����>������-��t��>*w�ux���s�s}��gX������8\��y�����ɝ��^\�_N?�)�3_){�/gj���NGj���s����~��<���ջ��=l�\��b{���������?���>��p���;?ٝ�W���+��K/_]�~v{����vr{��}�����w���Ý�ýޯ{�k�^;5��y����N5v�}��AZϟ�][�F���5e��:�+�	�.�ui�^���b�{&����t�L��#ꖉ������ng�?:E8������sWE}�)�/G�cJ9����F?mrHI�C�O�S�(����1Q_���w�+��V�tJa�F)�Ƈ�a�i�P�(K'h�p�� ���4���>��}�l���]
�&��6-e|��,�kʁPKĴ�B��Y��!�L����m��u����M�I���&�D�!��"��i4��@�D��Շ�=�MtL���#���p�5�к ����R�19�)���'dJ����ס�&���1�,M�����v��<�z�5��6q���!�D�b�8u)m�rmE|��U���/�����(��?ܘ��L=��
�=n޺H��%�4^p�>�ΰFR�BjUA�8m;ߨ�("W�U��g-Qh<#>t��t;�F�e�C��Y��{0������.���ıԮ4D~HQXrM`]��)��)�����"�H��7���E��������s�w�����5^D�2�����0ן��8��?������ų�y��Ío}����{w���W|�����|	��p�z�+�诫�~I��~��/L��eخٶ	��.�ׇ�Vt�o��R�i3�6D��P��������%
Y� ��$(�@�5���m�\4��x�'���d	bM�P�8/9NR������\L|>�S�1�6ШQ�P׌�YMȔ�rf�p��!�W�TE
@�<�K�
8YSL=�d�{N�u� ��\nUt� jX��ݖ�b�_�Vрz��ȭ�(#�[f�rm��OC�Potj�1��8m2��u�%M�ݫP�h� a��(��3}ڇ8�[��9B���O��'�S����x�|�����P���$�)�d�� 5C�\�(G]da����Z)kx
�B���v��RH��@��ܙ�'��tR� Y`u���ǈP���7��~�Q�J�}�ߴ�C�@L�?��j=(J���4�ڊjCE����^�Em]�B�h�����"h,)���|ӱ���ᔎ�	,�f��Run�,\�5:Z���ńs ���@H~���IY��b*Iǆ��~U��R��Lt��)����N��!��L�8Mg!@Rp�:!~��op)RT��Aߴ&�*!�ݐh��Ƈ�ҳ")�#%j����as
m�}�@���c������g��7E�Ɇ�C�%d �p�p��d�
M�EME���J�>ʣ#�gg?Ӈ�r�
�4�J�Bz*]�Q�lN���s��hUZ5f rȴ:U���*�Y�9 �jq�Pe%rt�QQt����C���k2Y$�
�m����&@8�o5V"�G�U���\:[c�|!�8�ƀ)��Ԧ1�;�F6RHJ�Z/�J�+j,D��	I�ބ�Pϓ��ZB�䳺���rk�r��	��	��cB"�� ��f���
�+��i*��R��#�S31����WSL�M��2��p��X�@�~*$7MQ���@��Bu����D�N\V�*���k�,SY��8D0�O4��3=vj2�E	*�Ɣ��#�Z��zp��
A�p*d*���D�I����Q?�a��N�&}�t���@�b���ޙ�ZR"@8���J�T�C�SN��3�е+�Z85	DK�5 q8�T��;mpF�f�x�N��i�,�A9����4��Z�S�m�^?�C�vC�C�m�j	MK��9�e�]B�Hn6m���\]��>Ghj.��jɅ���_
��Ư7���"�-%�9���N)��*���j��L-��[]�|��kCc�4��v>|�Ќ�*���L_��)Z:Z��Ӕ/�EF�B<^Vdv��S�Z2X������Z}]��4�Y�D&+�Z����2d4~��E*٩;��4m3    IDAT�xD�Lp�\
�(��&�%�
Rk���n�r$6L�ę�L�����t�#�����d��(f;�9���?�b�1YU$v����o���G�����d+�f�sf-�*�� ��G'@�Z`>S�T�R��K\�{Kȅ� ,ѭ���k^�R8����,ʑ��AVe�fd�̇���YP�)�^���������>��n@�Vإ�zv�����֭��Qݯ����{���?ko��k]���My�>���(�C�;i�i��:�<��5�.��=��;���:�_���_��_�����Yro��\���+7�\#���ږǯ�}����To]g)k<�������_/�pv�����~~����K_~y�Z���y8�9W�/����kp��?���γ���ѽ��ps�߭�+�=x]88�:�xv���3��~E���3��>Fc�o;-E���k�t�\YN�;3��.�kj%v�?�e]�ȩ!pB�3���C���>Din�zm&e�ƿ�ۿu�ܽs��o��]y�� �!O��� �6�K��w���z��C��=LMj��w��}rF�{tn�T��"=f���eE�-�4)�D�6UN	��X�R�c��&Ё����$Հde��}�����k�\�Z�i��M�"��d9h�h|jM-d����)��B�-]n��"�@|��غ��ز��㺔��w���`;l�m�8ߛ��#AD@�@66�������J*��\)��9���#G��9׬*�֮��%B�D� rZQ���ƷWv/��8|"�:����'�PHg��k�z1���w/}�³��Kot�ɧy:	Rfj945�tR"ܱ�Sy|Lj�ۛ���SuE!t��ѿ�g��{�,q7D��t9�Ά�����\�����N�n��H?Ռꚱ@���F	�����N��n6���NM���y�H�f���O��_�k[�����4�Dp�m8AR�8d ��k��e!��1�(�aM�JOD��@��B9<Z���[Q�DJ�D=�U:2Z�t:�ж�펕;��)E��_���St�P&�� I:`u�����Ֆ�<r!'��B���n:�p��$����B@ӭ\u<Q�ߟ���<%��{�ݍ|��Vp�	���.�|��[��|��xt�x��u�ǻ��7?~���������7�^�o��a[�k������G�2��?�цVU�=!��o�U=C�,��Ĕ��QB�oZ�b�M�B��&�A��Rdy����=-3�:��w����&��M�A�,�09U��g(���)gU��4:9"iڨ����R�AL� k[3��׃(��O�M	�ei�*�&��(5Q&Q(M[`��J�A� ��-a��@�lE���Y;Т��ӟݠIʔ��z�bBD$B��Z4&d
���A8��D(ה8��M0*d����(��2�FY49-a6!��FUFG��eJ��"8`𪈪%��.d��N�^��z���ڴ@~״�M��6��UK�&� ��W�e�̕2E�,ė�7Y� �6�D)�Z/�S��*
�w�) jup�%!S�~Tbj�2��,��{J/Q.��zPp:ϚѼǈ�;��l��VQ���^{��h
�XZ�6���c֘(b��p>NjEcE!e�pJ�fTh6��-G'��[���%�#&N"|d�6 ��O���4�jÎ��p\;>¤w���V�u���puKI���v M�P�uuJb|mD�!��Z�)���?��?tf�2"��>�9�� �Rj)ݶ{�D!��1u��(1�S��'�hHK�Kd��[E~L��9F�r�4�K�d�"�qJ��i|u�2b�C�����c�CpF��̩�v>M�����*|(�%�#��L�'�T���Bz�"Bơ��i��ܺ�B,5Nm�I��C͔)�����(�q�liƜ@dS����Ɩ���0G���V"}�P׮�E���a���hx=�«�)+'�P�i ���BmX�i�V�P��k5BՍhF r=�B�h4��&~���nE�RK�=�1��r�=��!�@6u����T��T�_u�����,�<vȦLdS)�=6�B8�?��D[u;`��SA���d�M�|)�,NOw�� H�~Nk�Wޮ�ڜJC���3}��'+Ȩ�J�&�=,4)ʢ\E|{���S���8���4M�`lE���HƁ�Ɓr*W��)�i�(js�z�e�N~|�i:rM�1O	�Rίd�� 0%8��5���Z7B#<�t�L�r��?>���	U·�V�7���]	��.H!�
�9"B���m4�3J�s���B&�8C����J��|5Q��,RB	V!n����负^5x�LW[�%��|RF'��ff��ƌ�S7�*u���_
>��m+b��G&��I�X�)?�:	!ǨaL��@�r�v-"U����Ô��T��S�($*7�hFL'2'N��`r 9��\�Q(�)8��iu��f|���^= ���q:�� ������dh�����B+���4�z8ď|�A���X�,��I�EK��BX��Od��`���hĄ�d�b�޴�^��i�g�
�	� ����B��0�Y��F�Ʊ_�W�EK��E�uX�\����.�e��[)֢��4�3��	�D(�~+TX�~����TV��)7�q� �B~��\)�J�9�JdU��U^g�;�9�q
�K�}N�wk�g =@¿C|���c\��ta{|�5lR���;����{�ɼ�\���D��^�v|x:N���$��g[���I��������~}K�۞W>'�ޮur��ޤ���:��>���hU�i7V�����Zp8�_�?독��\Ȳ�N��7�O���+�5�����w�5�qX���<���g/|2������������o�;��>���տ�s���jf�ۦ��5�A�yqv8ܾ҂�rC��&�ƥ)��:+v�1�-E�t���Z��g�*wU�~X۾���}������}]g���>���έ&�N��r��V�,��������w����[ﴸ!JG�L]d��_��2�ޡrCH��@n�x����ٟ��w�d�u�h��M*�HV�Q�Q��jۨ������X�R�ӻd_�X2}{�K	�&D
�c��������������:÷	]5c�櫮�B�B�B�o:��rH�":)�b|�22)Y����oL��#��#��	|�����zVQ4�(ddr����J��;��Q�WH����ɟ��_��=g���%�����>�'gWM:}'�Y%���H��ُ�����߅�8f��'�B��ΰ����n�3����p���O?�8�|�թ� =.�#�zu�I�Z�ci�=UZ�N�{!p�4,��)�Υw�c�X�C�y���4�����\`�5R��A!j.�z��2M����g��1>���4�c
�K�C4U���98FE!F"	R�.��Bz����b8��Lg8�{�6������+�Q�Aɑ �ъm���bJ�@��9@�e%*FB
�_���d��
šY-4���&��b*Q����^Q�̷����k#�{qe��3��hyu�%��r���E��}��x���/r�v����O���?9���y�������[��=Z�-�I�'���iXW��aMZ��YԔg�� ��e�h,|�M�m)�D?G�ic�Q����a��)���h����Y���;�=b�����m^]k� �Z��J���Y�R�g
Y��z��CE��@���9�tpL�f:�Lc%0UԤZpc�b�g�)���[i`��LE�Y�\S4��j��h��k#�s�BSYv�,85�#�O`j8@!F��DNS)��V-�Ԉ��>�!E��JYH��BE��"S`�	9Kp�� ��@QU�5)ю�FQL
�Ӓ��e5,��0�R� {i�� ���A8�k�`&��Z�\;�� �\�(�B�Ҕ�j�Z���Gi�$ȗ.T�z��R��f�9F�|=��i�a�^M�HK�TO��F&�c��~���?�sQ�M"Ӄn��z���&KTW� -ΐ�X�M�|��z~<�¥ӑ���4�d8��3��$c�Zn�7��.�W�u��s������������N�!#?e��,
F ����c�t�5���XH���!�d�6RQ�p:�v[3m]@���+�������f$�����: ���³r�5l��iNY�6��;0^�SV��Ȭ���j!�A�|�h����i��5��I��Qj8�a���(���O�GT����P0M��mj���iմDc}2�I�V+j���):Y�����z�r'Z�4��XA�&�����>\b%��"�i'�!0Y�MO51�G�s�c*��*���m�Gk*k�DLO�+8>�K���-�Ԥ�3�L1��4ј}��M_"~:�����a1��UoJ!�r���!q��˚�����8U	�7�Ӕ�O������ȆS?���[]��1�ȟ���9�0ݪ��jK���JC(s��m4��(�i��M3��JT�&�Jvrq��L�Ӷ�1��3�)�B����32_c1�c" C��o4m��0���U�3QAc�%�#7mL�B�)TndR�^׫�R���@d�x+2�k�r#Д�cD����2>D:�vfF��)e�'~��U7�UXnL#<pz�F>P'�{
���^H)�E��FxL A�3%� �:KM�@��u�O��@#��ȩ���vYi&$�FAD��ǔ�%��T�%�� �Q�F���e�-�'�U��]�(��◂�?�O���`�/���Z̢�$�
�ړ�ߣ[��U��)����)��j�>����@�4	�hӺJҁ������n�d�l�hB�)v y1�����
h����HE˒��D9!�~,'��I1�1��+��1NYu�H�b�*�\�Hc�P��y�6���,)=*�U�*F�o�����Yu�:���B�TJ]�r؈GF`�����i{c=I1M�35"sD��1H����C�D(1��V�g8Y"��L��/�}��uu�D��1�O�t�u[��]�|jK0�V�A�>�t������O�1���7��qt�&N��R�)Y:5`�Uix�L�	uE
�b�|�O,�M���_��Sq{a�8t�s�5I7�6)�/�W�o~zSt=��x��;�1��{�����)ȓƢ���/�{��4��9G_���G�fw��o�}�n��S��9�n���j}��ڵ��m-֊-G��6��w�My}L��J��V�o�����p�{��M����������?|��/�����U�M�ͳ[+�?��o�v7w��_";�l���Y��-ۃ��X78�E�[���7���pp7�y��#���|z�jsl,D�(q�|83u�lEW��E�~ A5v��r���n�?�E{�у��:�T�q4���0S����7L0ݡ1�@[[���)��!�\&���~�3�B�9~o�x�����������A�{VЏ���CYԝ�D<�9�*-�;Z@�RԪ�ꌎ��-#���"�W�i@��;���-+JD"U0Y$���9�:�|�)�M࿟��,]�ӈ��LA
�iZ!���) Ӕ�@��z��� �t�
U���W��I��F�xZ����F�S����,j�.�70!��p�ܗ�uG���?w�\�+�*S�48�k�Ѫ�,�6��QH7� rr�%�,M��C:'�(�a�� wt��T�z���g��_����ՆPs3�*:oj��yv�!�ޖ��P�O��D��\QMVS�F���
j��$D���"�4#H����M�f˯�t"p �@��H������U��	���e�$Ym�v gDt���pcR�t$jؿ�02�R6�M@��ܻ�.4d�W�)-���k&����h��cBp>���m=pN����j#ԅ�e�8����_!c��N{���L�C���)M
^x<�xY���˛����8g7g���xq��:��z�
O���%J��勋��������_}�{�֛�;����L['>���U��ڦ�l�ӻ:a��[{ض�������E#��d�I��R�4��I�R�ᕳ�e�x�Enl������:R�����?��?E�P�*��4�ќ�u����(��!�`�4�>��Li����5��(K.)�Z��=`���i@nueq�h5fĔ��pf|�m�֞��z6����a*2�L�I����%��U �(q�x���gIQ���+g
ɭm ��Wb�R�NS�~" ϶�R	#S��e�(��j�рt��pR��V�qH!K�:Z���8�C�\���N!�ɭm�:��A�8�����+R�|Y�!�<(� �I^���.������@>�Z��@�#��Q�6��^yr��`�h��i�"�!���>��z���������M?��S?�q��՝��ыn������=�	�N�8����n���K�V[B����7#���?O��(���ȍ�D9�.e�,���~�����@���d!�[�1�4d�pf�F`U�|`�Sá � �8TFQ;/�a43u��S����έigե�'U	�)�k�����.��0�UK[�U��㼵�-���#��pl8
�������*m�o�Nxm4�eJ�����֪)'�rH�&�GV��Ls�@h?!��G��S�A�O��MEUI����m�4�:�1#K���sV���3�X���Ȥ�n*�Af�Ml�qD�9Ӑz@����T��୎�Vvh��7 ~����?���)c)C�T�N�DV��ɑ��j%�&�td�Yr8��X?�@��YY�D ����P�i#NE9cIM.f����A�)|B�9�x"��9��=��M(Ycs*�fHu!i6
1��/%��	r6��Dhj�Yc� =�J��M�0�-��]�ȍ�=�8��C(����X8NY��p��T�BUfl]�pSM�ʗr��g��%�#��3�ͩ.<0�qR�M�������c�Y�@���F�X���������S1)S4>��ڛ&�3�s�^z!���>���E%��	t�:��\Hi䥵�'J�Z�
��At�|��iuH��,�� ejE�!�X'1#l]�]b�RR��T3�c6��ZVQ�4-���T=�hj���E�#"+�V����(��ZHA�~�B��hLM'���QP���l�eI�6#���5l�!}�h �m% �L�4?���3|��TbKZ�g.�$��D�#�#چ��J��G(Z_�.�T<����I�rFmv!L�4����č8D8dg��8@j��+�~`�.��h�(�t�Fb,�,>G����E�+S0�g�;-	4�#�{h�� �=�1}#��j�ڍ�AHb�� 'GԘl=����q�$A8�(��	S�gT�z�M⽬�Ul��&X!�ЬE�B\�T�@�VK�Ѥ0�p���<�w.O�Ɣ�jyW�c������&�޼�^i4�� �����G@f�U�kF
�!�.ǧ#�_�\{��>��e� tcћ��g]��s�>��>����������[��������_�v�v�Fԣ��i[t�f}����a��ŭm��l����*�ڽ�8uu��ڗ����/߼��P����-X��߯;��,`m�:���gnd�|������ꊘ�3��>��Kq��ᣏ����o��Lo���/_�c������5�觶>:;����>���lϮ�Q3[�����v���٦y�~&9����ei�H��o�t�����f�@�K̇3�"ζ���vD����C05v8���m�v�)���D��wߔ��t�����%SR�3c
7��J�*��v�ÑN���X/�2�ړU����ƧP��5�!�t=S�u7C������Y�xS�F�|5:Y�# %��Fͽ+�O�,"	��r�>��9�Z���B�[N)��J>>�q�����u��ϲ��'�M���>d�z�$^���9E�\nQ�����ψ�h6\��7#� �����b�QSRq�.\!R�*�MD(��ɗNV.���YQ��C��ԅ�D�����!���3M�D Dh�HM9�~<QCL9��"��;���đn�f�u^oE8�t�b��jG!R5�O����Y�EMe%)���    IDATZƜ�����|"��k�T�Xu�ꖨ���K��E��D��&�wj��v���7{e�1 �ͩ�w��]l�k�A*�)���.�����AY7p�B���T"B���������1r{�5�ޖ�H���H4*�×��[��{��M-����}�3����K/������K_z�N�kC�?ٹ���^a��^��^]{)|<�����??<�:��1 /���6{�YW�|]=m��'A��ֈ�+Kku���c�_(pR �R3e�r�BN9��
���ܞn�Prq+���Ӻ^��>@�)�q���ՑED!��N�O�Jt`0k�EAcR���M�`]�z�S�Wѕ���G@)r������4vB�g�s<�(SpB������e������_KD��@2S�����V%2��uR!�L�5zRK�T9�(>\�Q	! S=�*���q�:S"�hD����b�AP�}��F��N�q��@��%>L�O�C
�5\��г$�ڈߊX	�
QNFA�h�b�yY��Y{]�Յ ��@�	�9^xt��X�Z!�$D�fD��>�3騔"TT-�ojT�Sn��D"Ą�{����������O�Oa=H��fJ�y�*���­��X����4���cd��ѭ>��|EYE�ȭ�Ќ��`���E��J��R'pS#�d�g4�؏�c���^Y�u�:�R�: �@1"j�1����@���= _�)Ǵ���/Ũ�J�)g.�&�J� ��J�9<�8�� �C��mbOO�҇�!���;C$܈o��JP6հ��thj��W	�^>FA"_4e�ji�%>��txL����p-q�5����>�T�r�fd1
�m�O�8���C�z�B�%��r�RJ'�8V.M�c���cR��S��Ko�E�bj]z��L�
�!`��J
�8,��-��\�ܹ�Z��h�Fg�ӵh)��9�FE�84��u;�R�9)D.Z�	�q��ZV!Ҏ�cmL���R��Y�)�M��4բ 7�	��P.ڮ��)G?p�LSbY���#���Gٲ� T��Ө��?��#���I���Ǚ��L�!�h��?;I�P�j�Z���E8m��(�E�V1�a��#-~c�p*�d@�,�gc�P�l�5(J*���B�H�KPT"�)�,dm��ֈϷ
f�)YS ������Ӹ�����˭
�녦%))��]�J,WHz�C�t;��|&%B�38Y��_5#G�/]�#+gE�$F�2�\S�,�K�/��?�H!>���uA��i�ܲ�nd��ܐ�A�8)�,�����F�Z�<F��$6k+�f��M�U�o�5��x���D�q\5׶��Q����)�e�Ɋ�R�
U�fN�_b`�i�a@"u��O�	I��H%��� Cf&��A`*d�7�"��i�h
D�Β���)�``�8B�"�RS~G����i,��c��0:��sQ�~�5Bj/5SQ���Cj�O��J2�i�|6:s����*$��ԭg�K�\#�(~�ݓ>x�-�i8�<��f��`�&D
��1�B�B��0��huU�8�]�.��i�4�[
Ӳp�GM��?!Ω�`��WnZ��qR�U'��f2��Ğ@J��C#ЃQ
kQR��|�
U�o�p�ߪT�X���� �|rH��8��$�'X3���$��z0�<A) �X�zRE:�pꇓ�D�l[|k���><�w���Z;7���[��\���t�I�c~��y鳗o���P^J�W��Ӟ�@��g&�O�?\��{��W����'<����N<����˳�W�������F��/^�m+���f�^<��ț��VlU��:W����;<n�}u�n5��������g���ˋ������~�����ώ_����������M^o��vy�_�az槶�����u�ק��f�Z/��ֻ@���z�\������f��.��nK�ڀ{z�
u��J�v�|8[��|M����cl��)U��ܛ�#�m�g~:�SS4�45�5Ƅ�e�^�!��Z{Q�|�t�&=Rd�p��]f�t�WG���GJ��p"h��j����� �Pc|Q�S>B��Í)GP�M
��D���%��@�U>�5�D����E0�'�!Ӕ���5M
3g��ën��ˍ�S���Ԯ���y�2S�={7Ŭ�1���h�v<"טA(>2g���C0S3u~<	c&"�\;#A!��~4�� gr1��P�i��>i���� ;od-h��QSR�J�j���K�et ���VǤ���oE�B���yY@L����|��I����ʊ���L%��=S��W�f�[�u�p(s�Z.GK����i���?��)Q�`���o�>B�ә�&=멁djT��b��6�^=LS`��?��֥�Q�JwQ�J��O�#�ؾ8^8�/���<��o}!���x�Ú��'��%������p�yq��b�k���_�q��xx�h��ӗ�@�^y|���������Ͼ������`�����_���=�N�=7�dF��H���BZ݊of9�+e�IN�l7������R��$�i�� S���U4�Hr[g9B��٥wVܰq�?��cW�M6�ߩr!�Կ��r���A�8�1+JJiEDUW�3�&�������RhZ&}�@�X)��gSR��J�QKi82P�pQ��B�d����mEk�E����p���pZW�Bt(�q��hdS\:��d�'q: �UW��fZHK0�s��(eҩ1Y��#�8���#s�,A�c�?�($�r���F�������!D��cNS)���q����R�5�s�j�ρ['�i:_-���AP��4!
]��R,j۰����t�YF�j�j�A�!5ѭDQd{��U��K��ҵ'H�Q���U���˿����~���d�.��~Ԡܶ|��'��Q���1�׆� ����F6�6Bg��LS�^'�����[��I�BKw+� 1j��=]�b-8�ൢvF�[���#�����CPz��P^U��D������ Z�\u�|L)��,���?�fz$��K7��9�u�d�BR�B���_��:���["D]{b�,+M4���qj8�~�H�D�E�_n��Gm�B��4YS���r�/*���FS�L�8��D3��mQ[���2"�'�N>KG
��X!��Ȗn�ֹ���"�gK����3~U�[i�1�S�h�J�4�BE���ďƑ^����̓�-���*�^H����W�Tp�8�5s*��0�n�(��Ǚ~TeS!�,��p�"��bQƩ"��%k G.�s��1Δ�,�Q��d�S2�XnC��9[��� �X A
��L)CXm��i��|g&5#�t>���=Gϯ�Ԛ
������h��4~�Fў�� ��_����I	t0�^�O�!d|�,A)����h���t������Md����ΰ)�Q�Rp�Yl��C�� A������p��X Y~!SY��L�#��zƱ��Z��PK������p>p�A� p�:�Dd8Ј�f�1"�U*��+ڏLvi*�d�E����\�c):�Q����g�V1LSR:ACfE�J�����
��n��� ��G=���u���<��F�Q��Z�(2�iڊ����(�)G��F�ǘZ*$��єq����WH\��t�8�Wq�y:e9�󛆐�Ԁ��i;��A$fK���\�18���Mc��G�%�Y?�FQ��_BVQ��h���r�O��CJ�@P:�=��)�R��O��S0��h�L('����N�H?�2]���.G)�:�z�'�6�	r�R��-�43�A�$�1�0:9�۪�un����h	V"�R0�N��jĉT0Jg��q�C�h~f����G
���`:=���%��8F��3��y),�{ĪT���1EM��(���ג(��"��'~Yq�uu
i��O�'!N/����9������4P!��F��N3���X���p�,R��[�Z��=t6���
�-Е�g����y��n��g��Z����v{�������won���~�ݯ�P)v�{��� e����Z�%����:WBF��Z
���%����+o;�9>��������m�Y��o�ݾeo}�^�Լ�]k7�/���ͳK�Y}�T]�Ն�\S\[�~�=�ͯ����(����a��8�~�q��ߞ��=Ϳy�pxx�?�{��}]��7ܾ{��h��@����
y�#�1�`Q�}�k�po-V����-�.P[m�A �#�َA�p�v�Хı�Λ�ĕ+Q
���2&_i�Mz�!�΀)PV|�3���c@���h�r�x��\.�(���Pg[A�.6�s0k�(K���ȊP	S�1BY!�gL(jզ��,�Ó�E)�� nJA(ҢD!��M�&��h����q!Y���!}N4c��*���E��2�Q�NR+:!��mR(�ڊX�����b�i��8R�j��_�����2~|ǃc,ST'l�:�̔՘�,%Z�&��DI!G�]�
�B��Kt��)��t�D gh9ĥ;��1Z���u�Ճ�&HA'K���WTJ4c�"���Ɩb
�^W�#�9��#�!��j�H��T�ϤA��T�=5�E���+Nd=p<6)�:�1�����s8v���@걼s�J���*Pt��!��<�p��7�g���4`2��;�V�lZ�+��8RD�mzEi2�B�
y��mW�n�q���ʁ�{����GB����n>�Fg���W7珗�k��Vp���߾y��p�p�o<������זQ�z���'�/���^�=^_��7���W?��w<\�ۣy�F����������#����������Q����z;�@�������[���×��8-���j�Q����i�c���g���Lo�8΃��$(�Ov��"Zۜ��`5}�E�9��WQ!!�V����!�� ���2������5C΀��"���Zk���+��r�ᮩ�����6N�QB��B|HQYp >�Ȣn�~D��d4�
:��m�Ƙ��!1�r�0>ӕ�	b���6�Fˁ�j�R���h|�̊d뜾͉�r�-��#��C���aU7��p��q�ni �O��[Y
I�$G:ʹ���~�h!E9@����]HO���j�&ey�����=�,�t,.9e��h��j�#�ej� L��d�g,J`�+��4��aMYz�eȘF��|�;d)h�������Q�ȇ`��g)���jc����cZ�p!�,Ĉ	鏐��l/�@ʖF���,�[����E��Z5ʭ���!ь����՗�<���6U*��0�X�����ǡ�n�r!L�@MS�,��B�p#��@���U��WL��ɏ WW4K��`*D�T�U��U��ʹ4>�r9L��xY	B�D�N�8%�t�V��=x"�Dj ~�Rj~8��m;C$���وi$bdr���Nj ��0}F�9�R��Ɨ躠%8�BF�������d!8]���5
=��	�ӴD�ܔ#�ͩ��D4S����1���L�B�[	L�
r�Hᜂ8,N��^~�G#�A����̐9��A���̏��R3%�d�̺*Q�%��q�)F�0����r0�5���c�9B��5D�3��NR3�R��,�)�a�S��D��t�F+QJW�{�����\���v�� �1�\�1S�#W���zh�H�>'].�u� +�f�l�B|�\ms���Y]�=]��\T
$���,)S����2��)�^�DK¡l�!|�,���_���l������~�$�C��S2�3��C�
>�S#�fL��"�����Ki��uRc���k;Q��t$�V"�_��2~M#�k�H�8�|V:)x�jA��:�����DY�(�O�|L&�_HJU�j��-�+2�s{^�t�%�p#�ŦO���h�J#��	/��Vc�S��ƚ4��dq:l�Vh��� �L�F9E�4��5�?�H<Y�,�,���k��J��81фL�:�"���hY�8IUň� ���%�mѱڃ��_��!#p ���Ls6�Ӄ���c��i�:Pz!N�uqj��d�3q�Q�?��!|ۘ�(X]=�?�w�SH?H����	v9�7���F��٬�tF��u��N$�e�g!f�=�"|�)��h�4ֆl����i-ơI��i�"c�Ap��h8�o�Q{��0�ֈ ��ѓ�_[����ȍ LJ��Wk
QG�n*d�=%>))����0�ů�4�)H�����U�T[����Fi�.Q��)L��h��U�츻�����չ��vxد/�s'�ߧܾ���u��u}
3[���n�'��{|���W/=�\���R��޾��wA�����}ԣ�G�%���B}�r��՛�[�G��}�뻫K�>|u�z{o�q�ov^��>iy}��e}K��ݶ����X�ԣ/�%�=P|����zu'�b1���_"�]���W/�����~h�!���Wj��|x����ŵ��=w}n�n��ǋ;A=zC��o�~������}���<��O��@o���A��G'a�HX����Dic-t{�s�E;����Ģ!�K��m�N&���nVJ��.�����g�@g�ȏә�.$�pF�4�A�VāP�"��S0��l������sB
@��PF�~��)�Os���p�mv�rd9BB���=x��DQ]y�e��/�>[�D
�e�	�VNՍ@6��0XH�=iE��NW�9#�4���L�Ԍi-a��\�]%U'�*���D8$��~� 2��
f�U��&
��W���aH3�U-#d�ouM���`��ӄ�2!T�@
�uE_��롅ǧ��Ϻjj������+A�O���q�& �c���U=h/A4)�4Ƒ��P�&��7�[z��B�SEmpDY�s�T�ߨ>�?��[V�X��V�15}2QFD�^�X�u��-*�A�f�Y;;�;p�-`���Y�O�5�L�yB�]cZ�Z��3����D؂k��8�8j�jG�`ǘ���j}�5oˎ�����������]_��{yu���Ɵn����c����w��}��z��~�]�O�|X�=Ig����̫������7��ÿ��������돯^>>����y�tC��賡
����z�ӡEYH�s�O�H{BB(�c����v�,Q�1_T-d�'�O����� G3�Z�L�]-ˁp�m;����pL̟����3�Q�+d���$�ӑ�u4�F�u��r!�S馵]��(��-�>�qŌC�WQ�ꐚ$���qjI?��BDXP�(��f��%X�4�$�4Hjj�=�i�h�F��4�r���}����U���I�I�1Rt$�"ȵ(�1�Jë�5�� �b�^V��b�Z�tNb�YQ�F/<�*X��9T��H�.��"�|䪠1���������� �b"+�kd�@�E0;BFI��sr��Έsz|q�\�x�FV��
y~��g>t�i��d������h��]�{��F�L�Υ�����������@A�e֭���D1��D���o��F4����&
geqD���r�����h4�1�u�\�X��Η2R����|����Ϙ��A�4�r�iR�4�77k?;K����=)v���B��H!W%}Q>��G��)Z*RF0BpH1|d#BVb�ԃ��� �Rp&]���F���8M�d-��FLK.�H!�hZWh���t�8E��252L>�Nt��)A���i(j��F���<��R����p\������^�	QP�=��9:B��$p�v;�r뤱N�L'��Cd�) �4ORϤ2Q��R��Jg��
�1��_�,(t�9����3�N�Kb3���A.����� �d�7��-|:��r�ʕ��)����\cF�+^?Rz�Uq4cR�	��A�����9,)8Á��e�����Җ�.�)bJ�S�,8��j7��8�����zqBrp8E�5R
�l����;K�1��:K��d�D�c�4��U��	�J�b�����O!S>�?͘V1�Xzi*    IDAT����_V=�ES�Új��҉�O~�j凇Ĭ8�!�>R	SY�G%S�._:����Y� �
�Si���LbD�	�t�t�F�5���q�~~��R���x�����`�$��QX5N����� sh�rMFP]��{e�!P��
m煦���q�4�keE�T��e�7#���I3�q���v8�{{^�p�g��u��=5aB��_���g��FxcV�h
������0���Y�3V�N�i#D#g-HӔS��B]��T�'vo�����ޔ��s �dh��9t�h�s��Z��N{!H+��L�K�i�M���I�N�j�	>_Wq -'LV�����r˪�r���O�R�=S�F�i�Ŷ.Q!|c4�Fv|N�8F6U&=~S"RЦ.g@��Lj4]~�/]�B���(Ph���D8����O��/��u-du��]������r�A.��R臠��|�~Z�:��r��I|�Z�QH�u�W�}@��VA�� ����<K�)H��2�6Gz����!�,#$�)ZN�t�$RHQSYd�\U�_�]����L��$!�:YQ~�A'F�MeAH�d�g��X���=n/�V糎��3n��������Fr��q�rwv����u��u�|1�����l�s$���ý_����}\�K�����^�O��Y��U֝?o��~*8;�����w�W�P睿�����A��gw��Es{3�1�W�nh:���/�u��������	�s�E��pO�r���Z~���g5��n����?�.�V{�=^�W/v����{�1�n蹿iv�߮�����˫=������}V�Gl�7�rA�}�Y�Q�]Μ�.��j��>��V���a�.\Q`Y[|�YG��(*�iYWp;	� ��E|��6���5V��t�!%ԡ�Bp~8B�J`r�©h�v��&��9�Ȧ���@Y-�&߈�$�aC(�\]UW�7�[W6D��J�*+�������fZ�y��B�stb4�L�i�n�]�9-�$U�B=upfӄ���v���i�\L����d��3�XW��o���,�)Xo�� k eY����.�%�2�,�YB3�TG3����
��!8�!p|�,:"|�k��(��15�G�O�z���ZD	�3YD�yQ��eD`���3��j	R?h��Y)�7�B����zz���3GĘUZ�#jd� �k
t9�F���.1&'���P��Wy�A~�ְ%�L"�nzc�{��n������H2��(�2 nt�,��6kIF�M����6�!�E��J�6�cԨ�|�C��5�?Q�7�u��7_�~��������\�-�;�����~��$vؿ����������r�����H��9Vsw����񃫛?�<zg֋�n�c"_v�%���7�n/���^o���K�S�U�«��<���Ǉ:[�/�wu���v*����_��]]cK��v�ϱ�m�hV4��F3��#DN<N8��?4��c�%V�1]�l�5VNor��(�n좷R��eA��ZȢrU7:K�Ðj�(8_�5��|)nO+Fm0�5)L�FVT"$ǔl`{"DVHiY�rM�L��c�C��Xl���a�ub��~��JK��*�Ө����d9RH4B=�c4E�RVk����R����g)L��/�F�p f���C�f��8!�(s��Bq��Lls���h�|8����Y}��8�d;c�jp�s�T�3j�VK�3��B}�!��&.E��L��L:M`�8�8�dSִ�G뱉�z��s��p��*��BZ�&��,��M��~'5���r��(�f��y����QY�NYQ8�CG(�H\Vd��b�6>�8�%�ǉ,�c45f�G6MMW��#�m�+������Ñ�l�V?�~�y��UL��۞��3Vm�m�3U_�
���s�n����8��y�σ���p���w���u\g��/��yi9�����Y���O��F5wq�N3�V�%��%���K�,��#��ʦ�d��F"F�c
ɚ2 C3z�����p-��8�z���[�*b�Z4C��Kb��r�������_�Uc3]i��*�Z��V�f�L���0>��!���Z�?5�.+&+��`��FG9>�Ќ8��u��z+�_WDD�i���Xʉ��R��g�����T�`4%8���C!�B5V?�p ��b'KO�bu#UF�"���$&�HPt|����m�V
��|x�l2)�E���6����.��7��*LY�8��b�q�L� ���􀉚�I0�F��d�W�X]c�I�m#�i�~ t��VO������8F-Hu+W�8ڮ7�B(J����Y���w!�|����.�rąj�ʂ�[u�\S�R����nZ�E�	b�Ʃ'�B�ב����+�+᰺�@DM�qm��Ȫ�P��7 Ĕ�✖��:��Y��a4��hS4YF���]B���pD{�S�	DH�Q�B-d8�o��ѶR�mSj����|��`LY��E�[]mI+���
IIj*�5�XiY�C�#��zar;�r*ǆC��)��R�$e��S���+�����+c)��b*��_Q)U�
�Y%8-����$U]R&J�H���Mq��*��&�5�J!�U O�y J���_|�G��'r
�dQ�|!�kC�jE�1;���-p�I�/w��!m��	<U!�UN�Z��SA��Q.�u����U"˨ A@��h�F��Ө�Դ!>�����PE!��a��7�~�Z�c���8"�� dF�z�t�d�`���&#h�)2�l!��O�J��jF>&s:T+><2M���5i̒E.�2\V�ƺES���4�Z*kU}^Z��"d��iJߔ�1�V:B�>�8:B��i6��@�Ư7�r��sp?Q1�vY� ~"F�8�
�1�B�4�.�<o�ժ�tY��T�* b�Q(�����?S��rJ7ɧ���B�m�>�P�+��k��x��ǋ���m�����7������\��$�C��d��ɞ��o�>c����tp8���:����%��`��K�r�-Mߢ������{qs���{�[�����l~��*|�C|�G�8}��_}x�{�V�3,�����o�n\���s��>$�ޒu-��������.�}u}�컻�/��z�������H����W�E�ϻ��+�O^�ؽz}���j�������[=1�9����6}S^n.�g���Yo{�Zƫ�\;U�|���
��G6���l�ݔ��⅌�_��++����\	-�*��c�F�#�T��L9,G.2?�c9=�VVS��4My�\BE�)�cf���u%�!��X.d���VeQc�@�T)�(<���gZ�gB�	1���Z�H)�0�a ?�h"�NJ=7Ξ�d��C�TE8�����!U�.��B��E�T�hY��|8�*F�s�(�d�~L5�gYSdQ�����9%��K�0Y�]��!ͺ�U��Ѷ���)��LW1�c��D��*F�����AR@K\!��3~P���"'�flZ�چc����P@��[)�p83�R!|V���േ��OsKZ�n�K���������d$�Zsdq�F���	�I	���I����#�fw��쥊l�������l:g=`���VO&-Q8��R?�Jﶫ!�ʍA���uB(�a�U:�R�p�D��)+���k�o@_MZ�W�1�$�3�_���w��s&�����{��g��;������Y/y��b�zyv�Kg��?����>���������k����q�����x�;}�����V�Uԑ���g~ ���������_9yk�'V�́���o�-��ub�v#��l�گ�'JL�7�Q�Ԟ4�,��k���6m����+
ɉPTQ��w�Wnu������:Fd�:���6��Eд�����a���U�d����iQ�w�Ƙ���.��U��s �ǤCl�Pգ)����# � -6���I-2e&EX���唆s�T�>p�ڐe�l
1QE�(đU'��.V%��2�SK�(���3�0u�i�h7��3J��@c=� '}4LƷ	��E�ШD�)_n
S �DS�9��O(ZK4�c憖��i��!�T��
U%�1%��E>�P�7�j>2��X��/�Q�����_?����áF�̿�����/٧�]/!O�R\ǔ���o��%䓝��"�ˆ;���#�'X�}������$+W�p|�J#�M�!ڨ��j/dh9�6m]��G�גЩ_z�v� h�8R��G�>@\#;i۝�\��ͤ�J��?�K�ky��S/~�;�����k�T\���ݭ��q����
�y�ŋ���ֿ��[��~����W�>����w/�?�ɿ������¶�~��_���kCK���0�i�ǵhjQ�u�/�nt�L�������4�HUB3��VW�O�p;i�L�R�4�e;�AF(��� �� Ƙ|��[���@�| f�@Ӳr���7�U�����$�i{�Ԍ�!X�����9�:IM!�q�+�T	f�jF�RL�OgȥWX:G��Ia�Z��ۙ-���4)H4�On����� a�-A�Ѵ�&K]���!cVwX�M	:�ӡl��ǯ\��[�ӭI~K�P颦uX���Ux{z	�cZo�nbD�ק�rH4E9��8)sB���B:ԹP�N���O��9p�Q.�ɡ��1�L���Y�ɪ
0��Rʊ\�|�ɪm��rj`�R e�wiL)��5�תD6�SQ3�E�Y�|�5#1����Y��+`���Z�����ć �3����hpv�~ �k��7V]:�CXm���&^
�3|QM�eJE0-��5E��
�-�������yY��c!����d��3���F��������Z�81q���5�'�d#����Cd����M+�4�ԭ�:�S��$���R!������稲$6>�IH:8Rҡ`*TV]UȈS��1*���|KJ�����:�̯Vm��R�ҥ�\�Mn�*�W"�яgBq�jɔ���$�ͫ��(�6�r�'��Rdې��*��r[�i�Cl&$�Ul���~δ-��ɺ�&ٲ��9DNw,�@JlJ�@�d&k}g=�Lf�z��jcS�HJ P�9����+9`�|/_���>'"n��8�HH]񑫒�GM�Z��B�*��[Jx̐Y)gdea��2���?���N���5d
��=Z��S.�,#|� ��"D\��*�!e���j���BXuc����,�2!d��B��>��n��v��D�*Rcz�K)1G
|�9h@�B��!>��XQ|ј@��Nz �	�nd�b����L�-�l/�~���҄#k�T��)�'�ЀC@�v�6�D�aS������BX'*�(SˡO0)�)'e�V3:!��8sXq�U[�X�)��A
G3�+$W�F���>�Ƕ>��կ~�|c�^�9�X��kt��1�� �5D�B[���rݒ��X�	��,�C·��}4�~��yp�p�6�������Ɂ�̺���޶n����Z����ჯ���m��vc[��D��������>��	�n}���HNNO��\�4_HsnE�%��U؋�E���}Fk�e��c�����)����Nw��%͛�_~���_�}���a����]�4u��7?~}�ϗ]i��d�.���v��X)gw'���(�F���7�t�殫�V�m�ڛ�th���Y�o��v>@���Ĺ$���-K�jn3M
��1��Px#�l%dA�@���d;��{~N�Zȣ\�9��Mm����y%�������t�#TH�/+��+�&�g�p�G
��8�A,A�_�t`%2|c���c��I_���t�i[�gD0�bJ����m�)Z��L�I1&�G�'bl۩�PR�j:�|"���IRhE�l_D�����1��4<|ߩU"���Ɨ�!�H�E3e�m~��b�0�!j+�e���B�2�3L�K�e0���a�L�>2��2�� ԧ���Ϟ`�>^:�>�b���=i��'�]j{9�S�礉,�L#��ǝ�r�"Й�2Ρ,'Y��8,�3�Q���Xi��d|�c����}��������_ s<V��g����u�'S��>�2���c�^.Y��-�*ײ�G֢���K�@&��W����ϋ�/ׯ'ڨu�z�ٝ����G����w)��V�M����ts�E�����m
b�-O�';5���yw�����K����'�����?z������������W���^��v��oU���\�XW0��[wT�Vj�F�J���˴�!��爖�4�#MA��4��������~�)DYȖR`W�=���!F�/=VEM9W>�7�.�V��R|h�l�z��M�f�����xk�w
����ƀ�j�t媂��s��D+j�e��J�O3\���1�N�ϢAD��+��$F3�h�ZB=�(��z���v(�q���ﰮЀ5�c��t�P颔]�[禑�5���1�7"�+a��ON�(DǓè!h�(�_�t�`�Jaj9F��t�v�H���N�
��Ɩ�D�L�	�3��� ����GfMe�-���GC�mSLS0�bDұW6��'V��j���
�Ҍ�A:%RP�r8B�?j�So�@>C��%��=s2d�}��g4��o��2=l���b��5f	8��|�K[Z�u���N�MG3Á�0&����������c��
q�|jFQ����wȥ�![�D�k~6�V[�]M�_�QS4�qk�mE���=�o�*�]�ݭWTez���9~�؝�ν+��Oml��_���{?��> O��Gg^�O������������7Nε���uz����E�� lQ¨�Nf����F:d��Α�=��*�ȫ��LbJ١�@��zjqL�ďf�I�n04Y�����OAј���Bs2h��i�1�nӘJa����_?�ڃC����8
��� 3m[����|#���'���S~+Bȱ?�=�	�JHq�A�}�
�2吁���)C0�׹f0����p&���l�Ʌ�+dd
�J���8p�*� ���)���>��)�>�z��h�c�5#ى-1��M��FY��>?� ��+�q�W�M�Z�ә#�N ��ԨSj|d��e�X��B�������M�)f�FӖS�!�2
�����@*�#8����t�,N˧�o��L�0k�?�[]���,�z�|�U�z�8�)+N՗��/b��P�T"����p��P:��Rc�5�1���8!�ZE���'��L���v)�6Rk����1�D��g$�_��h!�>���7�)�!��r�qj��SW|Hj�m���c=�RN�8�����4�1S �9�?'��m�lh��~#~M�E3~6��G'����o�7�c*ڒ��cj/�v�)eN��[�Z������)�ԓ�?����M�|&kv^z"F6Lj���s�M�U�.�M�X�Z�'8{[�Ȕ�����ˢ/�B�t���J_U�n��%N����M�AG�8F4��V�o	�o�u
��w��̒��8p`:��Q���o�B�L&W{R �V�T���U�'Yc� ��z���$2���4Չ�)�%#&"D�s(�i��嚶.>BPzʍ��B4�CcT��S����ES�^8B�;3�O�R�g��~L��mf�;��1}�^�L�D:�����4>���[�b���V�|"FL�*���PV�q���A|j�3ibN�V�ӆ��×h���]6�#W
>��3�!b
�܈Y]�5�t�~~���}��E�
y��I_cU����MϢ5̩[QV�Q�F�N�{�_���}x�8��-s�5� 9h��vw��>�	�}rwY_X\Wu�t6����t!ŷqt�:9^��k���]�t��UC� ��W׷;v>�]��Lq�;~Bs���]t7#Lwg~����eœ�v}}q�Z�;���G�p!q������5�lXkw߽u��u�8M|�c 9�n��.mk��ѵ�GH}����ٱ�<9;�=?��W��
=x8{��= ߾:���+��|�敷�w���K,۳ĺ���Η2��ܵ�����ɝ�nGm[�"s�����ѝ3����.����    IDATS��oi��=���c:8�X
�,?��жM{>���������X��"N�Z�I��[�i�Q'1K�f[ꐲh�[�zN6��s`{\���4eD,߈�|�Q2�_Q)����-�O͘�a= `F�ɏi��F�D�)4�E�#w�^�K���L�#��E��2NՑSÄ�� �k^zH|���\��s�E|;����?���7�G�8��83\�,�RC�-ć3�D�M�U�FMrؖ����ʕ^n��E���0�?�%���-���:�zN$�}Ӭ�*�m��H����r֛_Vc8G�&KJ'�h�l���)�MN�����n��|~i��zxL���$�}�i��k���� ���������]��ɶ�����o��y?������$��>�5%D�Cԥ,Z*��(�-sm�.T�A��:N?�@�Zbʕe��:��1�0Ԁ������z9ٝ�[�?���??������>}�����õ�?�����s���4�t|��v��6�ߟ�>y���'��޼=9?���5�}�^����gGop����o>�<\�N�������oϾ����Y�k}[���M:p鯍jrZ��9��R���M�(��7����#�h6�=䣥P�3���K��s��鞄�~����N����k�����T9F^���6�Ot��>崧b'�Њv܍4g!B��-��6�)N�B��6˄T˶`�zV��7Ji
/W|��c�8|K�,˔&�q�h=��Q�)��-�� pY�p��8-J_��[B��"���S#�L]��?e�j��p#f�}GH���٪!JC��CAKu5S)Ȣ�rF�4�Ve��(d�w>��hC䖮:)�ҁ�60�J�GS�LL��D:�PbJb2�Z��4N1��4�,f��"S:�}|SS"p����W�L1�ƨu�UQG��F>�r�)�����)!k�3p>�aj�{����[�vgo>P�Jo�����,��L[��=�2�rħgj�d���Ǉ��t��3"p�
��nZ�Q��VJ"�)�K�%��jj �cd�8
y�8U8�')(��ٍ���~����{�'���y����pyu������޻�;���̵�<�G�n���~|��^����i��~{w��8�wO���PԊ�Ϗv�y�� ��p:�tطr-�p��y���gX�m�Q��%�
�z�+���c��?�bu��(�I���(�E��F�td�z�ԏi���kR��iʦ�)Wz���P�1S]����t��B|6;�Tb;o$K9!��j9@�� T]�l�$���)w@��8E5�:���U�`�̧�e&��,R
��M�i�̩a>�,J$)x"�7-dD�3S`x!��7�̆��hm�4D(2��Z�-"7��_�/�Dv2�����a�L3F�ju�d�L.h�6�G���,�Mp�O�*�I��&p�x>�;�pjIϺ�wz�7�U��%m��d���$�+�8��A�Bl�82�G0M<�Q��0=��H�t�0�q�L
�r���<p,}ck'�&�1�G��x�M$���)�N�5�a�"Z- 'Bu�3mo+*�ь�4u���DM�����B�M����Qq���1\��rdq(��)ZE�8|"阎A�*�����6�ZBU�"�h��;�'=��J�Y]���f�A���0�)TzQ���M�6�D�|���[�?qj9���->�!ҁ�Cm49��q����pc�� pbz�7E�����[z��Zo�'I�I)���NHR����R�)�~u��t��W)8�B�i��KF~�q��nI��G�c�_mm�z��FӔ���)4�z����Ap��I��)Z{����S�2˚�%�m�1Yc�I!Ȓ�D��q��V&4�e�'�?���!dCXQS&�	'�Q��R65:3e��`���q2 q S��)���"@�q�R?M���Ud���%Lʹ-~H� �]��S�t�I'�c��i�&����_�h3�@�8Ί*7���b�2��kʦ�B4k�Z��91C�%���ƏL�)�7"�SbRߡU:}#��">Ǵ* �Ԋ:��-D�_�U�֏�(���f���e�<K�HI
��Pb�ԀSKF~"��9�gw>�]�.���h�%�N��
�5�:[�Hsc"W�����Z�y:89�H�݇�q�h��X2k]�������uEѕG�)::������R"�����9��v�>�ڌ�����~��l��c}�G^�rYԗ%}�����^O/=ih޾z8��>%@3[)��� �YK�������ч'��C�������z�9��éEdk��V��Û��G�E���̗d^_��ﵱ~y��ַ2�0�'�~������M7�]kwv��������4O����ju�z�����#E��|h8pS���E|d��f,j�'�Ydʯ�j��`��BQS���>���+=�W4��D�BSh��L�M����s���0M�ҁm���� ��8L���
>�Q���%�����O
�TL�S�B�@#�i��22`u��Ҹ_��Qb�%��/�����4�g�zA!��ӴZƖ��#Kg��J��L�t� �f4r�:��YK �Y�,���ڸ������9���i��ӹM!�Z��)���� 1ģ��.���P�V��i8u�2e�B�i���{��R�K\Ի�b�����>O{���D���Jd@ӪHl*�������CN��G��h«�8�w]	�5&��o�L�'�F��0��t]��FS�Ⱥ%��~�ӟ�����'?�� $L�~��E/���];�hZt�x��m�Ė�	�m���,�E'+������U���'�7��:��~��O��O�����_<}rq}��׷�����+������?3�m��L����޾�����~������պn��/q�*N�������󻇋w?�����W_��u�}e�pw�����k�Ij�^�s=P5���� �/�z估���!|֮R`mA;�n�m#r��H/��!�7���p���>�6��w=��Q�i�+G��+�v����6B�O�6E��@Y�S���ֈo*�a�4�D� ����m�i:)T���:B�3��0�)*|�O]������J_9R�FV��� �6�����ղ
��fK���)�&n���H��IG��ƀFH#{�I�);C��I�@���9�U�����R��}��h�~e�h:�P�n�_�(D�d9Rڄ�A�.�u�&1B�*����7C`@�
���'�`3����[��2�,k�!{[��r=��:dE��2b"��=^L��===*餠.G�G���&��|�1Ȯ��A��4Rk!hv̨���
�hoj���tѬu~U(����>9�FY9h8�鐢�m�Q?����b����b��n��酌��<��_YR�g�G��sO������w?y}~����on��wg�T�_p⯟�p��	���9^!�)����wG''���'�����������Ҿ��[i���:���g3��L�iu�6�T�3�Aazf�QC�1B� 8n�ܶH)��	��,N�Z��$�@���5	1JA�c:m���R�$�Ҥ���B%9VėU�!ScÄ
7Vh�L���TD�gU�I!Û��_�)��I�۞l��Y:����X�~�uU	�P:��9t�*�Y��~�� z��S^b��bĜ(5�,#�m�o��4r͔R�͗��TB&8E[�r�Sh8��R@��D>#���f���q��4I	U��� M��Ղ ���\�뎊eA�$�I��9��Om�?w.�tz��i&�G��7}�au����"�	�g𘜢���R�Y�i:e��/�d����Y>H�=�D֏P�a�!m���E� �pRMNsDM	"�X
B'2�6�@�)� s�f��ےVĢ�Ц`��xO���%2�Q:�Q�����?d��M�c�4�v�B�qu�)��!���'qH!{(�l�|��t��42�D�aJ�f��8Y(&)���1��`B$r��J�QTV������+��hjYW�`���E�#�,gR������0�1���t
�pO��Z%[��ZB�75��'���r�:!&=�h�a4���Ȝ8Q9U��@�w�Z�d�Io�Յ#đ�p8�4u�%�,�V�F6�0�S��M����s=�On�	�Щn��/�H�Aв��ė�Zid���!@J�45�����[�!Iͺ�A�'Ę g��tx��B(��T�v ~�	�&ͨ�i��Ȭ*�:��O��-R9c����1B8F�H��F"�MJY�����rZix=�p8�g�<�S�<�#��V���05`c�|��j��Pˢᘦ��$�i���1�,S�=k���%V����@iV���7"��o��\`"�m]G�Tt�o6G'YYc��c�98̻��Ҽ�6Rf@�TLЈ'���������_�i;2e+-�U��)�Z���s96v��]���������zpy�����rί���)�����dJ\	�ճ{߹��;%vc���t6�I8�/��ۺ�<ON׏sz��n3��t�tpvr�����r�$��\����+�e�����<W���Ǉݰ:���֥��#�����ӳ����;L�P���oxʽ{�?98�?|\�i�������ޱ:�88����>~�v}Wu}at�P�z�������3h���^��� �Jݹw��s-v{��p�]z9	;�>�[��)&���5]��!ٔ�k ���:@
m��p�.ʯ��*m�~�Z%$>��e�V^ǫ%�k�_-S�9�� �i
�Ooq�sQ��F%j�1���<���p|6�H����1�	J�P�)q~�ts�4Rk]f-pV���g�6��*<ǈ_�u�����4u;�4oi�MSMܴf r7�L>Z)F~�B!S}����h�&}D8��t
�!)�(��t>'~j/`| ��iJ�N;V�q�	a�=;1Ň`�?#\�f�FF���`�*5H�z�p4%��=6�v2~+��N���>����bgɫ�mE[G�ތ�rh��EK�K|Nf���g?�����]���l�8��|lB�?'\�bB|S�g����?�|}��#۾��ߺW�o�xtuD2{�V�cj�p���6����ÉN햎�ڻV�"�q�hZ�~�����*������_���_����������gw�r4㖳O~ӍfO������/��i��s��.���^d�}�E��l�$p���N�~���WW.��:~�|��?�W���Kp�7��*��u��g����������nɖfl����=Z�l��N!�#����IR�"�B�L��1"�J�1��w��B��u�s�M0�N���i~�rt�W���F�!�aC��w�1�c��_|��ߊ�4�zH�HA�8������uĩO8�ц�PE�4��dF�e�����s% uK�S����m#_:qYF��V�N�q k�W�BFQ��'e���ZB��W��8R�p�5ơ��F]a�ɵ(&NM�V$�����VQ]馤�pL�t ���<�HgȢ:�Ł���Wzdׄ<AqzjBP�����R�T���-�&�*ּ�4@�I�(��IQ)��fDPQ:Y��pR��D͔#%�6A-%F�Ҟ��e�r9�j�ҩ(�d=���=��a1��a�P����{����Fȯq�מG�wD*փǾ��|�QE��u��u%��O;F�ވ�L�(ȱjNkO�QH:���9?�tL-��!%��lڨU���R<��O��F�ݬ��E�Ɏ�*����ͅ�p_}�p������������o|K����͟��_�n���/_���w�g^�<:�\��<���?~�'��h~w{p}�p}�/VW�o��o�����O_�p�z������\M�z���vv���o�����LH�st�h��ۍȍmx�5� �pE���L);s���V����\�ÁPK���^�
ё��aL�ڐjI2�R�S�"*!&0����?��	*ǁ�N�Dr�
��6v���nP�#�x���r��>'�(��l�Й9)�ar�p%�lxͫ+��B�	��(���N	䩂�_.�E3JI\�mC��e��ڍL��D�CHՍ�4��
H�F�E�қ"tb�	��a����SE !)��Il	�!����BSzj�@SYh�I��>B"��~ |#�π��q��	�-�Vh7��^z�!95#�$5��8@��s�F�΍�!�1�)�S������W��vA���*~]�s�)�%:���'}`�Le1�Ģ|M8�Ȓ�$.b�$��� �BLہ��_�TASt4����.~��X|V-Q�0��2z��~9��Ҕ�fJ	�oʈ�ϟN�P9SGK��3{k�ѱ�9�r;�p~=sV՗gr!��p=�C��ALCr*�Ծ?�v�NR��IǶ�So��!22$�,!8�q�_�ڠ<E�4J�`�!K����4�|�{9ikشtY:�����BF�Z�&}����XԒ~�e�J�V�(TV��J�?��4˟PY��Si��K��/�"G
~�ϟBl�DF�J��,�h�d!�����Ïi���HD� ��a��)��s=�$�Y��R�i��Y�S'F�)Z`Y�e��N ���K!���I�J�k܈���#�1&U��HQ��i�ڇJ ���L�t"K:QoK�C�ΐhu5(oɘ!�Zj/��h*�߸�_H�~K��&�(_�(�^��r>��Sn+������46�A�G��.�8������7%�4��Њ��B�����!O3�!W��3&���T��P�8|F'�\���9�cZ2��8?0��R�WC�Ch�h�ICV!��Զ))����p�ޒ��m:��J�b��F�R�b�ZZ>�a��U�9�:�:L��F�čz��,��݃ߏt~�k�}4
Zm�����`;������n��.�@�=4o�}\]��.Y�Z��ߦ�.{]��ca~8ӧ�O.z=u���ʃ�ߥ��έ�r'�.B:�����[�1[ݬ�Gs��m�ܢ�{���Vn�W��Euۤ�}|�.>C�i����������_}u~�����t�{��f�tru����ۇǓ�k��~X�s� ��wflɓ���l�.��\?���N�������֮��G_���@��C����PP�/�(�9�L�t���f*����1�,mX&$�4YB�ç�>��6�)>�鴄iZ]��19�ъځt
��&���ϖʍ#W����#0�Y��UL%B�A
y�q��4B7UQn�@���ߊ?�^Ąpj��H�G�305LfژH�)DS�P��A4�$
I1�c��3�R�]���Mz뒛~� �g�U!Lf�f��~ύ}�zE��%�����FV�Z��"HV4B��0>�S1��.��L�8%M��llg
�釔i�_��Q��B�ִ�VL K�4�7b��I"�-�9B|�(�$�Eփ��Q��6�T��ZYM�9F&��)��Q�ǑRT!2
>�f�"�Y.�k_g�NL�j�Z�dA~���|�-��^�5��-�z"��_�I��BQg<|~Y��Nqx�X� mDO��� p��a���+!��L��O���?}���O�]	xs��v��1��i?K��#��(;w��l�~Z����k�{��G��^�}ݰ��X����՗W_����~{wp��?F�_9�}=�����{��E��ʁ�[���B���g;紽*l�·�p6���86ak���ց8t8��f�����֩_EG
�� �jș�y�����������DQ!����-�r�=r�L+$w:Q��Ѥ1�oP�uѧ���tLg�KG]L`ˁ�I�0jp���4Y��Y:`m�c9�p �ҁ�q�p`ͷ]�Po�@`ȦF��NAQ+�=�D�Ut%�qجB
k�*���_����RA�q�雖�/��	��Hܨ�qu�Y�:̗H_�i�Q�Q�2:�c�h-z�BD
�K�z1�FSL�.�´L��V�U@L��s��+�j��**
)�晳5j�~4��lY-�����|Y��XH��
�
��Ѻ����Հt�ѳ�G���@�J)0-q��O��    IDAT5�7�]+�kI��_��>�����4�"�Ҟ��'.E���( 0�r�BDp�����*�o�!hpR�9�1A8����+gM���/~���N �����e���k��>�;�}����Y��/��oώ�^{�8���?��y��������ݏ�ٿ}��<9X��	�˄;�<����-w�f~��{�G��qsywyt{�͗���z���?:}�;�W��M}�עl���'�V����v̨�+$���pS���vGg �B�DP"K9��4��09�Q���v��8�c:�Jd|�8R�_nYF�����\HY�|6Y�U{3d�#˩%�}�hiV=�d��g�c�\oo�ҁ8L{�S!D�cjQ�d�M�rq8Ѫ� ������1ˬ�����#�o�J�pFV.���12x��r��dJ'�`K)W�o���;��
lF!�Z�T%���OpNB)�.W��p ��'k���B~G���)6A(�O�r�|!g8$r $����qXMҟ���3��ҙ=�	��WK'c�56!
��[i��li!խբpV	��)*'}�D�E���p�p�8�4&�)!En��a���� ��f4
hrZ`���L��'�C�T=!/���p`H4~=p�7&�d����e�jr8RDG�W�BkL3��<4R���b�ii�p�@~&�#���)�1����LcsD9ƖFӴ�8�Q��ƩV�Fӑ�0酀��$��T����)G:���q��`%�Ә��NNb��f�����7����Ҕ'��єMK�8����\L�q応����V�h�1��ن+��/A��O��H~4
��*ٶ�)MH�������h��`*�fZq$Vn��	�t�D�hU7"K��b�5Pg�[x�FV�C�>��2�1 �����L���5��5e|�K�t۔�v,�t��Rؐ'1�(��!���ؒ�����&�T�*�ڈ�r�y�៑��*�Ȥ��ũ��2���֘�����3)c�$���p���pj��1�J'������j�`�cE�C�I��NFC�{F�T���I�g7*�f�#��f�ǟ49���mZ�H7mW�2�U��1N�S+�W7N���!Y5C��I��������I�=	7"g�`�9���i���T�Lth�iD��T�B��zyJ�����H�����w���&�h�S4|g񢭴΅4��匵��'��:S�T�w��ƍ|t�;��|� g���f��m�����Ϭn\�|<Y��^ֶI-v{������'���,ۮ�a��S?K那�_��C7��x��=\ߠt]
��/�3�."��l�-���,sqT5뉖���"�ݻ�����d}����޿�n.�v�?xS������j���/|�����×������������-�����Ʋ�\}��x�ȹg���U���W�v��W�r໠>]���г����m��C�%��)�����x
i����a��/�Kb�r�[���k�#j�9Yhҁ⃈z�K�~}�Ǆ�X�����r1������i�u�2Y���q��,��DY��Ԁj4�#D���J!X
����,Z)�5�q����|��I��B!>�4rE�l�n
��t4��lG�Cٱ�ß%�Zmo��;����x��iZc#$�	YT��ΑN����B�1e:G�r9��$�*A|6��� �0O���&�vU��"�P����iF�qGG
�H�>�.]��X|cu�jJ�;j8D���+�������L<2�NV��9�*�@SB'�4�ȗ�"���tp����)��CS_��iQO�>ބ[�6D���$�#ܿ����a�G�E]����+�_hY�y�Uv;e�]�;�0}3e0���5��d�܎�^V)ĩ�)kZV{��h���gn	��n�&�klg���������Ћ��:s\f����g^��>8�ϼIY\�zU\�������mO<��w��rzw�6�#���ğ�3FS:_�f݌������mZ��=��ؖ7�CK��X�/��8V��1���g�W�M��#�I����7�\���1&�VUl�'5�O̝6_������љ�:G�Ϛ�T�g��3k�
E[#���^�2s�:;}F�iu�gEhjaVE� Su�t8�%kDP� �tȀ1ժmKS"A#�)��SV����?D?���	qT�I|LmH��HA(q���K�!iR��PM���r�&�|QS�5l:8����*�6�et�R���oE��J6U"�=�t��`�w�Je����>5Ӯ���m4I����X�B���i�qj�Y��sD)�BDۦ�a��N'���'��D<�rd�ŇX�TbC�pW�ɶ(K?h�)�Z(x�w	p>s�Q|Fַ0��K����o��o��!��?�s�~��{��d*�,
�&��S�|#��1ڐ��S��%�Z#&�k ��g@~�F����D�9�*��3[Ĥ[���m�}w�[A[�iǳ�7Y�/��·�߯~��Wg��~��so��N�.w�^)�����5*�u/��ͧ���g���.V>]�_�]~s�t���󻣛��������?��?����v�ګ�[�0�-ͫ��[/"�+���g��+˴��c���X)��h�� ��k�`%��1v"�=v\�T�Id8F�������Nl=D��4֙lc��yV���?�D&ɧ�gIqd�?��q�J#�tT�ဦ�H.N��-cZY���ïV��u��0NY9|�D��v� � 0@Ͽ_Em/��W�r1!%�`N��1D��p��-�h��
�R�x�
E��Q�(��e1
��rL�����4�E蜑�O��SJHUd� �o5��d����9,M���IG�΄ҔR��K/bڪ��LJɊF� ��Y��J�b��Y�	+
d|"�h��MK�(5d#N��8��z�Kv��ҩ=���� ����������R�5�D�#k_0����a��=���0[��ZӪ�H?�Y8e�S��	�ƜL�q�	��� �ڔ��Vɚ5rf����`���nZ�U'�_�,)�#%=&7�g�O9L~ˉcTH]d�Q`�~ G:��@����,f8�t�Ь����GP�)g�V��$��=��\]HR��\]>'?��ۓR LԔS���U�Γ�O�N�J�rD���C����H��|Ѷ�Z���g���2ed���K��P���kc�_�@�X]%D�����^j�ڨ��hm���~)d�0g?���SŔ�v�S��\]!�}�V���7�,F0M�Va��,GV]	� �7�T	��p�Y"U���1������P���B� ���7Y�[x�M+dZ
�h�F��$�N���J��h��ib7��V�i0�QS��O���DS@����D�r�.�f)FS�#+͢B�|����C���=K�㣱���(
�N�BuRW�wnT"5c4)Ü�T
���#������֕���d��)$�	Q�В�D�=��ԿN
���yޱi[(>a)n�-����il����m�ojmJ�я�/n�n'���3>�?�PQ��$���*��(.���z)F��huˑ>��	@S
3���(�{��wLL��Ʌ�� Y�ȉ����2�j��LQ�ۃÛaO)>
}Z?�پ�l��(�΋��%>�|y}��dqSYW+ŗ��`�k��-O����뻙ް���?>�n׷B�n���N�_�_^��݃��3rws��G���WLo���;�+��}E��D�9T�㦳[�Z^ϊSoX���y ����h�*��"'Ƀ??�������������˫����������7W��w��J{�n-��X��5������þ��t=r�������5}����7-��[�Z҉G�ګ�yQ#����ka�)�B�(�I�,�_��?:)���1�Hm��bT-��0�I�t����l�"��J%*Z�B�6��P�+Ē��ee�k���[�i�uՒ#4R�F�)|�C�Ģ	FJ�>3e�6���ρ#o��ߢF�F!N����褐9)��]j	����NDЪ��U���:�f��	�eCJ$վUy;՟�)~�U��V��R:R�iN	��c��,ˈ��਋@y��d8m]�[��*���Jg�P�vI�\�B�4�i��S���'R
�(�U�'�g3�V��) �C�<fQS:��B��ЄX� ��O�8�Gz�8S�2A��@�d d:L����y�*v�V%2!�p/
^���/�c!R(k�M�|��sxc_�����Z�2>��]�>��1�L��h��2T�%߇�B��l1�@L��VTJAJ���Z���R�s�q�Ћ�[�ݼz����7>�������������7^e�����ۛǛ�����:;ן�C�M���-�ɩ�+jsw��k����$Ƿn�w~2���p���[7d?���I����[���T��G�����n]:� �m�����QQhv�eB�+�]M1��q~��IgtD)��l�_S;��9�|�=t�H�ǝn��������T����Q3�4}4��!í��}Q��팂g��lG_:κ`#]3�ښ�Q��t��U	�Bđ�0=K1�ŧVE��ӗ�3͈�\<�p)Ul+�r1�p�4 V�(� a����E���(��>1�h�*�M�>)0H�YL�1�.qH���p4�8�%"�G��s�8� feMu�Q�{�q����!η@g�Q'��xêh,�V��@��Z=!M{�I�K_dk�ՙR�p(`j�c'G?�~K0�G2��*����D�cj��#��S��F��_ot�{G�=83�?m N{B�H��vn8.A��@�Q�(#�I�]�_;.���q�dh���F�t�Zf��Bu"q�ɒb-��L�D���X�'���3��t�H��ӟ���zc��������'Gެ�~�����ԛ���^�?]}��%\��]_ݞ��ߝ�=Y?�V��3on�������}�������?��:����ޭ[���;x���'���?�g?��������o_��}���9>9r��_�p��or�C�o�8��&X�琉=p�����<q��muS�� �&�+����������a�$r�N����J�h�U��[��5ӹ'M�d��rAX��+����R0��F��V.�ꪤ\
�!3!������p��VV�}D
pp��z�k"U�1�Z�Dk&�~�����1���yu��h-R�e�P!�1[o���U�Uh��LUG�O�	����6���M��i����}6��o�¥�'Q���vAZ�(NuӔ�E�ϕb�	o�����dS|�oO8RnC�ChF(�(�m�vZK���&r�8)�m=5M�O�i���BT�>+!�Sn�	dSOA���	��0H�����y[{��3)Ѥ$rt��� đ� "]�-k#.5NuKl
�b:�����m9���~&e��Ȑ%�����>�UՁ��h��� ��G��\�r���~���̔&gZ�O &�D4�6��3�!�Y/U�sF�8S�t����ҤB�rp�@+*TnSL�P+��1�l�/RW!�Ȓ�8x��Hr���q�V]Q�"'���l���3�1���*'eg�)���H�B��
��fg?�}���{��MjJh&���#�('2�)>&Mf�ڢ����!�Ď5���*
qr4�2�Oj���A8�cT�h��DbrRb@|N+�l������Ui3L)�җ�!״uY�ru�\#N��?�)g05`�#H��Y���V��~�5��M�����h	"��BSL�ê�ôp���dL������&�A"pLS(
���h)F�>��cO������s�虵(�)Z��nzς��_'3��$�T���_�����S0��i���.�X�(��$V���DEd}cR1qL}#���d#�i�2�� )k�>��@�4��U�t ���Z@����Ɇ�a�_.D?ӳ�D�:ə��"U�(+����g���������VWV;�T>�2{�拎�����3*�����Yˣ������_����������ۅ�աO`�}Yow�'{�{�%�J_%�}���nFO��e8�{�޻�y��x�{�_��G���N_{ʼ�}���S�ó��ow�l�Vc���x~z�����z����Z�:l���u�ճ����_�<=��`�������c�j?\�8=>�[�:��εǾ�oG��O׷>�}:y{~���z{x�x+�G�D����O��n\���Pߺ9t
�1}��6McF;ߖ���1�D���q�ф���͡WEH�8�����{��Y �8�x4�1.��z	������LE{�@p�䴮ʅWEbg��'HD��ړ��6��j�]2�%Y8���S 2���8B�Ə`ZJ��ld�J��q�ʯ�J/�V�q4�b�bEՌ���#ԡ�4}~���7ř�����9���U"�(�h술qL�4�$^��P"ʙ��B�*��[TL~�1#BP��vCn7e|O���e��U�����a�S�,�(��>��d��H
_'!f
o4���'�Sb%
AX�(]�Tm��Zˬ����v|E1K�=R9p|�a9�4f�H�c���D��duX] fYS�,�b�������H|"�%���U�B>���|��B�P_V���?�ܧ�D�j�ٹ���>.��*��z�Z��q������)��uܳ��!F��,�o��RD�!��P��s|u����~gS�g����}�f�Ɍ'�;Ϗok�g��:�����k�~��{��C3tzqr�ʫ��+t/l�~
.<�<~��/�}���oo>�����_�xٺ��1H�1���@��ab�f��������il��r��Gk*�I�hK��3>�H|5L)T輡�9.��9�ZY��T�D��)ᒀK�R�И�6��rr��e�G'kʻ�J�,�:oT�,k7���h8�!
F6g�C`h@F��M��\H�,���y�II��� ���R㈪U�؊���5��i��)�j���!��
��"���#äc{kؔ� 5O�/��7V��f��N&;|E�ጦ�o,� D!���nsl,�r䲀ei B�Q`.���U�ե��GTV!U�Q�@L�MM
(��uq0���LP�c����B��99�TQ7��*RK�EUZ��)�WWozP�*Ff],_�J���I)��IW��x4=^l��L���j��G�oX�駕q$ҁ�l9��P�=DP���B@��-2g��cJ�/��I�MGW����Tע0D�&�!���;t�¹isl�Ms�)����|���������MY'����^����ʍ}����z�sr�����u��{?P�<�^��{r�pxr~�~=\�<8;��ON����ͻ��^��o�??��o~��O��9���_��z�t��i�/@x��o=�����˓�jr{p(�Z��c�B�6�/=�,�"; �����l����F��y{%��<d(�gc��|=Ԇ\&��EX�(Ę&��p�f��� ǈS�Mk���q�@�um�B"FV!r|u�����6��rʭ=j���!�f��k�ڴ8SN:��T)�(j�*
�(�e��E']"�}������>B�M٬�/���\�?p��V�[���j�j����T?j���t)Bq���@�E�j9,�(��ɚFH��_�χ P�q���éĐ�|R���+�K��
��.̦�	d�wDT�պ��n
�W��� �`��+gd������H�����^Ś�G�e��瘪�@d���S(&�D[�iQ�*��pB93U�T=#�dmX�S?��BL	 �e�S�B�z��~i�[�z�W��ގ�mJ�W�����#��\!����GRH��rh£�����t�\�r��n���F��4��"�G0�ЈH�늓o�����P`���cm�V�/�F-їÔ_b% ��k*�Q�^�1�Xz~S����0qJ�6�%��>B�����$G�&�0R�i��1D��t-��iV����Z�:������O�%�6Np�m�3��ѴB)Oo���>����r���0�P�^4�Rf���Q|%8)j�,��C�P��    IDAT�QuU���J7J�����+W!H��|�ڎS3568�Q����ϊB��H�?Nu�9�,��-�48��ȱ����A[�{Y���*���L3�pV��G�~Q�D���c��@�/^�)$bE��cl��� 98j�PH-p����(�����(`�g*TKv�j	����M�[U�����pj,q"%r�S{!�Yd"h!��_WjM�ȢC6�wjMhl�pd�9|�,�NFS&T�S˿Z� !����J�*jlm��D=YI�F���TL�B@~#q]��QW�4�|�,��ڐEJ�IuZ���|�>22�
�l��R�&�;I_�\������ ��=�
�og.����J�sOڝG��\��Z��U?��Ҧ_��m@Ի�g�?<}��_�w�OG��⾺x�Җ���)�ۣ�O/N�����q�#ߩ�R�:}����uK�$]Aݶڡ\�[w�][�S��/�M�����j��vb?��>������NN|G��N���ķG��>?�^]���|wxw��;0���F}q����#�?{�z0_�u��	����?fV?/Ϯ�^1�ܚ]��:|���#�6|;ʘ�����f4�:`�E h�jJ�T�i��#��rM�%e�Fߺ:�E�U�UK�Bi�cB��1��^c��B��Q]8B%����҆i>>��Uc�@�1k#��ґg��3�M��qǄd�9�h����đ΁$N�Ԙf������$�}������oe�9�S� u��Fu���1V������c�=.�������_m�� K� �P��z*F)�B����2Q�D ��� ��*G�)e k�*
A.$]��!#+a��[���)dd�[c�)7Ja�9����o�L{{LIA���A6
��vQ��v�ߔ���ocg�pL�q���M���z6s�2�}����>�X�x=���q�B5�>�V��������WR1l�|Zʫ�)��0��_����[����*D95��(?�j�R�^����^�����������&oO��f=B��3����75N�N|����}���W�^����1���������=��G����������˯>�������7�S��w�Y����:D.j�p���7~�g�t�G�i�H�ي�U{~�lI�0�,�i{��ګ��A�?���F�*�>�z��� ���q��" �;(�
׉�f�ٔ������i��C32�l9���#�3[���[ڔ���\:qYB$Ӥ�#���p�Dt�բ����h8��"��>2?�4M #�#�
�q��t����)�������h@�'���l*JS"����Ǭ�U�/dl	zP(Y��� ��T{��(Loz^���w6J�Y+�Pe�4/�T=�E�(�}����1Q �_�0b�-�x"��;'��1�HTSJ+mo!]�mQ�S��D�����������)�I,[�'F�՛��UK�#hX?��B�h@9��Q�����?�f-��[/ ��g)4Un��)9�Sn��TE�[��!�N��9�m�.��}<x��}E߿s����x��ߞ\��������w:��~����?e��d�u]�=�uA�J���
��C�p��G�M����~��n�m[n�l�4 ��B]�������#�/=	��k�1ǜk�}��s���>����cO��}��3��'{���� ����ho&u�<;��γ��n~���7����_�οy���������j=�Zk9��nS~���ڛD=�<X��<j�i�[�,����VԺ��B(ÔI��<�tKZ����,֝0qg��;I!"���$�pS��-�u�k�V9:A�)���O
�g��jS:�ҁ�lYƜ���-�(�h�84k��F�M���\))�����<K�2�&���i�2�h �!;�[>P��J7V�\|�B���vPR�u�:v|��N��abBX� ���'-&3�nc��8Ӝڐ%J'N:j����i��gD��?[g"�6�~g'�Ʃ4�D�C�X���&Ł0)��oEE�i�	~�7�77IL=oe����f*����t0�r�4��Lx
�N�'�ImE!t�#!Go��4�@#��r@�3'�f"	bF���Ǉ�!�[�ҷ��]bY�3r�8l���C�h���#���[�,�����˦"_Ho�-�&Z�S���٤�YYiq��r�hՔ?!>�n-d��2�d9@�L��s�8��{�6pp;	� ��DF�.�iD�<'�jl4E���HU�,��ld��+�凛�1RV�h �fY8_���D Ӊ�4�OR.�:=�L�Hs���#�m����S�&��:��HL*� ��&V8��B��_�ƚ�s��R1ĨO�鐊�Nc�|�3��,c4j22�1&�#AD3��� q&+$5ஸ�����B��<ʤ �:R���b�W�מ4m��ԭz-q�s �e5��S9����c�� )pX|�[.Uh�խC!�I�Uv�[n�|k85�H�[l��%:���t8|YI�����Zܣ� 9�V�I�I�c�ϩ�+��r>Z= s�"�J�H��n�"+Q���؞��
5E�N�!Fj��k�OJ�T�])>��3�LS�O
�t�RL�,�\)�ϊ�-�#�8
D0=��|QH�p��gh�kϔ34�����g�Bh�K�I���|֢ �4(W��ޔIiDS]E�D��G����|K0�Md�{��)���QnnM8�l���R�1�Ux��j�n�r[��8�^c�MB�Mnwp�#�,�Oj��Ny{�WT��\�>�i%'�Q�\����z)���j�x]�Ş#x���/^9�����u���Q���G'G�>��z���c�/UO��_S�)J*�&�z��ήiUQ7~��]{���`#(���t����%P���gۧ�����;��yu|�~�gm�ݕ/�{����'����o._�_�o��ү�y�#�^#����G'�����%T'�CC��dW�l��?�	q����i`Bn�n�ys�
O�,�!��ў�O����II�O�L��H��-�Lx{�sR��]+fx"�@c:𲌬��H�x[��K(2�^�3mB6��eI7M�Æ��	a�ʈ4�-q#Pz�ꊲZ��q������p
��{�\T��8��tWi���;
�m���g]|��pY
A�M�pJ�Kf�)��D��F 'n�H���s�u�k5���&b�� ��2�k����,8�xG�T�RZ~S��~;p8RT���0"Rb³t�A?�Jf-�Mi�ަqT��AJ�c����PR
�מM��B���d8���v��X�8�B|:FӜ]$&AY:�E�x̍0)Jx��vn�6<���Gw�-
���>��5�+�~|�#��ҽ��ǎ~�����?�Yr,G���uS�2mi��5�X�t֠�u?���v���%�>M��^��6�_�6U���Ç~n]xx� ��>��R�oew�:=8y�w������?������Ƀ�-���HE�?�UD�������{�z���^���w�ݿ�zy�ڏ=�����V��\W9�JN���(��*�u�i��n��yo�BcR2!N�|��D�R�EmĴ�D"M��Pu��t��?M��0$.��&�����ⵏ�ti��hj�Vu%qQ5҄�6G�9�:� ����쀩D����sH���ᔐ2"��r��5ÇAˊLM4͚ѧD`�u�O
���R]A����@�a��"�r�*V��/��t~ʦ����#�T��!-&ЖB��,�gD4)��tb�v��	g�ST�(
��%W�Z�#�+��tcw�#�����-��nJH����S�|��|�q>KAf��<�s��ZU.ǥC×G&eD��u�H*5%8��?��tT�G��PLM����9���HJ�Q���m;�&���D��-Z��m�&M#��D��h�'k9F�VT�F4`4!~�|��t>�3�I��_�P)i��sL!wGb���ǒm�M�X�t��p��׏���_]��7�z4��w�}�y˕����<���}�����?{��y���ѻ��,��	zw�.�N�� ���n��G�~r����}������v���.���Ç�=F������V������ŝg���zp�M��y�.��\��Œ;,P�B�[����4����;p���ȲM����4�e@���C�LYH:�޴J\"����;�(�~V��U�X��ce����v4#BR9e�Y�(_ԘN��p#f{�2Mq�V�1f��R�
��p�q�J�؈ d�bN?2B�14� �i'�)E�#��#���BqV����Q��cT�Ç�?�hR@#N�T��	I�G�FS
�;�u��x�j��� eUTM"�3%�t'3��)���&/d�4N�\�q��Hjub�qv�K���&��0�RƷ?)Ǳ��W+)c�v˕�x�K�o���(�É@����/��c��V����`jS�Z~��_�q �8���V��_S�Bjqd�	>?Ax]���7����ش\LNK淐B|
��ʒ��;��P�)��b
q�!9�T��am�jC�:���1�,��g{
�4�H!LY��HwȢ�h�nzon>h}�qj N�8�NK����
�Ė�Po98���Z����9���R��t���u��$��,�}���ʖ�F??�������n�Ǥ�`:�h��i ������N��f� 9K�(��ubĄ3>)
!D��
���qFpN:���9%nu�<O� TK����ֱ��,�8)�I�1����T"��H�����'���)�xoon�
��H��$�/�!P�_N|Lx��J��I�J1��|�0:��qԢIU:$)�t��>�6�=`�'��O��iʑhd��@S#Y�	q�%v��"rOV��ќs��&���)L"AUDq�S��B��|~]�s4�m�j�X'�*iEEIA��#L
Y6d���l�r�
���c�&��Q�-�lc�K�>�i��8F4����2��1�*TJ
�z(J��=�3x��SV%�Pi�^OiJ!�����hڮgʹ�ai"gh��U~g��J$�B���� �FPE>&��ʥ6:���'}��я\�BF&_�J���B����%��Od}���u['�C��⦭9yº��������N�<�v�P�g�����Z��ȇ0o�z.}t|�s������~����9�o�]�<�aς� {�G1�X������y����\��U��"ZZ�\�$^p�^�v�W�eY�Ճ-Z�WkQ�	��c�a8+n|���۳cK�
��q��]y)�����3=x|����{O�~usw��O��˓�ӫ����z[���ۏ�y��凾�֛�U��o[mmc�;L�F]N�4��YΙ���o����!ń����$qs z�N$�)j$�^���
A��I_{�p�%���"8��{�A��0S~R�t�!���/B!����LH��=)@�G�R#Y}*�ЀB�|�JD���X4ڦ�V7��0�d��|�i�ȅ	�P�1�S�S����A�Ȉ�Rkj4�4��|�d;���p(�[�UȪ���IA8e����Th7K(A�s\�Q�M\Zokq&ͪ��"���p5_n�gsr*�[�A�i	�\"�BpV?��*:���B��缕�2|[��rk>M7������C� 8p�e��A�E�OS�j��_S����Ph����t`"���Hn�)��8:rMw)�e)��XE�>wh�b�:ӏ?���?�)����Onx����������a�ڷ50*�Pp��F�4��V�vG+ڪ�1�B��rӭț''�"8�=��S'�c}�ꅷ�������q�zG��.O�^�\x8���s)r���������<y���|��k�����c����۹�y�]�\��������O���w��3�Z�.7�_�ٿٿ;R^W�{H���,I�a�1��6�b���9��I�P���f�,_{b�)iʚD��m�iR�H��ʶ\jw��iXT9!ǅ�q�f�dr��#8"s���4b:ÈT�����%v�8�z��g�H���R�|!�p0}�$'�B�iR0�T�mZ� ���$*mS8�c�ɪ���q�N!�(��h>��t`MV`&�Fq��8�D!F6Hj�����,� ��!�:�)W4Д,�e4�E�7�5ic���s:���d��!F~���!�T��0��_-
�j�`tX�";Q53ˉ��j�)r�&��t���\B����
!��q^᫥4�V���o�rL�B�UK��+E:BUL����
��uH94Rr�u���6{k'�g?�����[M�]⺓a�QEfjD֛��ZTݶ:8�Z6���N����Vo@�[�uA�`��0e�h��=�(����+$�h�ˢ���������7�WO�����wpr���~{}���g�\��6���G����3?O}���������/y�������{���~wٓ@�w(�]�����wN>������������ыg_�J��o}�����nO�}y����'�J��C���pX�у�c���vbs�hFS)�b,��ⷍF!#�h+�)p�ˊ�ѡ�5u�:P'�*d�l)Gە�M��	�Z5e��[�u�Xc|�||je%k����&&�"�ң#eL)L�ä�����F�!��#Cֆ(_J�7���,$
a��c:)��!�V]MQSY��,Dz�JG��Ʃb�ъ�'�
Nm�o�U!.��}N:�vk�G��,�i��:g��$�gdE[ G�qW��B�i�D�[��4I�F��6
�RL�"�C(j�!�K��d��[���<�#*+f�'$M>��CJ��#�X���gc�Ი��z��38dڀT�Eވo�[D���%�B����-dDn����<YU�g�ԕ����GP������i]�JOJ=Љo*�Mc��G-0���G�۹��U�F|#>|��n�H`j�50����	[�T�
\z`�C&�\���ޔ��C�\ �c�:�ck�t|��FA��3��(\��iQ��I�� ���Va�n�D(X�Dx�F�J�mX
<^-7"�-\!�)�n{JK��![B]UY���_)�����R8����Y%��B�),�@�u#�̷4H�T"��O?p����uUQ��=�Łg8d����HNmP��G6� )�K��tt&�M�w���3Nu�r��K��H*Z��@(�f�wX�!�1 r6%zfm�#$�ҎA�Iy#��*d*�fp8�C���lGʙ�)��ҙ,ۂ0�x��J�ßD�n��Ӄ�Z����h�h�FdH�Z��B[YGk;^���J�A*
�\Q���.C�,^(�Ghu���F�"����l���ӯ�15`̪���S��vU�]\
DH'Ĕ5�4��#�`6:�t�?Bj���B�ӄpD%�7��?B���I8���+�/�h�sȌ�	�A&jt��M��5����Y�qG�(eK}Ӱ��'2?��"��TS�4���|c�pp���a�@���E��F;�q
I�V�Ac�{��D���=sw��.\�,��w�FYv�M��©��{V1\���ٳ\/�hț5�k//׫�Gް��������g����Y_#�}~s}��K��{듚V��\P�;8qq�{b���˺Vz�wsq{�w+�}�R+�uU+Y�w{}�ax�->S�^/����m���=u�NN/��\$]K;:r������ ���}�����w�ŷ�{y{�ͫ��8>�]�־��x�����ׁ>XO��O��J|h��B��:�6c~�B|�.���9D����g*�4NG��M�f%�����^e��)��~���g�h����-���.�e�*
��A:����9N��Y�tUڇ��'��$���1�Ɨh:R%����EǨa|>Zȵ���Y.?��D���ԊR�C훨���� %"Hጥl��8-0"��^E�J���-�Ժ��t��U��M�*���!���)1ǹ7���B�[�,x
�8Z������J�tTڔC-�4D5��\w��sƪ2�*TuR��A�i�S��:m0�H��IT}�ůc�1Y�p�w��Rj��(    IDAT�/Q'���xq�I�hp�W�Dsj{�8D���6��[G"e��xE�N�&)�̑!)NxˬU���3���^�׏���/��B!�o>������7����o��o=�{����W��bݐ��VXm݋֖Bjg�h҉�crL�K/��:�c��<
����x�d���m�Q�|v{p����w�u7�d����[����<>}������"w'�v����u��ޒd�.mn_*�q-�����7��ש�<�����P�@x�z�S�~}�����������+�	���k�����*���h]�H��U|ۨ��曶���THz�v��%(��B�|Ʒ�>��@�+�n�����fYQ��ig��|���:
r�p�D���ę�I�9X���ӽ��PO���KJ��Z`%�)�oQsQNǈ)]"R�Y;D��f�WB.K
H�����Տ�����|�hR8,��PJ�ɵu���k��,#��-B���!� o L��,�R-�B������3
�1*$�ae1�9JG�J�E����,Tu�e#f���L�S0M���T鮠��X
��u����#���}�)
wR�Z4MK4�I��:�-�5U���*F��9���*�r9��L���Z&���U!!�W�d�u�i]zp��駟vN��e�������a��MS��&UI�lFv�i"E.Z��S0 ��A.�D�^c��,Y�%��Tn�M!M���G�9��6�	��>���o�PȻ{a}�r��/���O������w�=9�ݳ�h��͕gR�7{�g��>�y���{y��{�'��_������y>:{��/A?�?[2��i�i�c��n<�=���������~i	�.��O��c���/�9=rԔ\7^���hg,�A��	V���0Jğ��3� qL�3Ζ���%�m��<T�9O�9����AnG��ꁃf��v8õ!$ר�J������1�(&���eB���ME��P
)%�f=�r:O�J4������KV.+d+�R `K�b�ɚf�6�!2��n��F�U���8���mL�ȇ�G�\��pd�:�L�t鬨iG����BF&Dd4�͐���!�V+>
q�Im,�ϊ�
�Nz�0U/�� �-DVQcA�4�d	F8�	�Dv	!�*ј`�J�	_��IȀS�N��&ޚ�f=�h�p��~��)TK-��! 3Qc� ���(����r!&��ޚ�ar��3d!N`#�*�a�4��9	�(�A�U�i�:D��D(7���t�����q:+�1�� �u�ޚ�n���i�|)ݷ�K�#Z:��*a,�CD�巺QN��,}�[�j�)_�)�)$�~%ИP��G���
4�K��9�ǩ�)�S=8����Q��ʯ�i�Z�M�&k���V�X�V�k�� H/+'5����S`:qt(T-�>�I�*J��#�,�U~%���lE���4U��5��UX�L'U��h��p��|�Pi4Nc[4�KA!
��#0S&��eBpuMk8\"��2�O�>���t�)#� �@8��S0��Z�Dm&(��A�t���O`!c&���j	n�N0��n4ZG��6��֘Ԥخ�Ka��
5�r�p��uU�h�!�����|���@�H�Sݲ�R�*���?�B���Ȑ��>K��A�|���]2?r�هZ�՛6��p��O��-��3�L
�i㐅����X�|Yh�Mri�ϱ`S�G��ϔc-�y�
�W�i:�VH�hZu��<δQ�t�;�����FǬ\���}A���Bnu�P3��O�M��-�LJ��|����d�z�J��F��ʭ[#�84!�κ:�"��h&��.��E�H4�JH�Kg�v��UM+]�����Z쵟�:\�$W�{�J鳘k�]���ě��O?���]�*�2�g6]'�9�lx���b��s���kׇ=Wy�by��.n���.\�������������aۙ�~ ���O������]���w��gQ֊|���@D9�:&n��
���k�|�s����~����y�z�-Ǿ�v�������,���ë㗇G�'^����P��pપ����o�x���f}��v7�>��X����9$mK�N����e��َ,��!$�&QʐzH��d��ۧ��y�~s{G���L:�����P�8M�%�����&KQd8$2�C����*�i���0"BL'����_�t㾹�І�rt"
l!�b�ٌ����ȅ7B��i����U%�ʥP�CN�(��%��3��)G�|�g���e��"Ӣht���ʯn#�E�7
�2[!��6y��l����ۻD�:�ށC�#���,�U�5u�S
!"znQ@4�p~-���(�m��I��!��C
�����CV�~R�d��\T�T4EhD�7�O`) �X!H��hFQ���S����pO|�XJL"�|�~=�+n*T��@��z�̑B�k�ބ!��Α��Dp8_���.pz�7�~��'.gB�~���Vd�z�)�"s2����t�f	i�D��Ek=Φ���fL��PEѶ��=��ˣ��i���%����G.��|-���Gg{�9Z�c}���G�~ͻiO�֡u&�҅�l�z��6q�j݀��}��C�����Ww�{<�޾��{�{ys�����������ե���c�v�~����z]���۲��v[W�86��12�%�o����mN�|�����lL!��m�N���)�w{Y�� ��!ݨ�%;��I�ԅ�Q��YK�,�ZNJ>��h��%^�8M 8@ǿ �+�B�$�o�T�	p���r������p��)�gB8)��Q- �Q&�1��id�(W'@KH�c�1�m��A&�iԆ���7�,��~
�HS��XT�F����)�`���ɭ����pj�~�[5G]cg���1*gj����tKPt����a`�[�ϕ�Ԣ�M��dZ�5��Y�S�t\�r�s*�7&D���}F0�O4
�$���)�Z�SQ)�5L�f94�h@4ↆ\]U4#����E�E��"מ݋zK2�������}�o!r��#�@�>MW@[W�B�cD�h���&���ǜ�S�8:^���rlS�e�m��/銦U�(��������}���>x����ۗ�>����D��yv|�V�͡�W�ŵ7���;;{��;O/^=����]�:��˯�xv~y��{������
����'�����9=x��nx����o�~��K��=yp����������[�"���?�W�-�G~k��>ݴ�}C϶Q�:�u9������˱�v~�p��&�9�slN;&d��?d )L�w>�o��:-��I��V0x�M�2� ӡ�c!)h-
n���rJ���D��MC���ē�,ݘ��2M.�(ė؊�Vk��I�_�Q��A*����YlY���)3��ր)�qn���pLK�#��)*��LQ~�
\JG��	�N'g��ߋI�M>K�Cv�� �|v�6���rD#���R��M#r��kl�qve��愴!
������H�i�%���,�Og�8�K4N
���e�Xi�K�L��c��rJ��Ip��8j#U�9����z�c҇�4����ee�#H�u�R�0����{��䲌J�%[�@�8:��p"�)%��8�E��XV�9R��IX:��h������AZu�r��@v���Lyc�&hK��M�q�YKu�_�G�#B�(lzo�+�iqv������V�~�#5R��4�hW�%6�� 9L����&׏>�R"NHN��9m&��q��H/�g��&�Ƣ����̖\	��H�8�̔_��)��	l�IM����S0
q��B��S��9�|�X��S�+������Jp�3r��S�)Cc���Zr��
�s�j���1��M��E�G�q����E�45V����ȱ�0+4m��HDN6�iݢ��o�ϦM�h�����MW�Ư�3��N�!@X��l!�JA�
�懠���\��4�m�s�֒,�i�����3�:�8uG�4ȧ�D�#�O��|d>����f������YѺ�e|xʵ�|��v�����b�n�7��Բj�ed�L!��sYL�L�Q:�a�i������:�Ά+� m���W�c*Q{E�#����I-�Z����������Sۑ��EG�}�Zj��x�@��zb�ڮT�����P�����n�V�]�\S���7��֎�w���UP���n������;o�=98��Wevt|���]����=w.����~���'}Ǟ�v�i9V�3��n��)�+�.R:�~��3������ov����^ׯj޹���U���-�#%�u�������\�W8�t{ptvu��˙��n��qp�-�w�'�������|�����'��^���M�y^+���.�u^߭oȵol��L���[{�6m��|]��#�j��A4혖ۊ�s���!LԔ`%�^�`�%d��*S(��0��v]��0QV?����p
�lɝ�u�S���T׆̴�#�%Y%�֧�*r��!�N���	qjiC���JoJ7=Ph�~k)��b#m���m�i���YxR�'����Ù\L�`��|�6��fuB|�(͘�q�[E����JIm�JO?dc��V
q|Q�B� s�(~N��8UAppM�/]h�h��G���q�5�5�I�r�M[,�&$���eq�\K�#�X��t�A
m��:Dh��I��j�N���2L2�MG�h�FQS �N鲪55D����m48M"ʭ�[b�ث���Urk&Zj�>��2�r쐵a�*&�˒����y�UQB?��1�
�G��h�"�sT��u�-~�s�u�a��544>BL�)���Q!u9@�V���k�|���'���3���%��'�<xo8���\�1=��L%6��y�w��[��=8�v��H��Ww��a��#���C��m�)-�c�k���=�ݯ����`}�i~���Vd�r�)_n`�!2{_T�h�a9�Ju#Mm�O~��7*��+ڮ���N8�Js���+�ߣ#>��ٲ]MX?���L�̙�yBA3��(��Y06Mz�H�+*��YA������s!隗��h�����W��	i���� U�X�h��BP(�r�2R��>�@��EԱ�e�	ASYF��H᧓����.<��꜈=�+I<H�(&b]�L���3����)к��J��Q]V��K� �iɘYW��4���~R��E�lSzs�π�8v�)�q��MD	�,Ai�8��59#}m�S�h4T��6�9�*��O��԰�J;��8p��M�0��C�L�*f���lk�m߻`\�s��w�w>�Ϭ�V8*f�r��b=+��#�L�B�h
�8����%BXQ���|`��mo��h�+g����:������uAW�[x|V�\G�W��Փ�����;<�ӥ 9���o_}��鳯�>��ً�ó����������}��ӗO�_~qt~��Ƀ�˛o__�?:�yቯ�yv���{�?=�����xr��J/~�O�����xy�΍�?������/��������~���������x���ʯxޭ��Y?Y�]�LKv�J�x�q[Q��jM1-6��d�F��l�D�� N[�1-�Ȥ咵�Yv���>I���X�Mf��4�H��;s�o7����D,6������o�,��%S`:1���1����ǡ�V�'�h7l]�:�U���>�2jt�I>+�����Í1-��j��:��mګ��� 5B�UEo��!����?�4%8M�N��j �+���d͹�,�?Fm�!�M��S"\�V��l�'d��0x!͈2���Jc4>�4#�2YD����ui����gt�N"�D8��*�fd���#Ȓ[Ke����Ɯ5�`̩��VHJ4�r)�aȈ !�3!�thr�)���!)�H�t�FX���$���gkh#H|���Bd�a�����wӮ�rIő����s&7�rm��%!�i:8Á�2S4N)���a��~�)Pn�'RH��U�F��@
�4>�r��/Z3#��P��)�o���-�I��F8��z�C� &Yh#%�÷�n�*�MK�CZG:?$&�r�;�q*��N(��=>��H�qf����J��H%#H�Q��&�ATJ��ݕ��b&hlJ��x='�S!-�Z�r�%��2�b��i,e�B��9F!�(��ZN�z�"3̎/G�=���1+���u�$"(�'�ǧ�)����o�"�|��Z]�����юx�fR����h�}S~-ŏYWF
�eU���L���1��i�a-Ӕ®�ʥc[��\JdR9B�2_�B�����^�sky�̢%H��ӑ�ǩ���B�|��r��sG�lˍ��/�3{�BS4�)
��_bd>2ݭ��z&U��95cD�X�I�M���.4=��%�8��#�_��ҐԌx��c�4K�r�)��Y`U��%����Y4EE�)�p����1�o���I���>d%�L9pR�����_n�ߴ�V�ij4�%4�V�Rt���r����V��ezy�$�Fռ�v]�ܿ�Y�L�%�[?b����$Ǿ��x�3�{s�ח�:�\*���顇�˻�ϫ�>&y��q�UH��к�ȧXm4�墳��]O��><;|�B�����<�;<�LZ�>���\��qK���Ұ��r�X������ˇ7��ѵ>kz�w}�5�}�W�ЮnΟ���G|��\��o]^u��_����G�/}�ҥˮ�y�󕖏��	��K76گ�����vã��7[��6y��m+wn_� E�:oڱp�M�h��cAʹ1B�j�1��M6}!cӘӘF�,�F���ٙ9阻m���@�����	�42��pL�u��S�XE��G�8��L&�q��E�3x�P��g>���Ӵ?F�DG�_!�t���8n�U�)'�Z����MR5S���ְ)��Af���AFB�q� 7��vL!H��h%J�����W�8@&��b���8}k���T�34SQF��DYJ����!}8�H�H��^+*�H����ҘTM������"MC�"�1�,B✖�4��6J���Kh��m�kW	ֆ�δE��$2:x=ӄ�G��'�1|`����c���^�<;�O���B7����k�/���E];��!�G��g}�uGN�JҌ�=�f�up��+�	�[@�rB,O.�NkE3�&)S�|�z���ӡ�W.9�_{�9�{ts����j�>�x������w?8�H���eFGU����6�8[�͝���.V����ýv�꙯^���w.���~#?�����Ҏ�m𛝎�Emg��ݥ�s_��/X�-�c��]��"�q�\���9e['nZ	��^Ga�|�:)�,P�3�#N���^.�!�Fv�pt4:���:�o_=��┢7�>j���ҩa8߈,��2E[c��"���d!�]��X�S=���#��A��u�+)� �O��C�/��i�d1�� `�q��kƉ��/����W��F{[W�47B䒕�@��r0#�TŊ�H\V�׶�$�A��@��,~G!)jmֱ�!��Q(�P}JG��Q��n���=����r���h)AR�C��[#P'��t��X ����.B���lm�9��~�J�EPHH�)\m�Ƙ��7 �����ט��$���l]�M�	�]���72�޺bT�=�V��O��C'�\��h��v�*�s�n�&������@��9đ8L�M��eMu>~d��q����у�%���B��@S~۫��[[aC�N_M�����/|S�_��_]^����v���o<S��|�����������{�����g�_|�͗�^_����'��;=��~��/~�|��7}��z����������wO�>=ܿ�����O�O�N^���������|����>z���<�����^��W�����ի/_�<�98�t���w��/���@=���������unXk����    IDAT'���(x�#j�� �R���i 丈
1SYpg��B�6�6B�a��* ����R�h�cAVRF�I��Ç��џ��⢘q��0��̧�o�ǌV-L��z��j��|=�� ��2޼kb�P[Q�	N�������F9�Pە���t��Y:F�����a8�zN
?AQ��C�联�r�1!�ES+��k/N��@V�L!	�!N{龅Äb�I�B�9���3�i���h!�M�a[��)G��i�zY���ਫz�4����-�4ǘ�Q?r����1���/d9#L�h
-$<c;Ly�ьl���U����~��g8�V'��ЀB���Y�zk!:�i?��!�Ur�t6�y��D�X��.Sh�p����Y'!B)���r#��V��1��b�'��p(gZ?
|g#�ӄ��0�T�*���D�	��:�ә�),E��ҡ��{t��F�6R��#��Y���'�i>'�RD9�a���4����y�ӯQ���[ʦ��V1�84e��I�4���6�D�U(2���O!_�4�_�n9��L��#�(�t��p#7��}#^X�gʉ��,���SN�\���dVnY���Ȝ�ڷj	%^��LP�"�R:��L-��&e���ai�SƄp�Ҁfd�0g�Xk�B(_>���YK��x+�3N)�9R��ֿDVKh�%�O!H:Urj 2q�OA2�B	˝i�j����r=#$;�1-=�Q�#خ�?dh�uQw1�LE#�X������8���Oj�oF���o�u�$�NW�#$��S�"=�>d�*T�)'N�a���G��!�!�L��D��(��)�JgWʘ�s||!��G�nw���3��j�X�4U���,��3;���5���\V��	'�F4�k�9)ش�M�eYm-�rQj�%���¤�tJǇ�	��[���(�u�ܺԽv`��G��������1��{��k��ZG�R����u�_X�a|�2��➋�{�|���륮zz6{wsr��+u��~̋ƞ��g~��b��/��<����3ݻ�<<=9}�{��ˊw�Gj�hyp���Љ��]g��:+�gA���%���>��+s�ނdn_�{z���+��c������8�>jj?n]��c?
����|��嫻�۽�G�w��n��t����\��y�E`�.�Z�m���8�U�Z�w��p��Y��q�fW�t�9�B�������T��IY4�\�|��
�ጲQV=��D�����b|Q�N*=L��S"*1eqTw��Ghȣ�[+MjI5&.Q9�%�is�d�mlm�ړ�Տq49����o;
�0��C�뇃Y!jU�b���i8>���1bʭP�| ?\-�5�b�M����|NS"|E	�z(To���Z8�|}����FJ��5)��zKS4N��^D5R��`
�s�W�b�,� ^Kr�
%+�z�Dۅ����^��qH�RW�5O�Su�1 �(fEc" �j���JC�Y"��E�H�x|���C�n�	�r�lD��7�Rfj��t�Z-![TVb��@>G����hR�C\{�KԴ���%Z�#�2�X��>�U�&�?��~��!��'�O?���/��)Ϳ�˿\���"�W��c*��Q�L犒Z�J:	�h�J��n��B�-�T̚F`�������l��5@���x;����Ƀ�㳻�'�gO���.��W����N��ۿ�o�[���c�(�4/2?������z���cqs�>S�����	z�?^oDr2:��,Ԃ���ͽy-��w���ND!��%��fCD�#Cڴ�E1��4�І�[���8�w)��|7��׳�U�wΙ:��c�:_�>�1"�1�U4d
��L�t8R�F�R�5,�\�X��&�R�A7������P-M�Z%N�Z�Ԅ�C��˅��Z���q��d��nM݈R*j�[)6��u!�N�"Zo��.�d4��j�r�u�:�8�E���>N_���F �xi�F
�|�9!jQ�?���M�%�`�A�8^?���\�����{'�M��\
h��CP�M�U�[��,|dN�Ϻ����'�-��(D!���򫘚Q�@|�3m	@�����̮���K��Y4�\��5w��hRVBE��g�T�{���?���;Db�ҭ�){?Y4��Q}�L�J��ऴԘ7��9���M�+�	��,=�g*w��%�/*+��8����8v�θ�'ݵL�P��1r�x�ܵ����N�埯o�M���}p��������~���O_}��˯��{���ˋ�g{������#ߣ��җ���>z������֏����<�y��WW�/�n�<�������^=��Ϟ囃������?��������{��O�>��O~|���'?������+�7w�S�g~�dm{˴d�b��Y#3�;�6g�|)�(t�l����Ԯv�]��Q�B�1�^��{qD�d~kBL����:R��� э����>�#��!k�P�n>
t� *��c��� B�zSŔBK��7�L�t�:�Gm=�@L�̧I��p
�q~g2�Cq��%�D'��Ɣ4�i�$KA��?+�|��E͘l�&���u5b2��@�d����J׮m;_���� �H�@�9��JQHm	Ƅp F`>)!�L.ܔcs�8�5#E����0x��MG��_J��M���;�%�k�t��#R4~��q:p���Z���A4�7�s|R�V���5��q$6����:p)��୺�fz�IsWV.��3�SN��	i�ƄRS�CDJ|#�D�B$Y�@Y|��iL�dD��}�P: �����|)%�sк�b���M1KO�Z�B�Y-��&�V�l��	���I�lm��
qXg#����&��I!2\:���4�n�8I�.�D��[u��Uh�$�����F\�T[7���L�S.��d99gv�uh��π�F���,8ek�%`&���v�r�FS�@N}
�NUL�"�\:0��)�Mh��
l�d�ќ6��T���F؄�1kC4���ġ����P���e*�b�'�����#Ǵ��c-�<N�v�����nE�id��h��L�q��_�+�Zd��̝� �F.T�|������'�o
b��ӬJ�˂[�є��r�րhx�FL`Q�Y�,��ajI���OP֜u��1[�)+qz�h�3�0�+���B��q���,Sd#����IG�`ҩ�Ŏ&8��L������d�P(���M�+:�D�F���o!�TMȉ��O�� ��pLc��Hj1��Y�D�0|� �t4K�gU�3?�}�������PR��L����N��6L�;���1"���C�k���4uŤ�:��9�h���GHPn�����Nց�:��l�Ȳ��P�N��k�Qz��2g!���˘�1O������>�c]��Ķ�&�s��E�� �7����HJ��FXi��~��f߷�z1um����b(�5�u5�τ��"��������ٵó���]=z|�wd�N��OO�5���9&~{yq�w��n�*��=��#�
��?$�f�;�����L��k���|�G����^_Y��<�"���=}u��������/^�^\�X������'A.��+�b��.�M�Mx��ەRem�v�_o56}�B�Z�=L�nk�������Ul|H��P:�+Gӆ8����h�DQgh@��@��pӚ���G��QH�����$��*S�+���(+���:���oCd�Yuf
g�U �1�C��t����(&��9Y1���>\�J����h΄Lu8��4��Ϫ�:���B��B�A�u��MQ!V?���d�n���5gB���݊#>�8��H_!8������V�Be�jL��0�h ���5Yoh�EK'��1g�<H�2)H��CGJ�N�p<���h9ZB�O��ȩ�5c��y�k-YzY��ј��g@"8����@#>��F\�p)�sjIۤ�3�^��sq0M�Ƨ�o�&��ʹ��n��=��h�W_}�1Z3�����ӟ��_��/~�5],��O����l�Ȗ@[���%S6]�]�8h��8
+_E[�nZ���N&�Y@S���)��d�j��+5t�|�{��������Ë��>s��<>rA���ؚ�7���}�E������ݫ�w�8Џ�yے{��{��c�z�v�:�S�Զ����_ݰŷosWڙӾ-��8�&����^!�v�h�	9�;(E�6ʘ��!��o~c3�ҝ�B��Fjkv
�y��9����:G�� 1��8��	�e@:|'@�����0N��;%��HN6��UH�cvsR]!��U�v�b-h�p�h�K�g�!��SQ�1��$N�� u�o4*�r���I��S�$eS�L=3;/���k�E�	I��"e|S4#C��Q.e�;�">��A��hi*)n�)D
Id�LHn����F�U4#���i���2��O'�� ְrBpL:u¯.����c"����J���%�Q0"��Y����Y~dd��4UQB��9��K��D���UA7u�%vճ%��ջ?��?��f]���b�L��7�u�`*��M+JM:�p�:�zz{ܑ�L�L��޺TGcB9!3�^jFS��f~xH��p>pz���QT�&�:��������Ï>��y��r�m|���������\|��_����Ͼy�������=�$̓��G���>�y��6��Ύ�ݣ�)o�o��<|p��������~�ū�מ�s����^^��/��$����ۻ�������;?:��?�����?��/n���֛�i���������-fVj!��;X�aB�l�,&$�mٖ���+��Ɓ��i���1��!��BN�n}�_�Zi3���Po�9�lZ������f�D��Jc�Q�tD���W��|�Js ��J�.��`�FfC���\j����&�6� �@�����328�i��n��vC�ȖeDf��[�&���L��MV��>r�EUL-��T����M��"D��s��U��!�X
�U)dJ�_Jnj�N	]�4���ćH'n��q��)�G�)ZJKeuX3h�z7��G`�d�>�3Q�D�էuU+�e�"�4N��n󉓅��4Dn�c�ƭ��^�42�p��4GW����O�t4P�B�U1�f~+**��gn/��5;B0��OS�#�i�����[)��q��lB�R&ĩ(_'�,�t~S�(�f� �t���X4�݋�>P������߃cu�C$�3��!���*W��p[���M��d1 �iWCL��ΞX��nl2o�PQ��l՘�Fd�8�ő��z@й�i�c���H Zd8��� ��Bm!}�3->���2
���ME��Ǵ�%j#D�rC�ŧƄ�s�\ro�8Ghd���?=���k��:�T�_T��8VnRE��a2 �����&����!]���G�Ϫ���ѱ�I��"���O�X�ǘQ@��djq ��)�W+�"�jl
|8�cZ����U�bYE�3�8!�d��8C�k*T?S��X�v�>Aʤ�2j�dqМ6��4~��rp�7*o��(�ZM�%!¯�֢ad��MѪ��r�����hd�W���e�(�a�DL+�^��h1�6�)��m����Ҫ�/��LG���Ɯg*��%��c)��PѤ������В�R��3Y����|Ձ���2���n{vӱ��˝���LY���B�P�۪@��el6���E�2�!�SoE�:���M"���v�g���ʾm�짟~�7V �֏(��1U�����]Ĥ*�K�Rl����>�᝴���y��v}}�Ihur�>�i���ۛ�_f��mȑtw��]q�sQ��Ϛ�^Z�(뒩ٛ3s���{����;�o�}���^N==:��M�>9m���O[�_�\�e]���ߢ����������:��*�=I������Oq��^���z�{{�C;�'�.=��{��t���]<=���޷/����zmx	__�^�I�[_���g����c���������{��k��C;Ϝ�F���̔�DR(�t�s���Y)Z�Z�V�$�t�M�R^��
�MGE��rjF��Gٽ��v]y~�G��x�h�H�%��BK�j�F�m�=�ax���9��xj���(���rYZe�D�"yof�|Ed�?�|�nEQt-����[��[k�s""#N�I�|�Q��ٛ�#�!�t��B�pkL������JбU�,Әxm׌,8&é�qL�fc�pS� � ���P"�)�8!��JD�I���0QӤp:�8r����hS��@���m�U,��U1�j�I�4Aե4IJ"5���O�)��*MI��p+�&�Ŝ�I)��hB�fk�"�C�Y	2�)�a>��f
G�AP}r�K�_Ы[�l.�/�h�UI߇��l{�ħ��i�3�5L\�t��B�u� ]�$�)�5L82C"T"�ϱՑՒ�IS)F�f��!�0i�5�a�]jd
�%bz�w!��dS��A���������39b�����1S>��M9��e�(��:h-���K� �ٖ��X�!�?�}�ʞX������~��[<7;����~��n��QUq�{��Us���o��˷e,p��to|��6�HX�&�=8nI� �d�:�7�{���D�z�r�Y�G#B��i1���4aɁ��p�����&�LGW�_�d񁎷E~�i����e)U��8��qiSE���后�L�og����| r�N#��Q{K�ȚEmMS��%��B�5Γ;)�@�6�E
�K�ԕ3.W����k����V�������Z9�z�� �1�!�������$.Jօ"����B��@���5�ST	`dka�=֭(2B
e; 
�&�*�[E`��V�J�����B�E�0U��ᘜ��BK�ޜ��|��gK!�ijQ�LE�kX
�:��"��=5����1�4>�VD��0�B�z�aL e��ez�kE�(&�����Nڬ�AJ�yBJW�������|���ln�Gy�F�#�ߣ޷9}7���~�3�B0��T�FH~j��a��V�hiq��h�����7�F�pjE�M��#��J��E{��dK#H�i�wy��� �o�<}�س�ӧo��yq�����O]��ݧw��>������>�֓�C�Y�K�k]s�}��v�/gxw��{�5r�����9Z=�p��K��<}z�O��p|�y�"���g����ǗW���g����휽�8�����ӫ������O7��fu��M���{�=~�]�S}\��iuv����h����
!��m1���uv��� ��m�=�ؙܲ� 1JAá8��јG�(DE̔�Zէ!��6���Д�ऀ#�U�)B��	J!Ҷ��M�'��cT�n@&(���?;�W�Tk4��v.$���,��r�Q�����R"N%�~�*L��Ѥ`��_J�&�e��Tݱs���)�¡�ɇO�lF4M��9��I�&k�M��6N=�%�g�׆)+�#H9ߔo�O�sC�XO�Rh��VbN9�h��8�j���h)	V� 'NG�t*k�eѬ��$b*����7ȗ�!Ԁ�SR�����DNx���OGHE�tƟ"�0��od�|YL��,=ˊoD�G.�ɏ\4�8)d
�4C�g�tL��t4�����CK��C����S��U1[`"�A��1�_���^��Ӊ������a�~����1�8��4�ҥ@�C�P�U�6�pjM��@�H��փ���[Q �����4����q8�y(����LXi~�j�ʕ[�<�Y���b�S�=U85,g*��aLR3ĩI����c:K����[Z��M�9��h@V��%S4u!��9g$A�M�iV����	r�2Y&�l|���$Ri:m_H�����%�a��)@=�ʪ����pR�E��T�Y��:v-B���p��*$r��d+��3qҀm�[�\�F&J����0%kT4�6$���%�	�"�S�|#bp��B��I7���B��4�L��!$h�^W)��3�рƩ	�<��3O�R,?�X�t    IDAT�rB1SkNS(_
K�ou�O����84�֦B�,��@K��h�D洢��;�3e:1K�n�Y'�8��Ϧ6J{F!�@V�,�	!�|LY��p!|#�� �2!Fm>O�L�T�f�yu���E�rqD�-z�1��0��Z��FY�l���x��n=D�4�d���z��#���B5�3�R ���_�'��(��*mD3B����w��l(���Y��e�v�}�Х��Ա/��}�� �:��y�#��f����zumt�ߵ�xJ�'�2l��0����k&�}O7nD{u{�����㧯�q���{��;ބzg���W��z�����໾��c<T5�Z�#2�7�J��ri�R}a�{������E�(_�q!t}s�Yف����f�wr��2�����_�}�ʻ����W޳o|һwv��~�n�n�rsw��v�ڻ�C�on�xQ���}�{�e��Zꁃ�z��%��l��q������7¥K����& �� ��A��&���B�Hs����G�"9�r�)�V���j�DU�Vc�heq�kFȔ��t��F�X'AN��"s�t�gQ���SQ�B��`Zo�|�M�՚]͔�FdcV���D��!�<�j�(�r�6��fc�%2ۛ%�E�v�B�{J��d���$R��L�&ì\!�j�'�Y!Fu���Q���_J���DLL���V�1gK��Z|��hΗH�������6-7����8�8�.���yY^D��zJ�A�t��I,�\�ƞ|���I��Y�UT�%H���Dh
�P�(�������o�9h�
�z�̊��
ߢL�쫙ݘP��.�S������?��/~�|Q����o�ە��k�>��A2��B[�:}X�fgR��YjV���a҅:�4]��Q���c���`�]%�A�/��d����ow�����wW�\"4��^do�߼��������C�uʻ�e�k.ہq��g��<��N�=V�N�jx�_^��s�@�Gh��v��e��Q�B���ȇ$ˇ��9p'\�W�\qy�_cq��p:w�
!��;"B�h��Bh�`H�C?YU�u��:�`�O��%pd!w���3D"#Y�GW���!8��F5��LQϹRB����M�(���	����XQQ%t�Q�Cb�ll+l�u���I	�ǧI�#d��v�XH�	tA�m/D�&��J�rЊ�a�d��g�RjLYSENdc}�l�z�P6bF��)J��BH�^:.�A�1��.d4׫ 4�;v����֭+y����<�N�J���&R��*]ź��.iU��֛g^�|c�H���2!��8X�@)�%��_��v��zZ�M_����MG��T��WZ�Rj�\��9�I�J��D�Y�UG�I�>9Iea��Bh�"����e��9�֩J��
-�/�:�j�E�3N!�	��,��o^:������?��vn��ݗ/�N/�9ݼ:���W/^�w=VO�繼���������ʶ�=:x6���u�ٛ��K�����ˣ����ݓG��O�����8|��W���>�����n����g�ݓա����7���g�?�/��7�����?�/���?�:?:~�s���Ѽ��h2G�ч����+mv88v ��6w�M3:��1jN$�BM:ăbno���D-\hJ�rU�3�0N�B8���ˣ����B@����(-#k�4V-�R��E�_H�t`j9|`�q��%B�cZ�(�Ҕ�@
�N��!�j�,��0EƜ[ڊ 8�Й��`Z�r�M20�L��T(RQ�E��Í��Sx-���}L�E�h9u�G�+�Ё��A�r�n��%"��F�3��ULq-����=�ۙ)ԀiN�%H�)K��1\9����V�cZ"�!��3
!��$��>SюѤ!3!��40V.pi��p�!_"YR|dY��6RW�zBș4SL�E!��9[�D���81CJL�D��l�pD�.�i2N�3"Ũ������В��*���Q:�$��%�����*�/���a��7�2F�D3�S��g-P
�� [��S�D�RH"P����Õ@K0Q1���h5�6W�Ɂc2S�i��L�u<|ů(&�ʭ.~�/*�Q�3~�f�Mg9��An4�@>�~L�쇏�Dq����g��cj��p�[K��%V�hi�;4�l�,)�S�q�"V�����b~!�֤FN�ϩ�p#~8�'�G���CH �Y7$���j���
AR�5�(�B�&��7!��)�h-�!f�3|Q��ķ��R�q�g���+��2ͩ��	�)j��rI��2�"S4#�6� �mB7͙�D�?P"���I����Mͦ������&�P
Z�&Wt)8*:�vOTQ r�8�zh�?q�5�_o��pBp�C
��B���ē�c�� ��A�t~Ӑ���#�V�2��+4	�DD�\c����?��C�_��t�5��0����AR��eJ�an�7��y���MB4麭=�tYE�~����!�6�Oǘ�oLG.���8�!�Y�ĨO����=�a�����E�Z�G!�J�[��Ȝ��{�ɵd��reE3N_�ӗ+Dp(/PKh����h�����ʺJ������9^D$�}c�S4�w̾[���F���������(�r&���Q��w�������X����}���|��G���cws���fu��{v~�:v�W_�	����;:X���o�(�£������WQ��q,j�Z>�.)-[;�7�7n�5�=zt}�ʤ������;���yy�{���`���������� 4@˿������� ��G�.�Z��m�4p��� m�<|Z�h����V�~.�9�\j��I�~w���P����|�-Y/�(QK�4�h=�q~���x)�0�)!h�W�>��V�1��:��\F~`K�P���h��22[dDf|#�\��E���͟{%J�q���Rʂ��ګ
dZ:�=���ҧ���JTH�4X=s�-H*��h!H�-><e!��?i�R@�H�/��j5��>A�"����IH�ɩ
�Z�QNú���)�V�YR�*ڱ3M�>� )t�p��R��R�x�)E38M>��2�5��᳖�Po����O��b�X9dL>ÙYV1}8CH�K�=ۘ�K8z���Lq�8PB|x]U����{
RWTHQ���B���F�����q�$����\��X����a�w">�W�q�r�K�|��:�D��d[�W��h�Qnk*�ִ\cn�r4a�nT��p7��6�i���=�v�n�n��������멿���us����GoȐ�j�>���􏱑�eQ��+1ڦ���ݟ���=9r��b�`�ǯ��N�x�{2����Z�`�_X��Ɉn��a�m�<���b!��gj��q�U�D6a�.j���O��5�V?�BV?�9���|"��Q�c��c�L���M��3��5��t����mJ��<V�A��@UE|�B�g�
��u2�un�+�hZ�%!pՅJ�kipS&��
�I�O9Yk�"d�(D�_���e�JWT�3��A:5��)��	|d���s0;^ESӒ,��0��:�%b���B�R��_v�&#��)T�s�B8]i#B��&�=G�YFd!q&�$�&NL�D
�F_]&:�#]ER�%�W�"����g��[]c�����B#t��R:G.e�k��iM�`ʵ
���Q�^#��T��ό|�O��nD��=Ԍ�ZU�%n�|'�9����I���jAtR��uK�)�!����4Z�6^�p�D�f�m�Ϣ�%�7�A�FN�B.j��kim,��a��ۻ�����啿�yy����mM��t-s�/'�6'��ij�~}u�Oi�o���8Eo��[�_l�����<~�����б�����O��O�y�뫋˳���ȶ����懷?�8_}��O?>{u��������w�������_������GO_�����.�~�W���Y��e(D~<�JǮ%�R��E�l�l��$�p2�Ұ-�Zo��^L�4cZ)e��t���):q|fJY��y��k,�V�����Af���(�#E�;�KL��ėǔ�!��9�(�a"p�sK�;i1�`#���Ja9D��Ę|:覎]����׭��sjX�$l�3��c�����CL�oli�J�t���[M#+��k8���q�� �3H������V�z���϶��E����:���р�[0Kjd.�5���ۥ�0��>2f
8�'��`�����r���I*�ΐ��!^�*����rD��d�Ф!�3�۴y"�tf-d ���P�uۢDq�E���ʕ�`�(�>xȴ�goR(���cD�SK�4�x\@�e	�(�N�BD8�,�C3Y>�Z����#�0Cx`j��V��E�A�?q�9)���	����P㔂S���fuK���~�.�����G2e�A�G�j���is�)O���c�n��Br+m��$(]�r�j�#L�t����*�"���������Ư1cNG�9�4����(�2p�SU��fV��t�e��D�e$�����L�VdZzY)7
��.�2��(��28K?M!����MBj��3����b�p hR9B�����1N�8�m��9�o'n�'�C�b)��Ԁ8l�Ijm��1Z
1���Cbά)a������Ǆ����e��c��n�M�9r���-rN:U�n_�3�R�B��|�j{�9�v�t
��8�Z�\�޶��-��+M� N]!��ɚ�sZg6nd�&A�l��f�k��F4��k���%Ro��� �*����|c���̬�#4��a�Y!c�F#��B�+A4�(jE�*��%n���1�Z�fW	�i�6ֻ�~%:�����S?IiU:��Ao=�eq���TaS�)T8��7�	鍔*݋ˇ��4N�\�1SdNYBD�r+'d���R��d���a䔍r�ֈY��K�����4-�G���������X�De��aE;��8w�)t�F�/��R��a�|��M�J��Į|�r��7��6��e��S������_�|�s|�r�зR\���zsyv�{#G{h�|��2�݇�.�Z�x���ӝ;��;}*�/���N-��d��v\����q9><��,?��\��ܙ�1���ç���Û[�����@�q��W׃}kfy1��	�/�<<�eEm5��ll�c��%q���C�Z{!�Q����̵
��4��HV� 5>�ybZ'e	�%�D��M���~��L�Q��� !�S�9S�ɯs>��^�@�B�No�����-�/:�� S��o�q �Jh	��2{4q�AHJ;��޶�7�̧���_K�|��ji���*"sf���j���[��5f���S�-�BB3�Ϫ�6��(W��#���j��b������L:�qz2�����"1�WH�4>��8��`��'���4ҙ=7%����a�8%p�9���Y�L7�~�L�gl~R6��i[����B�ͷk1�i�G���j�VARo�(T:��1U�4_:f�+�ʚ���,�ZF� �yx��MY`Y-���\#Aw��A&��r~����{|��*��L����wm�g	�ʗ~>��#w(�����Zu<�Ӧ��.p����|82�+P�|��0>p���9��h9����~��]���__�:;}u���^���j�������l�k�^���}x��ϲ��V��핻1�0��ً�ή/�ѝg�d���a�|#t9�\Zg�ÿ�]A���40:_�Bl���^�Mk�ڨB�16����eO�_z�՞7B��O�ʙ
!(�e�蟎ukt������+?>:R�p�
Y��Ĝ���S-M�4��?[�q;�1�]����ϙ��<w�����;��\mGnRkK�
�6�C]�m�1��4�(Q��lӪh묋�b�ц���� �([��EF��#�[�j��pc��7Z��4q��ogt��(�(��sj�TT���B!V-���X]?�K�L?��V	��b����)���F�VM	�l�����L֓]{���ɱ�Kۢ�bL-A�B��QVE�@�#s�:l׌#R�8�-jv�\)@>N����-�u���O����U:R�#���G?2��}���&Z��os���#ŷK� h#�!��)�`�z���
M�K4�<_K
��p>��oj�|����)e������]*��8�ײw�y�kُ�c��ư���Wvu<\<���#��
�ev������v�d���p��� �e�q��������`�A���v�!�_�}�������x��w��\z�z����<�ϼq=��#�Ν�&�y����
ݜ�嗫˯���w�o~�{���������������w��;o����/}s�;�����wF�y�d����ʺ4c[�CL;���X,�b�����k�6�i%�e����;օ Zr�9����ʈ頋";U��L�h�2�I�f�+�Ə'Pt򅔛��,4�:�D�j�yBbʵ.�����%�6���f]��0�"�ǔ˪^c�8�s�fY�\{H
�M��#�q��2!Ɓ�(S��ُ_�%i���i.��L!�Pˏ@�)D�N��6�H|N���$J1&�V�t��d���ּ�p,�rd#��ӈ��?��!�0 tL�5�	Qb"�č�K��4|TZJ;�3�l��D�hK�� ���B�U����� �E�*K3jJи�� �� �)�i��Tk���9�[��P@`p~&�95 ]W����1k��9P]�^�|VQ)��z'�ж�(��F:e�'r�n�[#��.K�_�<�)�P��k��@~u�s��g��iu�t~�E)��)S�_�5�_Xj9���DPX]xRS�u��|��1!��P�Ɖ��-���!�r��B��)�s��X"�)B?B_�={�h�m��Xu]��v�_�6S
~OD�pY����KdmL��
��w�/D�ê.�ߢ83��u�4L�>M�d+a,����S�@���,MHSN���Jwhl�TC(KJ�����1�i��+TȘ�B�AL�!�C�^c��Q����W���N��ȶ��S݊�PH
��0MN媅�B��M'b��B8DZ�K�75NG�y���+E[��=tr"��^k��sX% MU�":����S'3D�U��Yn���0��nEN���I��w��0ʲv~j�C�ъ
ID���'^(�ij�)d�(J��3�*���hXz��|颜��0D�cMFk�uU��8,}��l[�?A�K�S!Y�b�B��ûi��S�ё+o��|)U�L?�PQ�o7h�!om��1z_�T�JWE
�(_E�4e�-�W��o"���;�4\��S�O��潳V�{v�pF�U��Y.�J��1� 3�5�[�|%ꭢ�:D�7U��� ���"�,���N0������}Y���.�V����ۃվ�]�k�_�t����C'In�c�M���[�Ҹ����G�����;�.���닛���O����z�W Vw;�?�:��+�KsޤS�#Y�H*���=�}?t9-}���X�FE�ƪ}C�{�aˇZ�ׅ�=���z}�7��so�{�����.n�=z�d������`go������
u��n_�vt<����r6i��
��KҖ���,HS[�N艹!D���U�Z!��5�L��_�3V�ZJ�'%Q&�$ƟS
����*���&��,a�B$���z�5�|:�`����"�I�4��Ԓi��e�1�#Kh�[N-�Z��f�pLe�8-A��4��@>��Q��E���`�@!�X"f�����%�i�:4���*��>�Y��pȨ)77��ZEm�,E�N! ��VQE�������h{�AH�S��ٞ��v|�X�:���P-���@&Ӟ���7d�r(dU��#7E�� �O�V��r�IU���L�l��j]^�L� H;L
R-���AW%֡(�^u�4%ʪ��������5��NiS4#�e��9�����[|>�*>���q�E;�k������@��W�W?��O~��_��w��>��0EZ��{B�Ϊ��8i�V,���%�    IDAT��C掘v�)��j��[ N!%�$����վ׿���BƁ[�ovW�3cߩ�˧�{;�����/q���H�����~;ȕM��1v�����=y㟜��ݤa��{{''�����{���q���.t����)皧_s��Үf�X�a�A�x��@��k�JC,�55"l�� $�QJ�t��7�䓚d�䆧,��p�v������p����CL��>�䓮� Eֹ��X���S�B�T�:|�2ђqT]����3
q<Z������#'"Uc�;�!|!�8p�"@2~]UB�&�D�.*���C���pLƧ�� �Y�GY�_n�1��P%j`�0���kw�Bu�׆ܙ�Ú��ǯ>B��Ѐm�r�|{�/�����dR�
%"(!ݔ����j��4�-���Ʀ�l�D�?��R��*pW���$kO�`L_Ed~E���A���o��x|�)�Ƥq�4�#���E�u¡�()V	d����p�{*�^H
>D�u!P�կ~��=���
�Ð�֫+��3�F����[o}����!�F)LJ��e��Ն��IQ�8AM�ȚQd`�#�������I�t69�����C,�i����+��y~z����������啧���^�>=99��0o�O﯎���㷤�VG�+o®�n|u�:>�y�ԯ8�s�o���:���?y|�����w�{�����7p�_����ӗg��<{~|����G��ŕ_)���8�w���W�����/����ǧ����~�ۃ��_��/�<��:�?�����[{=�F��,�6�^�����v�)a����
��f[�x�u��s/r�od%���J��cg����&UDJm@Tg�P�ࢦ�*h���C���+'f"r�PcxR�(�<S�B�37J�Z��&5C��B�H0P��E`���ڴ�JG�n�_J��!�BF�F|c�𙊦@�zB�f$h̦��r
�p"�d���آ�hF�h�0eI���($AS%4Yh{7��:�gv;)-?����QX-�jA�em�E��I��[��B|8�$bF��$2D(qkO�D+��a�o?)�=QOMS
z�ԃ'm)���0�)�����Y�D)����8�EK��L�6��M��N�Γ��*T->#ճ?2�[�Ŵ�L����n�T���26�Ǵ�%v�bZ��3�>Z�F�Z(�:(S�m�G�6�Q��X�F�r���b��#i�9tjU�\\c�\���O����DЀ�)"Ŵ�:���J�ʹBY�@�5��Z���1!F�6|�PQ��Ӈϵ�0m�&fMr��jlZ�J�%�Y��Z�=��9z9�&3E� �L�!5͔C*q#-qk�B�ϙM�+�� -[	�n]t��e�i��e����T~��M.�h�)niFVT.���ƺʯ�i|��)�<A�,�3kqZH�_s^�D����ֺ��uEK-���c:RDS6�w2�@�R�)��8|����o�񑕃7�	5��iR*��E+�x
���0ѦF��B��
e|%�@��L�"K�8	%�����3�#$��[%�D]�J�YB��i��*|[ǙR��G�d�����4ZN=�9F`xʘ)�EU���l2�����Bi6�l-�,Q��q�\'���_�yΔ��ѳ}m�M��*-"�Ԓ�F��N��L�Y��:R��L�#˛b�~��n�չ�h�����4�+%5N�iujŤVWF*��L7��.�h/�`��U�l
��Y��q�Dq��ϐ��$�2>�[�[���oFz<�2!���9w6ͣ~ܒn|��~����k�Num��>]�W5W��v�;�`�;�.�hu���~|v���Ͻ�#��r5��M����M�h���x|���\�^]\?�7=}�z�������WO�ί���+����[�6����yw�d�[�{k���򸵭/�,OY�Sz,i�w˕3�R�z�������9����Ƈ��j�?s��'���./�.wVoy�r�Y��������ߍ[ߎo��)yw�|��[���ˑ2vd9�{�m��u���j�/�������i��s|���r�y(�ٶ��EV��?��뇏`�TxE�Hʦ�і�ƙ`Z���Z�3��ɀ�,r~%����g��|����i�NhJ4ń�~hVZW�z(+���Y�*dT�(��H?H�Bғj��A0�T�a��1��~��Ī�Jʔ_nR�A(�����cm���hB����i��B��`2 �`�8FE!՝j���D0:=视)���A�p�|�10Ǩ�Nl>K�S%��)0�Ӑ�UW퉐\S�B:1�.��P�G+R���-����o�d���D6{�Rhl�-8�՜�|&�rh�&���D�Jћ~������m8��#�kDN!�i%Jtt8v�`E&�l��=�˕�c
�X�����bQW�O&}0�sl��Nܧِ�����ۿ�[�4���)v��I�D�"�߳�p`��ǡo���tLEM�����q@�i�Y�Wn7p���H��_H:�?x�����g��<y�����ro���:j�J���1����<J*���`������O>������{�_����o^|������������WG����ڭ5��W5O^/��a/���Q����}��3v�˭�
M-������jC���02���F��� G)+fȢ1����m_`r�qft���H1��J;��⺦D����3�S�r3��j8e|Y
y>�ą{ن��7��M�~PC����sf-Q)�F�l������c#�r�$K%J��}���<",-bԕ%HI��(��|%��EV()��&_���P#۞��C"�B��d���n�R�R諈ƧV'� B�B�5�H�壅֒SG���Chj�fAK�4ͩ,�F�uRzN\ԥ)dO5H�3Z7_�m���Hi X]�(�� e!���Vjڊd�֪�=�&M�3�,���_�z@�%_�J�d�9hc���$�n��|6�"��4q�J+ߊ<���/���-���b�=��;=��G?�l�
1�V���J#���#E���<�)'m-��_�|]Eh,%5���/�N\��|x�S���+�X�h7W���|���ށ�>��Gđ��"�v�M��yg2^YTF�] <h{K�wj��>;~r���'������do������'o_�~u����˗�����//n�N�9Z�^^��G�_�t۞�ۋ����ۗ/^~x����8����Z���
����n������ŋ�w��ooW�,^~�/1cW]s���`�[�U�o���u�%(�r,ʹ�Ϗ�d �6�*�Z�8��!���5v,�fN'��i�2^�V�[����mK�WH��*��jq"��m��ݿ��+�`c�h�%�ꭅ�&U�����(���T��t�H�mEp�i��7���gh�>$Z��a�
G4B
9ja�r�:(��ګ���Ԓ�O
B��%��1e�|�F���= �ƨ�AȘg��5�9���;.�O
b	��(�*�B�ӈ	L��1�Oa����Öv��ƤD������r��p���G�����
UѴ�;c�Es	S���l��4ƙ�h���\��&�:�a�!p�)���1�YZj]�Ԟѫ��9r�DS�T�%%�l���-VH�)�7���T� ��9�0Ѫ9���6f�j�����E���i0Mc���c��x�R"fKv��HS.NK���L�(7�1c���f�)U��L{�ńPN�BP�@~K+Z�@|x|c��|Δ�j���吪�Z�@�����$����ڳ(�D�r+Am��r�K���JCD�4�e���h�m�"T.夌3�F����̰��1��!�j eSQ�R��0;I_��:�><q#�j#�PK9��9~�m�8�h%C�Ed�ҏ������M��ʚ¥�%�!(�HNe4�Nr���*����X"N%LK�	L�09�KP(}Y�eEk�'�h�*�{���SE�>C��P
�c���Ҝڋ`J��Փ<|~x�Hp*�3m�ܮb*���̪�V�9\zuD%��M��|�'h�,G��E����9'e#D�hu�u�8��8��/�l�R3Bp���ǔ)TE�d��F���/
/j*�D��m`��5e8�e�����1��!�89S��+/��ړ��� s�2����'rL:I��7J�/%�tG�(��BH?�*�b̀v���4UJ�qA���Wb�����a����h���8����$���6�u��i!��9�t>Pu0�m�<#��K�j��q�P��j}���lh�շ7o}�z�Y�(�[�n�w�ڬ�W�s�;gq
N��u�;�������J>������O��M��c:n���+�~|��I;�5r�[�{��qEswu���O��=�܄�����;ޡ��vu�ؽ��x���[���m�k����]�����GBf��:�^�|~��������q�ds�ֻ>�������׷7�q�׫ၯ�����{�{{���h�a|r�-��
͍�mn=q�UFh��|[`ύ8~(ZLc��i��z7mtԼ��Ƥq|��,��QH�rԜ �%�*mj�AH�T8��Q�&�n�YUG�/$���2��gz�����4a� ��3mө�Er�Ŕ�1VK���N�i�6VT
��s����gF�50C9��Rf��6\.�?�z�3>e���,���$~:�s�E�_�2Go�|L���T"\.N]q�YR�8FV�m�N��_c��UI��f���|�m/2��p�r�b��GF0%�a������	Y-ҹ���UjD�!��-�fD�C��$��&J�Ǵ}��_��@���G�\Ѧ��J�g'�)�%�F�̢4z(�S�|���I\h�~�	�N�s]@Q���J/�i֏��BH�p�'�C
h�3�c�m/�_��W����߸���_ӱ�>�D� �M�N,Bը���F�#�A� ���!N���� ��O���)���p��j����`����y�3.o���_���������k�=��=;nŮ�:��y�-<���f;�7�_|�ŗg痮Y>v{�_���ߟn��~���勣��{볷��޾��>:<zz�Z��k�͚���K��߭�c�K����8����p9Jm���a�kێ���)�M?�
���0�ͬ�)��}��e�f?`9(�#�,�9@�9����"=J%2R:������ė.��)ݴs��+Lp�6���M9"�?ht���`v�"H'^K
��"X?Rz�r�)��� ���Y
ré�񁦳%��P�fB?�_]���J$�b��0N���))��_���g����=�Ȣoʈk (]9�p|:�V������#c��ls�_�F����!p���,)�BiZ.2_W��*��l��Y=X���Ʀ�D]�ᠵ!��4k~���D!E�%ypj���W���7J4"�UHGQ�+}B�׳�˷|�7�%�"��;"|����{W+�&e�����T�C��駟~��F ���˙��jR9��j�����8��I�t��ϔ�
��8�D
��i��@�r�C|����S�,�F�'�k�gg�NN~k[l����}���73��O9�=�jq�]�㻷s�rr��/���^���t���ǿ��+�������ѿ����������_���������~���۹�9���/n�={���Avo�O���_���$w7���׍jǞ�ί~�������_�o��7���Q��z;�9��>{�㭣u9+�E�x�m�@K�E퉑�E�������}�U�/���i@D(+]"�v)4�]!��:ʵ����ǿ��)��}�� %}S
��J��'I��*�Α�����AJB��@�dR���QZ��@#�)�ެ�?k!w��Gtv�4�~���҉�f��J��k��͆M�B�T!�,Nc�(L�89��E+T��fW�C�h��F� ��Q��Έ�R(3��зdu�ĜQ>r���(�y�d����i"@�Y��ƩD��hZq�j���O���kD6e���L} �Pz�*F0�g��L|�~��JRp�e��5��1q:@�V�P[�>o��,E:'2qM���=�j���,Z�R����\bd���(�*�N�fh�ɢ!#`��h�iJ�Ut29�k�6�����	�2bVQzQ�^���̖��Qn��D��-Ĵ}FP.�D;d@>$�%�,���ԭ��ZB@��D��Y"K
<0�15�\ &�g!�i~jh,_��iUfæ@S�O��<
�~J���M�_]%�L�-�Z���G���Hm6�x�@S)4gnd�D�\�ɚ!N%�8~���B5/Ħ�Z�i��5�F�
�2"!d�@Sd�!fQ@P���$^�B��NKR�4q�Dj��a�EFcIAҩ:~�����Ґ�1R0V:���i')ӥ�� ddA�%H��4)#�O�Zs�5CG�i>�Qt"�� ��B-�ե�C�_����39�t�&�� K1M���
����������T�Q�zLi^����gb��H9�8�q:^@~�f�mi�c�4�햐�	͖��T�_�I�X:uX��ড়NK��,ڪ����X�q.
��b���B�t���,�U����t8�ӹo=/�Or2x
�DN�i�A��O�t��ЀX�����D��#�fL��zk��M��PP�A��J�r!����Y�S��� Lb8�ȵ�S�B[��9޶k�9)+>�C���-�R�9C��ƺ���d��!��t��Oq�`��k�js�#�ѧ9��He���ܭ֭h��Mr9os{�s{�?�;nT��S/�~xt�޸M��]W���q��eK�l��_��a�k�����ˋ����C�ڻ���m��խ/z�����;��<�<�����p�]��vX6w���s�i���ѱwʾ�B���� �V��n����X�͎�2�߃q#&_ ]�����g.[��g�\��p}��?9R�z�-����ɫ�;��n躬��tݱ�_C��񐱝�l1��[m�&ȱ�@!��A)
aBr;|J8.>��A����P�SY��%��DN=M��N���=�>v&���6ud�ײ�S��-7>��5��H�h#Y+�RZZ!Y�D��?>��?����τ�%rZ�ҭ���W�E�m��ɿt��E �8��2G�������W-��iE
\u!��M���"���&��l���5�h��[VT��Z��ThH,��Ȑ�����P��3�g�qN�� �t��v���d��p2�8R��!�h[L-�r�����)�\S>��s �D" [��	i�#�>���r�@��#k�Ȧl#��S��&�2��/j��A��J��^AJ�?����輳B.B���a��u���e����D'�2͘�V�I�[om�ۈ�2�*�^?t�)��eD �:dhM�5�'�>̔��Ǐ>�t+Z���}�{>����O/R��Kf5]���6m)Vs�|g�h}��K����L��-����_?½,zYu���s���d`�%�1������ݳ�G�^�=�<{�������mw�r��>Nv]��n�~��~>:�Ÿ z��|���?�������v�ӏw.�/������nvo��K���~���{�+y~��nǇe�~��v<`]V]nH0��x]�B�l������n�svW����v`4��[dl{�p)�^>�C8�91m?�q>[ZKG���?�E7������H�`Ls�9|�q엳G?�^�OÝ$�&�c���WN.�b�jFS
��T�j �Đ崆 p�r��>q�(2*~=׆�Y�Bp6q��'%��H��2j�|�oDP��BФ�r�W�B��2GV�5MAS���ϐ-�TQ�8FK@s��p�!�96V�����h��Z��@�q攠\ �p|���bN�hL!!�a5OMW���,"��L���:��-SQp��!��]K��p�\uuW�B� B~L�7Q4EsZf� -��#�,j���Lv.g��z$�8���O�U�x�z3er��&�aߧėk*dı@�x�n�4P];l0!|:�Tn_d��y^��Q4Q��`j9�d5fj�|��a�@Y��ȟ�t��7fp&�T��ij��fm �%C0k�� ���S����ã`�3�    IDATc�j..��Q�ӳK��G'Ǐ��N\[���x^^]���ı�>�Wg�w��;n#v�:�o<{�����{��e͋ˍ/������G�������Ź;�n���p{��]M��7vWǫ�盛���Փ'�(z������o������G����ޡK�{k�'����?�ƍ�g_Ҷ9mQ;f���C��-��Ɏ�=q�=s�f>�clW4u:�0�f�2:����U�ߋ��!��f|��NL��U(n�<�-�Ք�Y9>���o�pj�J�U-C(��i4E�e!�'_._���V�i
V��3��~k�j M���u�B
�[W8��C���,80��	���J!��
����T7����k/�M�s��*F"�8�U�U7Y�%�a�kL$�z�K1�N����:4muhK���?��z#X�Q��B%���	������)��H�ԢY�쇣sVTK�@�o��US'���'n*$�0"%�ԩn��"����J��� �ϙ�9m�Z�*�)�I�c�2$�6�MSŔ^?�)�8Lʶ'�/���_�� QԈ�Δ�K�\8&Dz�q��qrfnjR���~b"T��Z�\8rS�tT�A�!1ɚ�*�Ĳh���@�N���9�z#"��/Q����٘�x:Ɯh�Q��3s"�Ec"�F �R��p��K4�"��(�;Y��382�f���P�䧀� IA�tpf�l��������ln8Ax%J�D>fR��94E�n����ff�{�4GbF����� RJ�B4��01��p��2�bYkG��)�B�U_� ����`R"�� q�i�1Ŭ�D������,g�x8˕hT>��4Zgo�Ƙ���!��i� 5 C�7~��![�s	�|�[?���!�vNQ��TZr)3N BL4`��G���đ����-��J��gW4&�ږBFщ��%,�CQ8���pc�h�E�g���;+� �b�KDˑ�S��mLN�dc�Y.�rp,\⬕�)N�p�C����6j�*F`���7�߈\]S:��f���IU�=�(A�Ԙ)?BE�@d	��b�P�X��&���{���a#��iH:|!V��Õ��FMv�������F���cf�Ԧ+���F+�,���)$^��~2��K7��=�OT4��"�������rW?���l��ٛ���{��Y�7;�E�o�y3�w{�����n�7{�G�7���m��_���\�c�㷁�ݕO��9���p���w#�G���]��n6~s؛�C�o�}������u��+�?�z�>�JRӀ˭�J�.}���|��x8�l��N��w)a>��\�t�s�.̮v}_�VW:}՝�|�x��뫖}T�4�vw���������g���۫��˯����j���mRX�[���u��d?�s�#؁y�@:��|
5�|G����>���<>r:քfMA���q�D�p0�X�F�Y��)q�,m���P��4r�8�q jƩ.�|k-1�Gd&�M�g���G�v��dgcU
�:�H�����RbBZ8զ�h����Ə_.��p8���*�Ŷ��t"���?��)��/���)s ��!�듾fZ���$���g��(�ad�҅0�Uə�#f#Z�u�*|���z��RZH����s�����G��ݓN
�1M�Jc�?@�v&�h����`�v�C�U�1Ť d�K�ÙI�Su�D`���R֧U���R��@��<������FKR�C��@�ue�J!���L��!NE�ɢ�7b�9�FH�(>A��rf�<}�Pv#F�x+jj��,�2�7p���w��ݿ���z��!&�rar�C} �j��dZ�ե�	�^1Le8�|Ƈ�]8��L>s��S�.�ks�8a��^/���G{���'w�]��z��?����h�����2g��ˍ��mԯ/O]�|uq}���g�'{�^~s���>������/}��ѭ�s;�ls���w����ͳg{�u��p��9Z�]ߌ��7�/;�\W�=���[��ȋ��qq�yܑ�����,��Y��Ph��?�4EG���������#��m�:��D�[�3L��冴N��nvz�t�(��:�#�I�Rp^)��ӧ��_.�D4�5�܃�	p��S����q;��Cu�
Y���U�PQѶH.��V� G�5�D��ɬ�(�S�hr��B֥�ȓ�%>f���W��HɭQ��@2�\~��z������!^�i�Ԁ�E롽�O��j9!��6*'J_u��V��q��.���k ��|���84QOa#^9>P���cZQ�z���5�B�N8�3E�&��J�qMI1�[U�G�rrk&YSY86���vŤ�,�,�o�]|���\׬=:jCE-Q�P�;���eRp|7�w���\]�&E}�����w����QJ�gsg���ɺ��!p���s�������d �M9B~�͑85M�ۆ��Fj��D�D������Ӌ�B����ë˳����x�j���8y|���w7�_����W��b��__���q}}y�r��c��v$˲���<�GFF�PU̬��(R %���i���F�@�R_4�$���H�(%k�̪�Ȍ�gwsw���{�2%{�j����ַ���y��c�^y	�75�����wƗY���o�..O�7�==��鉏�xi�������{�f6wG�G�;z7�7㚨����s��>Jz�K��[�^�����ϕ�,�.�㼂����z����ޫ�/����U�r��jN�Ɇ�|+��u����N?L�tO�p&%��b��ͧƜ$�8>SԸD�!�c*d� �����Ĥ�b�i�X.>)>��_�
a�� 6@ɿ�_3_�����#y9���(��9}HS#��;�嚢�K�W�!.ںtn�VWє���B@=W�0Y�|c8f��R������BKWDf.�Tb��4�Y �PS"�9v �C��,�fu>q��H�qȎ�.��PY��ړ�Ǥ�E�$k���MBY�4Q�aR-�I9���Z"QL��[�#U�Ji��E�І�r�9�6k�S�ϩG��Ѵ��1+�l���q�ėR�}�h%�e����*���b��O�ӓ�(r�tʒ�c� ��N`QH+B�����M	��7F�K���ƦLsF�A�)+'�hS048�q����9�'��2�cQ���J:U��#]��=9���	��!@"�!�+�0��D��l��:(+\��8e�'�"� �ُ(�>�j*��F3��q�B���0G������\>��r������Ffg��D�A�m~�d���ϙ�������@6}��I���R����0���Gk���&�j�@�t��U�8r5��f� 1�c%��4M�LC�JTN]ǯ�T�XZU��J'��u�������Z�ZrM����� :k��#S@�	�3�pLӖ��)�_\|��~��i*���n~���цhf��t�/2���G���K�?�$~�)��H�f�TT4_� ����q��Ɨ�I
�錝�EnZ4ͤ�'A��0��
AD-�MMH�Ȧ�BJ`B��_�qn!&�)�G#տ� � ��(��4m�lUn
-��T��� �hR�H!����
�c�J�_��-'2�tF��G0�\���s�q$Z5�i#٤�Xuˤ����8FYF!c��% ����3Y@�ar��ߑ� f8���U~�*(+cՍm�����E� ������3`�����OA�_Ś2L%DAoH��}�҅�qc�m�W�o�<� ���-=�%Y�ue���b�M6o��n.���p��+��#>����}We{o��d=�-au}���>./�]1ݺ�<�ޫ+��w>��l��{Ae�pzp��������_��wn��[������ե�Ҏ_�rK���>L��S�~L��Y'²�ni���9z��u���~�HG>5x��H\E|S`���} �$w�x��Yye>�]w~g���}tso���`ɱX[Y�|#��yeQJkc ���o�����2o]�{��djD(�Kt��9e!̧J����')����������*�`�`T%)46����X�Wc6�cd3q]�+�T��כ1~����L���m�q�kdB������_����Zh�"NSGdv۶��`�Q����V��-8@��`���2���>j�*l�Qz�N	>��W�B��S�ҥ �0�/��B۷t��8���+�$=�_����H��
���i]Edᧃ� �9��A��X����MeIi[ 4�̪�'5�:r!Ȭ�j|��|�_��d)��Hm�pj9ᐪ�:oE�ȉ�G�7���*��1R�tJ7Ja߫�δ
!����s�Ьe�[֮˨՞ ���ǌjX�7u��F8Y���@��x�Z	�F�o�R��{�܍g��X:��|qs�i�q��]eL��&M��ՐD8P�uuQd�a�;�O�jUK���S8U��r�s:�4~qu������/>�����������)��CDN��~����ΐ���:����ͻ�7o7�������ꫯ�}����|����wޮ�5o��oǛ����=<=<ؾ�>�ş��GG{�.N���:\]]�=	�;�0��`u˿���zvܭeY��:6��!��:?�Zc�m�A�ۊ��
�I�}3�e��h�o�u�R0��,���ɨ���g��\d���r,�-�� KWK3���Y"�:Wb�[B��j@H��(J��n
ɚjL�N6�
�6���� �#�C��*jdu�)j�넂dH�v�� �h�q�pD�)�6���q���B���-�ZB�B�FU�5f�L�eƤj��Z;��+d���Q h��`|F��F�#�H��0��&�7�ί+��\Sc��M��I�	fZ")���(��ǁݐ��A��\�YW��1xg2�rF4��'-֔����ٹā��xJ��ų�miړ^]��6$D!��h�Ԭίd�L�դ�8�B����U�#A�,|E-��h7J����������/a#�6B�P�oBh��2���(Zo�#P"Ä�*)C�l�b�G	�Ĥ�BB�`��_��Wvc!�h8rї��xr����W������;ww������[��㞱�=/���?/��/Y��?\_^{}u���򫙿��g�;�����}��������W?�du}fq;>���������V��~�j�`g�-�����.����ͯ�~���UӋ˻���C��V~J�g�࣡����<��}�s܍�cw>������l�&�]�R�h7Z8����q♊:�N����I���P��@c�4�t�L����E9����WW��)re��(��c2S�R(�(��I����ZG�R��&�H�E��OpQ|��+H�)'�֔��3~g�f�C�"c��
� M.M"Zϟ|��(0YBn"rS��V�+�cL�c�)+���jX�M@�t%�f-�9�r�R$��ӟ�|
eͅ�O��C�4�_g6�TȦ�B����
a�w�fYU�0f�s-�uC`�9B��M�4ô��	Ah�5� ��̊SP��J!X���(s���l�*�DY�=Hm�lʈ�U��ݢ��E�l�8�R��Z��F��Ⲣ@�9��D�LsҩV��6���̙>N� �hr�s*jj���3A�Ǡh:3�&B�L4G#q�~��j@.��u�����S���~ �ಲEl,�D�JL���I$�Ɂ��hW�`,j=�\j��҇�D֏|�PQ�5l-|�%���C��=���y�+	YT�G+T��������J��˝�#@�꓃�
�*aj�w4;:BL�����r�A�(�h:Fֶ���gd��:~B�H�Y�%�M����$D.=�*!��R�.Dt�<�IGh:*��/�������p>A;�T�iE��v�_�A�{��4K��\��K���C��\�3��/ݘ�aBFY�)��`L3���h|4N}"EK��EU%�\f�*�H�BF�u��q��2�g=�T� ǁ���|t�2Qi��lD���׶В4��2��WRu�荊�!�L��V�)�BL#�hxR���)+)䬅(����O��%��@�� SJ
��q�_��B`���.ڏ�6d��J3�ƙ�B�'�B8'|:I���	�/�w�w�c����)�6]_Q"$v,8��L�(���I�EWT�Q-��7'҃�Q��Hp6�1��Ȭ*�"
�	�]��Z�htt���K��b%z#�1�m-��F�þ?��K����ޯ� �%�Ev�8-��e=8��Ǻ49Jخq��q�s|D��Mm�������������l���/[>x��i�������sO�-�μ��ڶ+��@�����7q~�"�M�}�Z�+���������;Ȼ��D��}����?������x'`��o�\�r��ؽ��l?�ٽ�����R�����k�]�6�
u�tk�[�[w��I6g<ϳ�EKv�3ض;(vA����SQ�ѹ���k:��Nd�|⤘�LA[�ghzbqV�S�$��F
�1�Z��G(=N:���,ڔC�n��&��8S��/Z!�h�+�!6�hm����"p F4N
U��aM5ДC��N�O���H�!@�[�)�7�졇�D����4�����o-��e	�dcE�3�e�h�Չ�} X�K�w�˕�s�9DQ��2���#�)ʈ��9Mg3!M�D�Ϛl	F䡻����L;'5�C�n�U��H�r��F��@�c:[�X]!�tcV�hn�KE�7ř�n�-
1�*� (�ҦL4r
S�t��\�nE)�Щ���p|�� ���1)
3%�̯���&���|u�8��%�N<;�p��GB�/�d�-��p�|�c�w��y�Y.�?��?x�ۛ��ML��H���(SC�k�9*U[>C�%G��c�h�t�<H( ���pX[�i�M���;+l����kdN�ۋ˳qKƋ�O?ع߽�>�?�_��zw���7�s<��Ym\�m����k���������w��g�[{��on�/�ߝ����ݥ�2>��ᰱ�:�9;s������غ���������l����j�������[�V◢=��l��8�mO���&�t��l]���,��:�R,��
�����3��%��>AǏ~Y��8"��M���w8�>݀�*ZcEkOT�tS}:�|g"VQN���/�x�hچ���T�"*�n���G0�Ap6�_9��芏C��ɑ�G��L�ހ�e�4�1��R"h#����Wѣ�AԔ�Ԍ@�c�4N+�J��2N�E��q$Z�����]�P���6J�+S�Ʒ��͙jp>k�-X	:���Q��UK� q�EU�Թ���!�jAt��#�2�3���6�BU��HI�:5,�8�Q��D��\#x�I��*��U�w��0�&��PK����9��>:�zv���ZY�Cz�� ���HMȓu�"�WE{hFf�:d�u�}�Sԗ�_|��'>�b�L
=luK���M������7_~���45/�7��E�g�_�fL�AL�*���!R8��c�P�"�	,1)cY��� %����X��i� k��C`c=D�����>=v^�?���룃흓�W���[���S>5�C�j���=���8߿�q�rO~�f\�t�s���w�'g���l��tw���'?x���ջo/�N����6_}��7�up���'�_�9=;��t���r}u}>N�]wӹ����>�s}�	нw|��_���#7�����ҧ{�^޺덗O~��Hlo��o+ƾl� ���v�2�ybg�x�mN;�Ia��1���	�Db�SQ�#J_.���)�ߑ2b��HL�lĤS$Z�)**��)�"���궬F8Y��4�T�DQ�@Y|x)|:����Gk�+�[���&R�����L�*-3��E�qCD�B��荔,�%+��7�qt�A�|S����-(˸n!R:�8�(�Vn�'�HA����P����b�3%�N��a�|c��9��P�"���k�`2�S�TKR8�&'��u�a�F!��y,�!D*:S�F��h���ɯ�@#ku������k�=1�h2�YNV:�hD:���ު��B3�Nщp�H�9�Ng�Msf?bpRS2S�RL�pX|oc��    IDATc�ϙ�?E�Nol�F!c�Z�X�*=�E��D�c�ޣ�~ �M���aH�P`@S +�h3�
�Ey��c�N�t�R��+�(�
MG(5����1#~��X�@j59���Y���Kȩ��f+�OYTzk��_$��Y,�%;�K��BLx̢�&�f��1Յ�>��ZI��Nu)8��9ą��h酪m��G���,�X-�j%l&��\Q�D��C�ub�����@p�CdfAҜ4�
�-d��I��U�LN�g��̢fC�2v2pp����c\�����z�䳖#b�2��c\��&Z�����u� �x�F]U+`jF�Ƣ���t�a1�;�e%H�>��;�D��FVoDX���)
�\��������4��V���t�1����y�~|�Qu��0q8_�98�iF.��o��I�6�0�U�J�(�V�m̯�9��āP62rR�Id6#ʪ�	Q��dq�@����嘆�fh!���Mĸ.�ߴ1�D�ǵ'bLVєK���Rh���`�@�J{%�P4A�cj�Y�(�� ְ)�B�E��6���^z�I�ǻ#����`��2e�D����R�e4{ih$�U�L��{��>O-_��Ay��~�W#�=�ǽa������I�
;�^�z�tۏZ��w�ż�-ٵt�"K_�~�e{��ү���1%�Gu�x�|�������G��ؼsK�#W����wt��b�S�W��o޺���Sj�Mi�Ͷ��Dc���[?&���޽w¯���"��.�f��9^��z�Żf]�t�s�铃Ó���ƺu�бksۯv�Z�;{L�m�_�_l?��?:��y|���coe�^��-_G�?��=*U�ұ�%Ʒ�AZ_*B���vP�S`���v�m�;�%b� T�^j��=�Q ��!�r ��FSYD�u�/���
�-����p�R'���,���t0!���P��1��3�K����zW$�EI,�X�<>���T:��1I���*ñ?�YT8�Du!��@�Z����?bV�h�ڷ�5���l�SW�j��fz�Ҥ�aJ��cj4���
H��z5�)���̔�kl�� �͍�U") ����D�_���"tD�����}�8RPўGhi@�eE�@����Q���t�8��e��(�l�pS�1S+0&���&���^W⺸�,��C���Z/\�h9�q8-���*�&����)�D�O\b�*��R����7'����[)C�3A�*z���D���"���.e�����-G%B����z2u SYH�t�y�3�Ư9��5-�ڌ5D65u��9�~�Y�g}6��/o\���������~{y~����������;�ۿ�8�ܸ<;�>�>8������?���os����vh�n{��������M�.������2��6�	g��׷;�����'?���_��?�;��꫗�oo?��6��0�Z�I��΁���^��1���>�~V���3;��y�յ���cn��l�E�Cl&ޱ��m�m��|�Ҙ#���"��B�	��G�4p����'8��AG���|!�5e-�~*7��	�� EVoӢ��C�����FL�B|p �3����A�%�0P]~gi����2���#�GC�R��џd�M�(Ŵ�4��:�����Xɲ��T�ˑ���=��VW
�j�$�b!�]��<�**'}NC$B�b�q,�a��4�pJ�wAE]��T�L��Bub!�F����1�D�:�K$b�D�Ek�O9Ĺ�V'@V-�sZ����s�r�<�M��F
Bb��.>p\*[6Szu�ޢ�iьDtb�g�����c��4Au"�����L[�����3�-p烺s���D�K�.g*ᚨ'm_�$EV9��p�ʪS�8L{E�:G��9�(���02�FQ �tV�tp
3!
�3J�j6M	>\������������o�����6j����Wo�������r�~c��h{�U��s���q>�x��|�:��l��w�߽x�y������۫��g����������������g����x~��W/���/��,?���'=��ٓc?1�utp����������xuㆵ>ʺ�uv�򁃍�z͋9l�
p܎��� �������7ܫ���S֊����V�h���C�����,V
[���X�W�8����|)p:@���6��?ߘ~F�-&���U��$ը%Yh�+�*���J7M?�H�H�ُ��V�҄*��xlL��3U�2�gE�3EV���l�L��9���?%��#�1�X���Ȝ�#��n�'��R+K-NO�||��p�H�(+�Vq�!"U�T	�b�zc�9L�u�g�l*ā����&�Y��Ei�ʪhm}!s���T���P�H,���<m���i�1�Z�>�
5�#D�9SL�B�@kO
��~�H���*�r�bJ�p򍓀SE��M)�h$��'���!4��3¢Q�8�&h4ř�/��&����WN-!#C�7�6Ҍi�����)�)�	��i�M9��Ԛ� Z��������ȭ"j�;�G0�����X�V��)��98@S�`�#��q�?[�1���MYOוSf�LU���)���r�)̊r��T�1��S<�Vt�%��	&"�O>���������`��ԙ����C�<w��r��7�ϗވ�	�}�����G
��R���UJQ���iF�6�
�ş+�"W�&�pv�qd�8p��dv��LS�jZ
�:�)ۇp#�P��"Ӫt�9+ ��8��V]m�Z�@`p&����/]
_�ic=���L����ki�Mk�X	 >VE��<:����S@ּ\䩉S�Q��1�ȊN��u8��j�� 2Ks(��̆Mܮ����S3��V!�Q3�"��:���8�M#�W��2�N�.�j
-����m�a�E���FK�&;9r%F3�`�/�#�t#e�����4
A�lp��g�֧-H�8�qL���9`,<�D4|��������J���B�^	"��W瓪�Q�W�^�גs���,&AZ�N�Ȍ3k�� f����t&����h��Z�Bhr���:�&X2�i8������?P�ny�d�d�#�n<x��ô�{��өz���;	��Z9.���9n0k�7}�����Y��!�Z7��m��#�UY��Ƹ���r��Q�eX��������?9�>��30w�+�wu�;�M�!�3�g�O�9.~���d_#?<���?^΄�yc�4�˔�˝�ƅJw�}��vm�ȍ��o]�ݺqK��~S��ǚw�}���}�u�s�����q�^N���w;~������~%��a�Ǜ�Ҧ%�>�U��Y�r��bۙ��p�;�[̀s\�ms@��h�bB:|!�􅊦��A挣�w��,�P�4��Y�䉔h����0J.��Ԭ�YB�?��aZ��J�d�AL�T�B��mQ����%�q�C���ad�Mq��O)r�댠yYF8K�6$B�P-�l*��Ls�{L�{N:�9J�k$�DSƬ����M
q�rL�b�TQ����%�V�2���~r:o��)^o�f��98E�
�
դ1��"h����!r��_"�2KM(G��i#�������	�$�N�t��X8~E!�)\�ҋ��:!��z��DpX���1ө�'��!��aJ�'�Q9��iN�)��9&��l�g�ڄZ�#�z=.�"8I�����t�sz����Uζ M����5eEMk>�~��BS��jP��ob��G?���O�|���ls�����~�������/������������l: D��S�a��z��ZO���s���h@�̀�_�\��r�?����;���Wn<��G������{���7{;'O��'[g�|�f�,au}���]��w���7~����-��=;:x��w�O��Ѿ?]{Ϟ�<�Їy��]]��w�ܘ�=��`��֑�Ư�O���������=��^�^���Trü���09�W=19��o9g��a�ё�C��YK]����#�8$C�|%X�(['�Y����å��Pu�n��<�%V����_�@|߫��qVA���;�j&YRp���cY��BU!B�Uw� ׭!)FF!�ϑn�ƹ��RaNK�j�iK��m����Զzd�$���d;:R(�kF��J�a5YV�BB6���Y9�h����?N8��¡�g�vC�@�礐JD
GVSL|`{���(N�|4>�V�.E��Nΐ+I��Z8��39B��α����"����h�BN0V��a>A�P'j9F}rT)�6�������@
�(��u�!�B:Z��]�e���6\ ���L��V˚ǽ8ĩ�8ժ�J mK˔b*jK9i6����ݓ{���	�hK9>�����Ϯh~���h�|��Ô�p�,f��o��#��q
�K4���VJ�JD��i�DL9��'lZH���=�l�W4}{�3����˫K���_�哓��7��^�<?;��Ʒ0�^�H/ܜ�G�[W��O����?}�����Զ�l��rGϞ|��������������ɍt.OO�������[���{}t�q}��~��=�8to[8�>{��Ǯfo���=�|}�z���/���W߮����W^��o���2NB�6�w|�ҝn��E·��/>��/�:w��Wg��Y��������1M�����c�/�Nzp��	��Iǔ���9ɀd����i�N�z��"%2�8@F�5�¤ Qf�-���h~ ���J�I�g&B>�:������2|,�������
7��O-�����jr�6B�5�p�9��6'?rӹ�t�jDH6N�zc��T�S�|!S��m	���a=ɀ�r1�!�mEE��q�|)�C%J�DGn� a�l��_9�H
R�t���8�3��5Ú�h�����3�1!���82P(���5��DY��Dc���&2�R��!pl�zn�g
hՒ(��E &5��(��ϖ��Tx�1��1J�a|��τ�R8�өtc!>�l����r�U �z�4�[W�b��@g>Ƨ_K�)[276�~|:�+�WK���Q(�A�W��3j)�(� �8�"�>��¤7ŉ��+!�ǉ�G�7�cR.�(�W,?���O[Z�+�Ye�h:h�p
Ŗ�f�1���������D�Ngւ��@ugn�	M���Nbv�E@�v�d���oL�1r~Ǵ&R-dV!����Nd!|.$d�Т��=)Z���R��)�B��O�&*��j�he����`�A���L����L
�eʑ2��%�B�#si��p�	�E�cT�����'RS`Q>2Ӕ'9�4�����w�d!`�Y�i�l	��LDH�l����j��Ҟ��2N.�P�qZf�s�J�G��3C�!����D�|��r&�?��VT4���-�4Bʲ���!�߳���DU�\���ζ��I+׈S4�8�t�x<���7U"��i��aM�uU9��B��<Ӣ �h��_M�0�(�)7�3����F/�ǇP�C#$W��ut/*�Q�E[~̞˝���xC�;d�*K��d͛J�㳜��D����C��\ޕu��wN���)�T@�
�
�d˥A�&���R諈~�ҋ��Moúh�e�î�t!w_���~���xoT��:w�v���ٺ��U"���Yǯr��M��]ߝ�Rws�o�Z����ޓ�}%�����mVttv�4�v���W�e����^��l{�i���&:U\1��_-����^�.�������'�O?8v�[o͟�]��y�xow���?6V[{�ۛ�L>v��]�R��t�ٻ���/�
�WA���xc��{�+��8(v{��q�Țr:"�F8P��Ę��J��'kt�&��>��I�Y�d��;�  �f��p�0�7�1Z�Q�Ѥ�N)��?����������a�τB�ɦR��4U���BX���b�����������4�(�p`���dr��a��8FE���B�9SG�������r�ug�G�e��Ԫ)�ͯUǔ�zo
E� ��|c��2�j���ű.cӊ�2�ɗ�^�/��YT��K*Jd@����Br!RXR�E��>��@#&��Ғi�l;r%����|HǋOJ4G	)=��M�SK89RD��r�F�d)8R�=��������(���$�V�\� ������F�!��
�JH���x���.� ����9���R���/��'�Z@+�׆������W_yO�mi�����}��{�;�����o��p%Y&���� j{?�H�I��|BՆ��tm1 ��Rj� �-��n��k�7���}����Ϗ?��3�����w7�!xq�����?�涏���������o��{�o�;8bne{s}��}�������۫�Oݟ�ۗg����ݿ�޺����˫��������m�H}{s�p~v���z5��s}s�V��P�gr���	�Z|���8Y�%��ҧ,�so���<n�@�%�M'0�:����q���?D!L
��Ɯ��rrG��RDG���%r�mt��!)�c�wYΰ�>����7��ñsT�w"V�BS!~m��	��ߋ�/.�o:�4�o��3�|#5Ɵ�i	�������M9�a��8�88��D��p���@�Q"N땮
BjF8�S"f )4
�b��h�+!]���t4!��s�PT!�F�i)��9eQ��1�lgR@k	Bu� ��\Ȭ�����������F��oi�v�f����\���5�t�$�xmN���hB�t JC�:�+8G��:� �
�p�B�)AV3�p��DLE���I;�VV�V!E.Mɀk���ǎ>���5�˓�.��!PC����
�ZU� )Yp%��h,�ZU̇#D�Y	9��D!:YO��8e!p�є[�ǳb�%n���o9����gO?x��.z��ŋ����^�������;���y�qO��p������7��6<A�;VwǛ[�w�o��?��Ov������?�_��ܸzr���������o��������ķ����_���3/���G;w���~���f|N�K����߾��ؿ��ؿ��p��}i�w/Oo_���}�f�p��}�G�6��_�u�|��f��mr�v�­��b��F����Tw�8�mc8�����IE�=�3�<�!D(k�Ccv�!�"t��'�(�~]����C���Dg�ʙ��U�]RN��tV:���s�����#Nug�)Y]�6ʨ
�Ry�h"U1"�M?H�#�C!�B���&W�(����p��-<MLS�tdaփ��9�U���̴l�Ф��s��7iZ(�j��H٨�P�I�f]�ƥ����i��!m,Pn�r�T7�Y��'P?�S_��,��X�t�F>��jE3���YE
_:N
s�>k�L��g25@���� �h��6�!�Z
F�D��ar��)h�3�SCGK?)�<c�k)qS)�M��ɤ a�*-� �=����)���g�����,)���(�N��BG�(�q�T�h����#�Y��g��2:�M�A#?ZL��ƎȒ7��iD������%8f��Ɵj�YȗŁSH��,qN���dM�����ܶ�*CnI7���2W��e�R��K��%�M�(���*Z)�!�8���V-� c�qڙ*�?��B�7Ƈ�٬�PKS͔�U)��-
"�lg��[��I�B-�(X���$sDU�g!�����t�?���b��h:�\j�g-Y�4EkF�1�Z���b֞���!@X�U'| �D�R'��őӘӣ�i��DR��,�OBѤ�/��|�J����)����4�p�]*�/�4M�|�i��מ���D
�#���(\��e�4Ef�s��=B���Qi�H!���BD��P3��t�!B��y�M#���Ɇ@XYj)�@�y,-�����"Ƿ\8����6����)�<���<�rE'!�VM�H�p��B�f�jq�^��aҳ:�QFj}������7o�Ha���DQ�DJ�o]ƚ4
s�^����FR��2��X���O���    IDATi����b���g�ZM���3�ȇ[�T�x3�w� P���ʲ����[�q�|�}
����إD7�����I�qUs|�Ļ��1�:��i�v勊+_���\~`�[�w�:�����ݓ�Ã��oF\�P�X����5G�6�/k��_��������q�\3}w~��K�7+SwnW^�lz���(���_~N�m�������1o�����eSGg��Elz�z�_�V���/�8�7��7�n����� ��8?�����Ʀ�܎�������������Խ �75罡���U�&xXY���ζ-i�Yf�<���9c�M��;�p�B���N�(2��S�_.Dt��9	�x4�/�c�b�����JQ��*��8IIjiF�d8�J���&�s�=^&�Ǿ)��<��U)�ʣ`*�c"������T��?�制�%�K)Tu�+�oѤ��|8�13>�@!�)�N�xO���d�n�/F감tu!����G��6ԭ#r��6�(�v8A"ґьu[�)�I _�i�bJ�3u���_�,̤���6
9f!`�c&2�� Yֆ(Z�O� �@Rc�����4N���ZhY8Y
��Z
�&�3��iF.��䴐�p���J$�'?g*P�it���1)G��A8B���;v��x�1�i
oo�pw��E̾$�`_�s�ӊX�_�|��9�_���@��nϗ_~Y�q����ӋV�&<;�SG�My��me�jݔ!���m�� �h�Cs��O��:����ssp��1�W��1{z�����'npy�ss�����˸��?����O�n�%�&�����.�~gm��\ Y�b؍?>�����>�������'[�7�W�7��gW��~�������U��s��9�y���{�;?�鯩���m�pD�N�X�������qǄa���)��,��m���B�-��E6�E�ӈ&D����fǾ�(v�*B�p��z�r9d%�4���,_{��?�S�/���I�OA��F&��HG6�Ʉ�qj�)�r�p8F��S���B����!4�<F!RB�(���B�E�1;����+4��$���0���hV��ӪT(����.i��l�ZJ��J M��d���j�Z��|>�@�G�,&��05�Vj5�;��4r�B^F�ir�B)X���9NYK|���Q�G�	��@S q+��� Kq�N)FR��9�d�(�U">�)G0�=�h�aՕ�1EA���h�����3�]��b�B�)ي::���h�u��D �f��T9��}����<���U�t�}"�mHEé)�e���)�9�1���S)5�T)�j�S&�4����鲄f�(�Pc��Q<��,2��=#�n�ݰ��_��o~���4�Q�jf�aw�K.7�ټu�pOmw��7W7���t�X=�=9��z���뻗^�|�E���_�<?������w7כ���<�o���܍���zr������խ�`�]?#�	���|��ݷ�����������w����/���|Y��zӯ}zAf^���1>�:�j�KM��q��T;Ʊ��{����S��R�i��̅OD.r�2f:Cxy\#x&�Ek�Gյ�`j�E#cB��`��$Z��)4T��@�h�ɧF
^d29���\&��'�V��V�a��U�?�*T4�dR!
s	E[B4њ��¥@�g���(���:
R�5B��N+���C�� �Nκ�F�jҴZ@�1e!S#AՋ�a1Kl&[�|4e����1*D|!>@4���B1'���ȍ���i�Ɣ��'��ܪ��(qcx;&j�f�����<�㤬N~Ek����5�d�29`#P"�d�E�@��À�A�M�*8!�Ԗ������������f4-w:M5c9R䖨��1=�����g�C8���HA�����45�98�6��NN4~�	��3Mz�t���K擪U�CZHE!S_:5��*q����M�F~���8�>'\W|H=P�O�
MAb�pf�r����K/y��`*��S?u��L� �girb6��>����(ԛ����A`S�oB�f߫��įsj�d'h*шP�60X��,��R�+�ҟ#r��lSՁ,D��S����L�Y%rQ|̖én�\ʍ��sEuKG�P�!��/4ێ�(�SQ�"$0)�T�Lm ;���������Ӣ�����D妾ܥ���'^4��)���pʜY����*Ԫ���k���C�Onj4��!��o��j�׏,
p��q
J)
�����@
%>��	V"=�6�lE!K;��_v�"��	�!��(���e�9�4u�e%eZK�̴n�N��M�S�ꑁ8�D?J��Á��bB)WA2�`��҄���&���)c}�rMK��(_��i��;(ΐ�S
N�F��h�z��_�����a��PE~]Y)GT
KmNs�d�l���M���KGkB(C8���8�i]E�������ǑBd�jq0�%8�*!SbYq���z���D�
�YE��)L�B�R�R�=lgJ�O��4���V�����^3~�1��ug��@�-��]~7	�G�Ӈ��	��`u]Et/�;�v����o}��1�lφ�7B]�tEӭ_ww�׍a]ش@�qno\����^�����%�[��<}{�7C}u����E1��W\�����%M�3��w�k�WD���oNH�Ie�;w�{������n�����������/�}���/���k���z$� w	�;8���:y�k2ޚ��z�=�*s���joܪis\�U�wg��Ds�4Tt�:��`�G'�9����K|0;ܝ$NKR�r:��*��0�b&�,�pج�_?	Ñ�H�k�!�)�iE�ZBS��au���:�e� 8@ǿ���	���ሒ�a������=�����h�Ξ�'�+ݚ�Ԓ,�7�T��b����[B�|N�3���I�BE�l
VR-S�,�5Q��� mfq�Kl�陹�q�Njf._>����3)�(+Z?���8���(e,c��5	����|���8�z��oxr�C��	�yu)$��sk�#�e���1�"p"��`�҉�u�p emB���
F�F��~�dSP!>Z���Y�&Y>�t���Yms��eM)S�O��C�S<��@N�sdQH?�zS�H1�;��ҍ�:��(�S��u�t9�?�w�����R���]�٪�X��*D�ΌzB�Q���S'�D8rE'��4-���^H�R��\i�yu����E��'���Ӌ����S!zz�s��O?�������]c���Y��q��`�ss�:���U�������������ڽ�����8w��gO��|��[�?��ݻ��)��j�;���w���ՠ�.�^w�u��=ݑ��
Ʊ�9#���/퀭��fl'�c�)H�鑀��\rSco�8p�)�t[#���c�)$�O�9cf��/���$�EP��)��:vhk��9c�H�JCj"]'�L�"���Ҫ�qX;�_	E�>�)�j�i�V�?0F��lt���?�	�y�JgB���U[>P-�9cR5�/}���F'kɎ�%�P�uX�!{.]3�8�!) �c�êU�h�٨�T7:�,4���␊��,_�2_c�Dum�|�yO�)%GK�r$2j���v����V�r�z��C���`*���Ԫ���)����I9���P�����M)�ա��t�c'�,�a�Y��tu�����8N�zޫ�'7m����yۧ�B�ש�Dͨ�ƈ�	��@	�.�r�3�uq��\�Zh-�}@ �bMG9#�n�`��XW�p���ZxR"�p������͜U44�2}�_|���w?���%�{��_����[�n��J����G6����7._������<�x�����d��NN>��̃����������U���^�<�x�v��F6O��mߞmܟ]�>l����>�.���w�g��N��y�ݻ��������}�ɟ��_��׿;���[O��5�Q�{�&<^�9��}����y�v >�ji����6����w���U�|Q;���l�(�K�4k�1Kw��@L鎔��4%B���XH4�QԔ�چ����&&��˝>'�M�ʥl$�΄0}Y�E��O���,~-�����u���h�hɆ�4N�B-�k����k�S�\U1���'��p��ȑ5qL)�V��6�(����TYF)��Y� �H����b��3��R.W��7� ���8��5D����Y�)"TKBd-�ȇ�2A�~��ǐ>��Q?��S25�����(ԃ��#�&�Z�|oi�*�BJ���X����85'�V=hi��8F�0=��Y�=D�W���9fJ�c�����g� F~�L�ş����D�?^�A�A·��8��_R`4S!:�LDz|P�MiB2��f��yt���;@�r9���!ª��~Ӣ|%���0U�(�۫��W=&�`B����gz����!�+u[`��p$fu�7��SK�A-a����Es	��R��
���%%�,璿�G�sN֩2+���La�
�6�	ʅsZ{!�P�k�X���T�L��Id��S��vQ@�ߴ�8:d�H)Q�\�#?��B���R�y�S
�V!E���v�&��
���B�_��u!�Tc��"4���rS��ɄD�
�8�*1�S���]�Hkq�fVx#><_�8��?��BqJ4�DS�n�N$�:����#PJգ��B�i�ь�Vڱ�3M��3�KiĄd5��zQ4'����)�X{r����M������ā�D��8�t8�+���[oH�j�Sbc�1�PgeN%&�SE���\!j���I�����!���b�L�Hd���p�mˬ��j�:�g��ﻍ�O
b�'�a��N��*r#1�uz(M\�DncMS�n����9�H)�N��z���o�pH=P�W����5���Yu#��T�E�68,�?F���>��z��FY���b�:o����:�㖰�7�ө����C�>�����v�����Cpu5n����;�o	om^���+|�G{^S��uxT}7l�R�4�m����‎G٭w���}��a��_nC�9�Gn��H+�"<~N�7=�i�ޥ���M��e��=>P�z�{2.O�N�x&/��t�ƫh������a>�������x���=v7ww�wV��j����过�������zk�~m�Y����;���^��F�x����z��HՒ�u����;�R�q���~�y腜r�����[)Uҏ9�p����Ru;�,ǹ!$Q�B��4�`�U��8��D���`)JMG�s�1
K�(�Y:Ƥ�7�Z�i�r�5�a��"�8f�8|F'f#D�Hf
��RF�������NY	V���U'�1��gr)����Q�>DƁI�rN�i�Ҕ�CDh)2�iQAH�'p��}cSc
�R��FH]�25�?�J�t4��ȭ�\��!�B@�g�0�a|� �q���$0�, �s�hZ9)$a)Oe��(Q��BЭ� k[�T)����Y'�[22Hu���(�
�iR�4E9B�Tz%�l�B�(1e�~QN{�Q�mZ�T���44�Lh�q��!η?-���noJ��fj�Ôbj�>G���_-7#�h��oh{��E튨��	3��Х�7�I{#~�Z��5��ㄷM�,*ٔ�h�h|Jp���1C| ����/wn�߼u���oe���k�G�/6w.�._����.N�nn����[t���y�|r�}}y��}�g�~O��O?���C���6?|q��ã�{�4�J���n���������ի�_���m�>_�����?���?�>���E��o�v��G����|��ݯn��i�Ɗ�Erf��A���>.�}|��BƐ|S&�i�|������ɎZӤ��/���n������od���
���%�N�.�;�sRh�3�Y��T]��t0;�=}q�I��I:����Ʋ��e�G3m[;�1k�)w�
��k�\j�z r$ֆ�\K ��"��i��,#&k�+Q"0��!BLE>�=$ȯ4�E�`r�&����ÉH1E�'��*!�G���9��BK0e��I�uX�����3��d�&X{���8�U7m	rɪ˱��o�b��O�������á��d�UgD�:3��[)N�cE��I̢)ǁ��*"��y!%�B�X2��p[�� ������d�7|�������B֮�G(���4n��t� x ����_��ǯG.��t���?��?����f��U�d�g�p�~�*�S�h�.����V��4'����D���R8!B��8���.[�G�{�:�-z�҇Z6�>��M���]O>x�����������w�޽~ssy�C/vb�η���./�^�ΏWw�;�w�?�9����߮n�WO��>98���z6.~��ӳ����������õog޼�vS��������'���;�>/��o^�����\]�no�o<���pw�7��>?:^fl\���|�tl��ځi-n+쏭p��ԑ�c�V8\�t�8Ħ�����O�t#Ĥ�\���"d0'.�F�T�l�S�N	x��:�OA:��"�M�!9���b��g6�.��Y.�iM�1�i9%R�O�S�j���ܢME�z��K9��!'��"qh�
q��D��r2��M� ��iRQ>�h���L��e6�J������'e)�@uYά��J���A��ɍ)�1eC��Y�y�����,�Ǣ�4�k�+��Lʦ�]�	�C�h�*�q;���4Ҕ���#Hl�H���� O�*�����:�C��t^%���q�����Q��['Д3ARs]|�FR��	j/�%YR�4��Y4�C͞�C���I
.�ř�K��C���dP�D5"0��hYi�����?�QM����IL>~�9�{��Tu���B�~
K|B����g45ҙQ��-d$W�����>��n��!�c�/e�B��*�MK�/%��i-Doe��1֭,�L��¿W�)���oj��+5EPe*�ӏ6;,=���S�4M�*F|�,׆D��Y�\mh���(��Ʃ�3�cl�Ȣ�U/�859� ��yȗ>m�I�L�\�ْdǑ��X�c����d�EvOM[ȑ��'��,���'������)���fm$A  H$r��="�g�i��0�}��jv���/�]:p����i@��|@��#T�����ƒ�c���iZ��_��v	5/=<��5PY�H��5������&<Z��TnwL���2�n�Й%4 s6ę4�h����*�$�CR���J�G>i��R�_EV{���f��L�1�V�yv�t�R?S3�RȦ\?8�*�(�Cs7�YH�3T�K�n!r�q~z6�h�!U�Uj �gmUI��["~U8Lb��W�,��6�D�!1K���D��JI��^u��"�6pv��^�Y�A��-K9#>߳T>�1g�qLgW�0�d��: �u�Mk��M_�h�S���hz�m"%���ÕrvD����8��fQ�>ue��)�)ޒ4^�hiLT:fm�950��B�������l��0ǀ�Sg��a�</}���i���+��9�vv�so��D�w��Zo��r���>�hY��Fу[�e�~|��׽\2.������n��JwU�(t�,�B.��y=��V����H��btl���/^Z�Z^�O{�x����v��损�A�U����~�����x��/�]ߺ�c��Q�՘~�lo�Z_�;��hk/��ű��v�x~n/���N�"��8jm>�Ai�acE��9�(�gl�r�(�P�R@�{6t�{�cџg��5~��S���҅�H!���Q`9c-
2��	�Ct�:��.C�Y"�&�\'!���dՉ���EA��F�r9,���+]VY%����q$&�HM���0���Bh���Es0.Y9�i=p��s�2ŔR��h;F�Tn�M#H$ʒR��F�r�&�5�f���4\��Ȼ|�JC�K/��&;|V������(0EhRf�&&3*�(tO8����'��5`+��HJ:�(d�bD�0��,Z(�o�    IDAT��Kc�4��%���+���l̔�v�
��ȅ��N?���I��%�q"H� Y��zk�k�_nYs��M�ZYpH:��lʡ��'�K&�����+�^9��îDƗK�/j{��I�;�ޙ������~���_y�ۋ��ӱd�2�ׂ�"�:i!�2d#�Q����B��Hԅ�ӡ��ZӢ�n���r�uc�����vs1�q�l.|N�ći�~�?y��ۛ���o���\o�o���y������/^�q���G{/�~���W��_~q}�Y�l���N��]yp]o�>��㋃�ˣ�답GÓ��~���X��o��܃ڸ��	�p�+iF�㐌�@4V�1y,z|x��|FiY�8��
��es����� �h�����<d���i*�,xd��"�ց� =�;!�:���k�}Mg����_r�]&❒���H}*�v�Qs�!8����u^v2���� �����Ј�V+jo+�>��di���DF���m��o�rd��8|d�ʡi,���1-�B�E�b8��ͅ��,��)5��`$h7එUT�&�c�iV���ݱ?-s��#B�q�R���ѣ��gE�)\��^}"L~�$�Ub�V$���cF��2M�3�Vm��Lh@���v��ԩ4��pfck �����(P����Ù���f�~N����唞%�I��⻭����4D�;���0�JCGQ[MHʽ�% }�/<>G�8>��r�N`���z�C4od��:��2���B8�b�Nr�z��ʙ>eQ��!�ƀF�LV�=�.j����V��~�������f�ځ��+�M���{�����x����o�qդZ>s�S*׫��O��ח��v�����{w|����ggw����������W?}��;'����m��'���ߝ<\_�^_l�������W���|l�|��ދ�_~�O��tݿ��W��X�崲5��F=+sŨ���������&�|g�@	�k9���h�,��7|���h*��/��Iu*�,�#��6��8��с;E����eU].�����Lu�8d�������e�R��A���p��Y7)K��.��+��U$����D����g��($BaV�H�I>����|�\4�� ��ٺ�ᖣO[� �� g#�7���
F�Ŋ��Zƽ�\cM
��Q6����4M	��5������DR�p2!N
��+q"��^�^e���6�G"�}�K��3!N'|�P������5�xm�r���7堅���V4�V�rbڒ�g3��&EMC�� ��V�ᘖYK3*�[E�)��`M���&5���"��.�z6��\�@�R��Ĭ�XT��uB�LK���-w����b�N�%�S�a���Qnd�%�6>Ĕ�1�F�3eE9�Z�'��&2u�*JQݍ���i�L���ѯ(�B4
BM�}�2�<	d�t�8|mT�}K{Ub�Ԧ?���TqW����LB��,���E��A��j]p�Bp ��NVn)�h�6��(5��RkD����X�t�lN�4�?o-F`S�ɇ�B;��p ����0k{IKSѺj���ѹ�R��X� 
eU�����R
�+gZK�ۦDp?N���v8GI5���T(kx}_�#�,�f�։�*�,2j@B�=[��Y�Ln�����R"ͦ�vA
��n��dR����f�Ñ!�z�Є��`�G�J�]�D��iB�tM'?e
�7[�,�����/]J'm�Ai>�O�&wC�b��%"����0�1j�,�8J�`�pZ�D>���Dvϖ�(�UzR�2�"���EF0����4�I>A�14
B�-��"�
H�Ԍ�49-��S3B�a��	�N�~���1k&N�!$PJ��*փ�r�s��4��7em~mW�߃&��p�ժ[R�M��L�r� �{:i�/W{g��M���"��A�ҍp/��#Dǫg4�"l�A�`�q�
��S�Qq�$s�^�t����nC����[G�C�zQ�������f�B��k?��)�7O������ܗ
�]��7{>|rd�C�10�<����qr�w�ϋ�k�'���������7����z���iTqmn7>p<�����Ѷs�]�9��v|��xsT]Ϣ��U��`5�P��j	/�ϼ�}�ۃ#O�]A�P��U�޹��T�$�:9;߼��:�˜�+�v����vj�����ێ��s�nw��������$1�[4�)]j�󳿯���b���N/)$���8�|!)��� ���Z�F������k#|��W����r���дfHb�0A�S	 �G��8�u�^E�"�̅5%�����|�n�x�LȒ*���t�r(����*�B�7S:�f'r!8�R�L�V��)q��i-�tr�-��j����qDM[�1Z�d�dU��,�c$j
�6�-)�Uǡ�VǷV)K�� �%S�v�y�g�Ș�s�,�]�*|x�ԃ$XiQ�#��j�`�69uM�U4%h�,��V�D0��H�:�Z
�t�5�唎����J�n�l���u���La*�(���r�|Ʃ���MK���i|�.+)�Z@U,P
�]�d����*���cJǣ���q��p<��@��yq�G?�����=/e��?��sC3F7핰������5N�RT��J���Z��kK�p�B8�Fj�O]ʝ�+5�g���sK9��q������݇��W'��1��on��wuvt|�C���z����<]=z���'>�3^Ƚ|��>�������ً��~Ns}|������ۣ�����������˃���#?����q-��ܿY�����=�{����X��5�s�h ��B/y���<�ZP���2!M���mE;C�l;f����Ȧ'�:	������H�H�}D��2�4��n����	
�������U���\D�0�>T��nEB���0�UQ�/�ɦPK6�#Hɗ�$&�i��l!
�$&���eL\o@}Ji�N�Zp5w%s]ݭ��v��J�O��8���-6��f�@�i$.E�6*�p�Z�&�#��qкIsDk�B���$�(s�lEM+�b|����.7)SfZTc��
�
Q㷇v�(Bx��ϐ����A�����iZ-kq>w��|I4V�
����T�N�l�3�tj^�sX)v���A��HQ1 >_(���Ւ���a��h�6YE#���M�p�~��_��&�!�]|{��#kU� ��H����~:FY�	5�CYrg�8u��y���wL�F����%d
/�hʐ���6��B��>$k�.�B5o[>��#,//���Won/7�����˳�??�~�O
�x�t��xXvp�}�N���zg����_�>v,����[?��盷�g/��O�����7���O��ŷO�������~����g?|����w�_n���Gۛ;���;;����_�����?�|~�������
_ksy�y�v��h�]��5�t|�v{rG�g7�ca��������j��`�tyl5~��'>���[o��|
���2��������AQ����SH���&�Sԩ�ǡ6�8�D�5��bʦ�ܦ���&Dj6#d
�@!'��q��i�mJ��M?0e����Y��9�9�m���)gJ!0�Sj�QV��D�pp+����A`�Cʁ@��� ���	! �!�Ӊlp�D�W�ȕ@cBU��r�M������V!E�|&�r� WŸ���n�1� ήC��ͩ�(�#�?-A4CΩ~�`!>SZ����ߺS����VjJp�%��ܚ�=�6�}��\��CR�Lf�t4)d*d��i�A�-�89�D�9��YLJ�]N;\,�u�8(4�ˢY?8���5#ʀB3
�f-L��h�F���)�X�F)�����)��s]��|Mi⪗Ub��@E��Կ,�_���~����f����׿�t]���?��60Yx ����ap�M�4e#�E0���H�x}��'UN�M�Ʃ/�Γ��E(�G�ɩz�T�M���h�u^�M�Cr�"�E� ���F��@�XcRD�Rc�B��"��q�u�K*�B���-��8n���=&��*����nY|�s!���m�5"@�9�	1�K�G����7�O�D�;��	<�&���`ZK�ȴt�ѥCӜJ�4�n=P�#t�D�1�m�>E�T%�P���*&_�@���>Z通��r�kF�����4E5`��i�!�%�9Ĉ�(3{�/4��5v�&Û��
hU�0��L�h#N~;���N ��|�i)��i{�������>�T	H��v!�����nE%�������c�S��@��4�4����������{��Y%'A>�l�U�6�:���(&�@$��&�Dƺ"h��0�H���1Mj�f�����^J��g����F��rZ�Ѵ�S[�c�E��3"�O�CYzH�D�H0��L��	
���h��ŀ���g��qM�o���^���֝����utc��o���s|��SR7�����|��k=�����]�y��Q��{wON�����p�^�����;�������v�������d��+�z����p}�z��S�W'�K�ى����|�t��a�p���~=��6i/�z9֟~\��޹��"�mY�� ]��/fܹw��ų��LH6��{�̧�'�-	�k����|���7�������^���x�ӱ @����r��n#:8i�9@c����IS�-���*�F��t�;C��p�SD��Zp's�J�	1&�B}�A��Tu���9���"瓭�J��1��˩+�-e4���ȝ3|�Ha��1�dC��"M/t3��x5�y��ˤ�$�0�(w�?�����勦_V�'���)���Ҕ_J�6���� �y�����\��3�m��%5���C��c#����S�]i��R�Ip��Ԙ�CP��ԕ�u/����M��U�~D�����WE��S@3�<�ۥ�.�zI_9"�3��:D@#�6b̄�D�5/�,��Z)p��q�˪y���J�&�UNT�Ԙ�#]5�Ԉ���t��f�O���H�U0�y��r�e94*z�$+�
�O5cQ��>�_�W_}冬���u+���'۲�hI{e����nW�hN�K��ox�����1�uYm��)��Ʃ�^HqP�GP!�G���k#=�x������%�'7����_�?}�o5�����ŝ���w\K�C?���%SG��6������_\��ݿ��{~>�f\1��ҽ�}~s������衯/�0�N_.p{u>��<�c�76r�������Z�������^���	7��j���
-g��X�r2͝ɱR�h��a�?�LT.3�������#����D����8�pw��Z2%厠�:���|�,>)�]���K��OVj�+�;U��ʑeu^b��v
�I��p�+'�g@!"s
a���Y��0����^�
�R�O��\��݄����Sˑ+�N��WT4�=a5�ì�w�TZ"0>�T:)!���N���h��Ќ:1
�e�k�R$��e���F�V���zÙ�U�d�Ɋ�c�t����A��)F��|�����Z�F��hLz>�4�=H�ֻt8q��,�W�1"hOu�� ��p�&��r�^��z����T��+��)N�¡`d-���n��6�O�T.JV8���B�@������4w�|K�:lQL�Ƥ�G��Ӓ���<�\b�9���EÇ�r�nLr�1GT��g?%��P&WQ�"�������.���p�ü�wzw��)������o��ֽ;7�C���/N��	���l�o6���\�m�.�O�/��'wO��֝'7ϟ|��շ�?>��l��o~��w�y����ͳ��'_����~����������n��ų������\���p�����]=y����ޏ�ڜ�|���Ņ�H��C�Ǎ��v��Gf~zz�,O@=G��Y�sϊ�cm�nJ�sW9Nu��v?��c��U~f�8��ivk�dp�e�zGA9x�/�z��	&��#��i�������hGP�c��,?��Y:+XQ���F>*�Zh�0���k �τ�W�jJ���!!pY��*T���O�?���O���r�(:ErB"kȗ�I���J�-�8��m)�,�g���IH?f��Ъ�}#GcMK���pQc!:uc	�A�*B�]ũ��jM!8�R���g*R���e����#�('3%;5}8B�r�UtC�� ��q'�X��?i8U��*�:��bjISi����4�Fk�����>�>�V�jjd%r�M�bk�����`8FS�ZFڒ�TTz�˅�ΛX�q0ᕠ��F�e�%£UqTZ�M�d$J��������DdS�i�;GPQ|
-����Y8J�g����̖�#W��?�.��͈���D�Y�p�ir/�I���,�!Ȅ��փ{j՝��V���H�u�,�� ��oĄ���%86�Se�a4V�'���X�Bq�����4�Ɗ��dH��0�jQ '�^ۜ)�We�"h��Wn�h�b�"BM���sCjI'�j#e�v`6I�_���$$ؔ�d©��g?-�4��gS�#]4p���D>M����[~S!�R�XW�����X�3�dE�'R�������_Y�=�����ψK����9��?�4k�3�Tˢ"�ߵ� ɦ0eçH�x��@S���U4e���eȓfZ��r��)��.)$�N~U�f��t�
NuMJ�֖v�D(��Ӕ��a�JW� ���
3�C��<$v�!)+gd
��/)'2�D�(�Z���|���I��R:����}�i�rcB(���$s�,Op��rL3��AE�+�׏J�8F!�x�$��JI�=?5̞�Gr��V�4����O��R.�ު�/J�f**����
eUK���T4AK0E����g)ah.WO�{�i�����w�]���P�I^�;~��h<��׽x1�������z\�y��IO�}ː���΅��e�/�^n.�O�z��ǶW{G��<8�g��r�����ӣCߛ�i�Uߺ�������	�
3~�r�
�v�h|����J���x;��Aל:��e����}�xgՉeW�<�]��N/�ܹ���c�Vk?8j[|5�x��i5~�fs{�>ٻ�T�#���=��}�Z������R�Oit�:�֌��m�|�/괱��:(�F��A�KAKӔ��8&��؁�$4�Ech�EӇӁ�
�UG�Ȧ`y��D�%�R[j���iXH�VM�<h�B6M��1�h���� �Bx�p����������ҏW��M2��Є�a:9D�Zmi��!5	���bS�@�rMk^
>5f�ȋZ��c:L�Tb�=W�Z��Y��
�~��E�j ���q���:Z�!�T��V1osɢB���C� ��j&�Uјr��B�4�4ʢ9%.�(����h35~m�3�K	1N��J���Q��VNzQ��FNLʽ�7���4JdBn}�N�f����T%_T�f����᳚7�ǔR]Q4��a�9�ڨU�6�lhJ���x(oZ"P��Kg>���.]��%M�+y��o����o~��ߍ0�����<^Gj�M�?��M�v�"(�^O�G[p#��8I!�8p��m/}����̍�<:���뛫��Ƕ/.��>;{���w�]�=:�{����������G�}���׫߾y���X��x�䫳�����7|���������{�����vs���W�.��sw,{�ܷůN�q��[o�o����:;:qLt�˸�{�!�:�>ߩ6���b�:��M�E��Vj���"�V ~SQΤ�a!��dq��@V�)B;?�8��~�ҡ��⸛�����@����"��-q"8���w:�)�%%+��r�ږ(���ەD�:O�_B���%�
Ĕ2#b�nd���^H���*�,#u2�@G��fD������FS���3m��đ�-���Y�7�`!�N�/Ω��T"͊j���Ʌ��o:V��*T
M��h�4�� �+�6�Z5$�|��    IDAT��L�d8�Bp4����,��}�����BpNS#�3�3�tICwe�LP����e�)K!d!8�*d��>��!*2Av�4Ç�ꔋ�.�L�M���w��1:h�P#G])(�%�\��n'5I������^�4�]=���O!���*@R�lV�=�-G?��r����S�_:����'���G!��B�]AG�K3�Y��]�����ԱgN�F�7���d�du��/��/����w��ooOWG{���ա�/>��=�����{�{����������ɞ(}���>���ӳ������ݟ����o�����{�ξ������������7���x�����/?������G����������~zy�Z{ϯ�y��;�'��`���v�MM?�y�:rf��o��*��u{�5��f}�p���ж,t��zq��vh��S�A�Q�mf[7u�{6����4��w:��4�C�ֶ��zWչ�<�����3d�	� � e!�"���Lkus�9FUZ5'�����W7?Z��n}�,A9��q�M)����ij�3��h"|:���be9@c��t�$҈P��1�设i��H�O�c��@K̯[!��J�e�Um:8�������hV��[>�)�lY7���̭�h��b&رN��D�Ё0��(�D�AjL>f�Tߴt=�G��
q��I�/n�?O�z@�����M[���t곶I��)rK�����H�N�)$k�OX�i�?S�v��D��qV%R	���I�+�8�NE;&�n�8��%HJ�h�H�-0MN�~����@(G6�B�%�U�gL"u(1�h)��fo|�8�x�d���$S �f(��ĉV�qV�����K�'AL�jAJ�\"Y\�iK4rf�֧Q:s�!�
�/���G�r��t�cm�mQ���E)sb&Xz!�%��Q�����;qz��orMw��PH���A�&�a�t:�z��Gc�s���ն�S�O�#%���G�[�D��L��͑��E�0)@V�1�����E(q�(MP2�꤀�]qLu���3�)s� rR8�o[��h"�G(�~��T�Bu�r��:�n��8���M9�8�� ���J�̨��e	qL�n��+$$k������ߒ�R��t�9��nX�QN'5 �`����U1��zF�D��,��&E���uXV[!�cEc�|::�E�B���ҫR����;L1�LL��#�\��LyN����ʍSW�D��%�,��q�٘5�O�-�׏P��B��=���ON!M�B�՚
J���f���gx��
b�f� �I���[�Խ�(�;O~�A�����p�h���X!4M\�\�����/��pXE���e�N�����'?)~Y4��B餀��<�e��×��_m��}��WTo_�jd׀:��zSԃ)�@��el��YL������>|�-����&]�q���_�al7�/o.=ERLҎǅ)<�˵�'4}����Z��%/�7�#ϵ�/V�Wޒ�������;��#�R�M����c�ZIq׻�{�ص)�K�|/����'����mLg���U�zuj��u�������W�7[?������5�9�rA�k0/���l3���8El��>�c�K`s�/��q���ٹK\W��o}8�9{ih�����'����c'�X�RX4�1R5+Q�h�����;^eu��\�h���e�	���2u�8[���4� K��5282�H���E�L�aeiC.?0fq��*ʯIj,HQN�:S4r�U�P:S\^3����o��Eo>�R85PŲ���П��\VSY�S:~#ж
!�Pj��Uݦ�O��FS�f:��#�2��|��O�f� �R3R����b�R�-nJ?`��5W'��C����8qhB�FQʚ����Z�S�> #�G�P���4)��/���hʙRR"�ճ(��f�QG�����re���ϊ59AE;�q���[k$�(k '):�C'���Q��;�B�K
�gȻ�gQ>��d�}dRq:	E��RwS8��2HS�� 5@�P�n���p�{��+�nѮ���O�	B|��r~��x���4Q��[8N[\����s�n&"Ǩ<�g�a�˓��a�O3�S@.�?Y�}�;���[�����n��ܻo}�����l�On�|�p{�ޛ�#��>O���?~�����������b�:�;���S'�����n7��n����ֶ>txp�@������O������M�vN<�z�2��`ܡ���e��{�k�1�^����ov�>��cg��,܁��B8�ir	�n�Y�t8�vR�1��{8no�ҥ���hj���?��p����wL�F��N/U+׋��Yt/Mc@#Ш'����ܜ!~������á�v���H�_=kI�mB{�Y���ɡ�P~8D���ܢ�O<A��|�/��0��eLٞ�eE�%W	�)�Yn� �J �FV]!�R�:�-OV�*��J8R�����>V]��6MQӪ(=�V�2%"�o�ʩö�h'�������@�PB
�Y|���E���1��`փh���3D�Z�H�@��42��su8-�TQ���$e]�h��(�*�SM��$~%��p�)�&MU�%kZ9��_]K�j9��A:�Q�}�K����==�9�k�w���@_��(C�1�G`�c2��>�t�dǟ��%�qH!X~��geq$6�d�U�b�z��˄�O��ܑ��3������W�'~���g��/��	�	��_O��	�}O�|[��%=T���O._<����?~���'_>{rw���������_~��w�x�������O�s�����������󳧇/����~��o�U���>�9���߮W�+�`���<~�/�]^����9����g`���gY�� >@�����_��[�nt��}��'�
;Б2B���%�i�F�4�D��]1���C�Q�=w�0S瘓�/��/�>��Ph˥����÷�Iu���)�M�ȍ�M>2�,#P��},F>�C��V�W1�,�ϡ<��_��XQ"I� q��U$Ng*���T%"2מ�����o$�!�{2|FJJ�(k-��������%�F�d�ʒo�8:w�AX��n N���8F����!S��vAD#`2L�J�Ѫ%LJH�Ip��E'y29���8�*��ѹ3�ǔ`ʁR(4�U��Te����i�1CВũ�����1m+�4�<�uR�l�4i��,
u+�=i7�g�T����L��	�~�-ZJ�6_����R�<���@ʉpj�ހ�C�Ɵ�:�sRH�\L���#��tD�Sִ;ސ�fBZ�bT��t���3�24��hC˅��[T�n����L�0�s����D����f�R�ґ���Y�(ʁ�r��Í��@��1q��3�����'�m�3S�ڎ�Ξg]|R����'h�b�NX(�T36R	)m)�c������MY������EUBnr4�y�g��S�j����L�S�Ȑ���E�eqJpf-�xa��(��I�RS�e'�j]�.n�g��7�)�G(�hi�語ˍf���S�[c��Y(S)�VJ�"�^���3q�#�K42R@VB��w��#��N��U��Nߟs����C�����hY"��J6fQ��|�7-��mE�p�˅q�,�)=0ZY�v�SW�>���r��s�E������0�E���ȍLj)��V�THt����S�/d�*a�̮�
��*�%��g��a���V�@T�+*�����aR3�OV^u5c�L~w}���p
�OM���q~z%��s��>���ݺrM�P]#�{N�O�"@J'�b�7��L��U��3�#�Q�L��r��FYč�yA3�30�=R5V(&P-|�u� p��Ưc�/�^8W�E�r%������+�Ѷgu�JI����W(��b�]z2�RJK��9Z�����v�;�F����^ySr�*J�z����`�9�pe����Ó������_]���҄Z�g��]������?0�-v���\=�;�X��O��CWvJ�o�=���������7.[AZ{��"�zI�M�Y�?9�*���WͶ�g��gW/�/�/O3��@t���;���<�[3�~+�Ss;�J����C��o���㽛+��܌�Lf�:�����0�p�+�����s���r('-����wV�D�T���"Z�F!�̝�(��Bn;���-�eQN!�?K��mͷ�zÉ�"~M���M����e+(��Q��g��o�4�+'��vۺ(L���k��H��\��US`+��5
qD�#�ş�Z5��JIߔ�l���DJ7"3�l����Cbɡ`�:"s�I
8���mR��PjƢ�X��p;q�Z3�*���f���3�ii�ь6�52��팱�p%��B�є����֨��.�\f�L��yH���q�x����>~LN�)�r�@�RQ���7�R���|4�v�bdբ�G0�S!>ӒQ'VAS���L28YM#8���3`�Y�q�U��{�z�9qSKc����d冘�n�p�s�,d#�Y��i��������^���������w��|����EL/7*��ڄZ@+7�`��L� jj��\7-�	77n��O<��g �+��q�������b�E曫��=�zs��{���ݜ]���¼�����w��Tpv{�y��4��~�����c���~��u�G��=:zsu|Mx��||������k�ͭG]ٗ�],_oMǫC�n�'�����I;�|nio��J���t������X¸u��;�-
���nc�^���4H#�A��!H�h�CnI��/��L��xR�W�]��M�������D4�r�S���H�BW�����+�N��o|�����$кh�(}�Yi�)�&j$k�DE �:LS-�1U���Hdo�Jg����ԧ(�H!GN���7%� 9�n�8���KNK���MmcE�<A�,~#q��#B�W�J�Bw.F�2���ﰪ�O����^�ЌSV�D�M��"<6D��m�sQ��F4����*B�6T���i�(dlKӇ�Zs2[���A#[nLjL����4���7��1�t��)$�/ћ)|�^H:^K�@�!�M�N�ir2K�H����QQ���At��g�|X�M��*ދ"�;B}��׿�5�,!ǂB��1�׃�1V�n� ��D�C8l"�L��݄��h5���BU�� I�wf�����ݻqv�����i���>���ݿ���;|���?�/���{1�n{��g�$�#��?��j���7}���O?~��}���x<���ջo�{�p��i���ǟ��WO/����޻wp���������ۛ���۳o?������<��_^��˃n�{���.�|y�_��8f|6����v<�O5o���.����x�3my���F;��t�Z@H;c�W�����9G���v-#H��q�8sd}��g>�"�����|í+P��,5g)?qR�Bl�^�y҄$X��뇳�`�e���Y��8F`����ou��8����M���9t�m{�Q(b�2��͊!M�ݿu�1s�r�O�Pʝ��h�ch��D"ҍ�g�.`�������+e̙�6��d`�mf"Bh
M}H��Dk2��wx)8pQ�Q�i"�5Ŝ���\H�c���H����2��gr�	%)�D��O>�M�)��tH-{h�'^Z�d�� �рN��[�nŘB��ip��4qc ��HI�f�gds�-} �*��t��q��85⍳
��gcKH��O�~��H:�U�SJ��H�GL��3	��>5LcU0[#�������͵$�R�j�.�����e�锋\��Bm��)�TdSS�M�X:g�WژM���sD���9uU{�8�t�������ϷR'�:�n5�z��D���r1嶨Y��JW��pj	�Nf��@jR�J������K��#�mX����%���d�Rө�.���"��nx ��$r�q)D�B�E!��U���b�p y"D�,�r� (D��h5�fj�i�D�9�1���v�;1�DD�e��j#r~Q�r��J�3!�u2���N����b��D���#P��'��8S�;.D�'M��g!"�u7%K�Ħ�pv��z��U7"s:C��MGn��0>0Z��P���@��"J��w��CL#G��%ʺ�(T?Ƣ��7�Uz�y���{!YU�+>DԨ��B�j$�Ac�Q?Ɩ��4&��Ʀ���aҍ鈚����.��':k�b*�uw	��,N���Sȑ>�mZ�9���&�i[g
�l��� �|mT�U����ȁCl�\O�q��^/��G�t��)��*���"���d����k�0��$΄��+�Z��D�Sf��|"��H��yx���K,�'i���/zd���4Jtic7��&v������{7�NϦ�d�>'��fu�t8�o#��:��J�;�E�'�}�WF����鷄�5(㠌�{__��d�	��J���v3^{���ۋ���;�ーނ��n��S��Cr�ۘ�����ܖ<u�G�:^���^�a8nn�[��v���#��I1����e��ً��*R���Y��C7(>׼=�^�|���f'o��;��^*V��-�����Eyu�1�!��׏#�9Ψ\4/\�"�<7:�BY�������y8v��L�C_.�l	�t{�t��F)1�����4guL�)���g�=��UW�*��2����LCJ��H��)�+d��>���L�ޔZѪ �b26%A�ܜBY�z�8���h^	cH���Z��5�,�?5K,%)#|}&�ǌ,�ޏp�*'K�a�[�|���%�
�r�X���@�KY��4�5 �ɻ�8,���B�L�t�ӗE�9 �P�ݫG�>�(˭`���0��ÛF�g��Ff���W�����!�n�A��I�A��-fuF%��3SY31�J;v�����[��o-r���כ(&'���9�d���������JC�3)F
��Z�n��ދ���L�75����駟�������_���.�q^֍�ż�I�ɤ%�F(���Xy��E|�ܵ�c������]䖭�y����$ay��^x���_�l�Ûo8����ɏ��_��^�m�^l^\�w���Ƀw�����`}�˗/�_�=�櫏�|�����*�k3���k���������ۧG�ϯ~��8�z=�E9��-v#�'O?�s�
�ζW��. �R_oQ땻NVr��8�6�}f�� ��Ό��."�El��M�%�a]-��nf�Jc��"d�x��Z˻���;�:MG�ԡ�;�׵�)ԉ��(W
_���r!�z�@kuN$�h�0)����v��Ek�f~)�҈LMn"�!������5\�NT�,�j[B�6��r���Q�t )֢L��t-E�h�c������0�%8"�9U$ncM9�Q0v�5�Dk�UG�T�,��W�&���Y+�����D"�#��\"R�QV�h^��/�����R%�j������JO�D#�3_���-Q�)5�p)�������hL�t���m���P���� 2��8�`�er�}��w��*pVuw���tw�e��ޔ���G}���4I�(������|�;Uo�8��8���X�!|ȟ�-I�M�b�k>
�#XN�EM�SR1&�V�ԉ��p�������g?�P����������7��4��O/o�_?������O~���G�ۋ�˭_��m3�����o��p�D�]��}7��KZ��O}t���d���~���?~r�㫳�/ίnWwn�m�������S_��:x��;���?{��7�8ڿ��?{r��O�o��W__>}����9�K��{�o|Yе'q'+/Ք�E�(9�9^��!�햒o�?��Nm�]m�L��xݍ�.L�6�4өhJ�9O�̓�!w�@2թIg@| ���@J	!i�T7��D�J1B�����)��HX�*��� �t6u���R�F)c��s�I��F���    IDATS(�pL3>�a�-�X��.I�nP�R(��S!Y�mN���>f��A��`E�$�p��rME9�h�(+��o��i"2���<3e�-~U�f��#�I4V��r)�_���j��b:sg���8!��b@ 'DQS d.V�*B�!��rz[Q�\&K��5�o��2^Ȉ�戽~�D��ʪP:B�mj���Pm��t��5l���Q[���4�P4�FӤ�p�1ӄL)=PemuG��'�Q?sߢ%�&�P���eW���w��(̢���1�~U� �U��3�� �*r��?D��O _"˟�*�w��m�(r��tcB���(�iU�P�c�`b��JT�ђ*8S^zRMCJ�
���!����3�/Z��6Ҟ��GZ����y!���n�n�o�!A)mg� ��
����)��&5#��(_z=�R�H���V��Nqf����cķEB��J?��Ƭ�4!��7�(�:�X�p����@%�T� ����0�hHd�Kz!c���(fˉP?���rT�I�Zt���@Dc��O�*����h�I��1�8ƤȶW�1�@c鵤O+ʱ��svs�*�Ȑk8��C/�Z2Yd{�/�]q��r���Y�F8>�-��I�`�I��~�U�jÔ�[Z:0�N ��R�*�hj{ZY�+4�Z�PN�S��I,�2zn�fU���e��|�X�g����j�#Pv ԅ�˚���(�\#)�A3�R��������2N��B�u�HYƦ�HL���̚���"�ws�#kI9>G�D6��Ɠ���uWB�0�h���e��a���iCVh��8%�pXx�#�6��d�������M_.Z�1���G���s�xG�c��t�S.\"�t�~����/1���W3�Q���P��tWH�es�q����%F���������N��]��e�.���Dq��x�A�M��U��]p��2H�]�w�f�/�ue�������G뽋���������_�z{{n��������\�&�ukq�t�]�g�v���p�7�� ������Ã͸������{'��o>������V�7��ՉW"-�x<��5����.�ڮ���:\����7Dח7^����F��^K섴{5�����q�ф{8������huȈ�U�$�,�_��n�8�#r=�w�kXKUAӕ���Q~����M�Pc�Lkf�.���C�\�&�Zu�+�-�W�Il70�i�8��8��v��:�&2�[�H���K���G���3�M#�$�U>�6�1!BScYVo��YG4�jaꄂ��E��D���RH�Zt��85SnDM$�����t��S`�t� kV��O�i��Of=PHߦA��8�V�VY!��#K� \�G��Q.���d������56u,J�	4E0�wn��p����9zN�YT�P�^��̟Qu�b�I���Q�Org���^������1����(�DL!ck��$^Q#0����bR�	��'}�׮Ӂ�d7�v�#{/���E��'bi�O>�~2�~������o�8�CI�T�y�B�8�L=r:0�*�����F`p�����4Z�ܝ@�e���&��� ��ï^��:n���/�]�x�/���7�?�p����{ǫۓ����g��G��-����|�1yssr��aWR^�͋����;�>|�G~|�������Gw�>�yy�u��J^^�9#��`���B�þ����b�7�����>4t�w�L9{����Ǖ�N���c,��;��Ԯm�#1CJ�2�QLց��� BJ�vJa��bp)\)U���j���])���0'D��o���p����F��ZN�W��D��ޔ@0j�C���a��� �ק6Z#G:���
�^��2�P-!
����� �S'��RQK�H�,�Ѫ����\��|�����M��#�1��\�z�Ƈs��趩�g"��n�h��QN!���/Ŵca�R'�n����j9�j�b#f�tH�FH�85Y�h|Q�u1d�,��B��(N�h4�I'�I�zk	M��RL�f�V'���P��f��pQ>�P}/��qH��t�<�māk.�>�IJ9��j�n5���Yw�
I�H�ffJ�-u�⻜�-�B�˛Z��8}���pR����;�w��_�����~d�>k��G��Jd"z���_�3����~A�������8�Ȝ�93Q��c��,&�������˵9{?�;<��\� ����������������ٙO�x���ķ�{W
�l�����]�����o�16�W�}.��7�>x�v�/���;<�n�x��ӯ������[����|����l�ƛ���{{wnV����ཻ�~E�#����r{����R��w��3����Tu���#��f�f7��C�G�jɧX_���6j��h�Zo�m��Q�N�y �8�L�h���4t�8��N�:�3���i?t:z`�;4�R6��D��k��&(+��/��ZF!V
��F��J��I���'hL9qS4��	�ȷۦ�P�h*�J�|��dgJH���e��Ǆ���jq��k$%���k�j�XVHS~��_4+��Y�| ���� �BF�csLA]D`�ޫ�$5��Z��SgF�p>�qF%�8D���@+��L�?A���B����)#� ��VS�D���E�F��N&_b�bʂ0d��q�#[)a�-AFEYSN`d���sӦ�\N��_uR��5j�b�3�������t[V)��+�p�[�AH!�o	p #kZ��e#����
!����@�)��J���G��.��l ^�45<�˅�b�W�>@��p��z�l7BDcB��9��n�4��r�"`�Sk	�c:��-��)�ll	���r�6�>���8��Eo�'�_Ef=#��1E!��'N�>9���S�Iά҆L���T�2���s|��չ�OӘO��i$�!R9���`v��B��Y�T�\)����1���c�C �Zm4��tԌS��)GcM�� ��Iٮ���8�i!F"�r�~�ZT�(f`՛B�3�4'^zRM�F���*ʟ-!����-��,H-�RQQ��� �`�Q&����!ֱ�� ��8�L/�82Ĕ_H��	��8�2����LK��ɖ����C�����d�N$�X"�n9tڙ�	�^p�8�qD!�ƶTh,�Qp �z�"��nn��`�(��c� ݔqf9�M1Gg��ik�L������x�4�p���L$�A83��� JdB-
ί�t�qR�m���P��'��{��9/G��&ŧ���5��j��^<ǁ��Q1���&I!���a8j���d�~�zQbJ�ͪ�D�T�Li:5iJ��D*�_�ڨ��4�l��ߊt���K�+��E���ҵ��GNNS�5��ݖd�=���/8����������M���x�t{qv{��>Ǟ��f<*�]���t���q����{�����K�w��y����KX�kxz�������{�.:��I7�G������#^��|�����5�Jw����8��o��=��מ<���S[_�t�>��>]y�u����{~��ՙ뻷���;ۍ-���N2� �����L�RM�TY*�:��0`�o`��+����]��q�\>(��*5))�R�;wǞ�7��8:�c~��s��n�΍o��`���Bܸ&�}w�6q|�};.?��+/���޵��7J�ML�v����қSڡ��9�(��0S;o*dc��<���:>|�;��Q���9�9C*5�*FR,)y^�M���M(Gʢ:�HivZƬl�he��R#���k�r�E1��c�i����
-͎{0H������,�t�~`K��VE>>��۔N�	��i"�Èd��g�8��Ӵ@�6�E��=�h	4e��2�S�_�c9�F�&�i��j��9p�i7��i��,J�H��n��ئDr��6B%И�jq:��85���gb"J�)$JD�,�B�*Fx!���k����t*��O5HkL����;jIi.*��P�ɏ�,�65��|nHLx �T��m�hL��uN'$}��p��߆G�H�Sf� ����6N��9S��EJQc>��Đ�̶��T�t4�a�#��Y]�!/`�K��'�|��ܽ����kR�����������jZs|���H0ݸ˃P�<�T%k�0S��қ=����0U�� P3%� 4כ���B w��乽�� ������Փ�7�{_}�j����{N|\���K�^_�z/��mzWһ?8�|�������}�������������ӵ�����]�vs������"��tmƫ����~��|®r��;N\���n<~��v��������8ˍn�̦�	-�q8-�mG�CL9�4��$��A4)��**e��o�D0:���xr��;�8��p��(���\��m��3�;�΍r!�w��5�juSo!��N�4M��5��\
t0��UG��á	�G�D��"������	SM��u&sB���%ҟ��"1�)@�6f�!e��!�K�,Eр��#|�8@R��r|`�;���\	��(�́�0SUqF"�%#��r4�,f���i��2>Y�Ѵ�tR����7&�&���7j#��qf6��,��|�8����X����,$G
R˦���eMg�h�8��"(��.2��z�����Y��k�,��5Ψ�o��-��R�n���%;HA�Tݿ�v���SŽ��_~�ɞ��?��O��o����O?�ԓ��WB��I���(�>C��#��2�ጟf��^uqR�%�2���U�D�Jw�c�n}?��g/8>|f)����f��;����������~���j���<��g��=?±7>κ>�����㫞�>v�G0>x��l��:޻}u}��������_o��_�t��`�����w?Oί���>}���Ǜ�//_?���js�����Ӵ;O�ܧ���z��9��^��r3W��qS7��p���S�ޗ�%�e��n�]����hw��wz8%�����bj���L9'�(&0\�<c!J˥Y	��n��1��4�ڠ��@p8F��NE��Y��Qȉ&T4�_��4dHu����`�H��dn-��!��rڜ�/q���d��ؒ��Hy"�V��ij�	Ĕ��B��B�D8�kE��:t�ь�Bd�&�cJy�ĩ�P�F�8�"��5��cT��l:Gr&e�'2$��BR�Ijrji�hۺ��Cֈ3o�p�)�(�H��)�}�D�Ҝ�MYu�B���Lb`xS���yQd�BѤ��G�Ig#2�q�^���5Vb���w���+!�T!)�"dF�7���C��4���#�i�X"2Z���3]^�Q�\c~�)��g�ń�c��uR�e	��^9�|!���_i�:LĔ&�lr�W@��g�LtN��_h�� d�('�_E��-�P_�cB
�K��<g�������U�pn�35mH����,�R�U4�>9����a@d�|���!�)Y�=�Y�UI���R�FQ�ՅpL�I�t���r��Is��RCh?cV7#�8&n:�`�F!�i�S�Jϭ^��g�Z)��C^��:j� ��5M$AU�_��?������_���8��c�b��G�1�ԉǈ���֛�8B�@���r%V1�>~�8њ�#�UdC}���^!Q��6�5�PQS�h���)�
�3 ��6hJ�f���ִh[�,�YV!#K�f��N�D�hSc�&�H''N]���P�D��K��)�~���\SY1}����Y��iȉld���;6	�m/�?oȥ�DJGK�{hI��kx����D�L�n�-D���U�� 3"37�'�,:��V!�m+""�1��h����j�J���}���<����~&�?��6ʴ��b�h�?�Ui��R�7\.��qG��UѲ⋚�T�U����PSH��'"�ԁ�g���ΊhS�,5�P�j_�t�!/�xv+:��\���]`���K���j���%������/��/�����+�hv��߸�΍O�� �]"v԰�͍/�욻���x�ǋb�ԮW'k���������Yх��_�x��~|�e|��۲���W�l�����&�Ha���}Mo�|��ʞ8t����>��ǈ/^_|�������������M��뚻k���K����6s�է�O�O�W>�{&}�zsx�웚��I;��|!��Y#p S[j��#e�*��j�P�׌%ʥ����Y���L��(Y�n>G�9"
t��*�TbmpЌu���<N�@���#Ћ^t**�f'�hR�;�M�p)�OSY���02�B��)�T�f� ��1���5,]�r�ɔH!�4��X)�� tp D���?_���ͷ�n���k�%`&�c�a�,SE�GCo[�B�ɢ�0�p���1�)��-�}0��v�(��b�hf	Y=��J�Vъ�qz�+}�h���RhJ7Jm���$�Ä4�!AY�12Q!ϗ���iU��|��7jI"|�9�f�Zj��I5;�l*�/�X
�hj�n90>��B���]�Ǭ���=�~�W��=圥9d;vR8�p�cOB'�a5B�6����s�Y�t4�Tt��5^oa��늃�^�o��H�0�;�0a*�J�aF�X\y+�� �L3gnǔ��aRh%@�h�),�&6��"�c�+��^�����6���w������w����_|��_|��7��!pu3�l��=~t�Ar\�}}���{���ul/_~�⛯]T�!=;^-��ڬ\��C�ѓ���Gk�ȱ��@��<��\��>~�c!d�J��c,z�dǕ<����ܸ�vL+��;��9��'|�ch��É����Ha:thf4�8J2#�i����Tp\2:��	:��C6Ĕ���y�J�Ւ�B�M)@�ֽ��[W��	���������LU��6 AӤ4 !5����D���Z�pj@z=cv�"�2�ʕ��!�E�Z�M-Ӵ-J_{���l9F�����o�p����6�Quk�L��erh2����ʲ.�uR-�C����I��˒"�Qzn������X���LG�;�V:~���+'�x�z,�׳�N���RpcKV"rmıƦ�((��F��h�j[,��N�4k��N{�/���$�Q�w\.d|�
Z�L�(��Dr4�����3�\x]q�r�m��A��>�����ݔ���ۙ̷�$�B�g�D:7�򋤘�T��!>Ĩ%N�I	�:� K��V� '�G(�95" �Iq
�9�HU4�*F��P��e�r���O>��h_�{9�}�������;���>8|�����L�g5=����=����^W����7�݅y�r}x�J���B�O}�{�M_�����ꁣ������W�Ͽ���ޮ����Ͼ�������}��C{����O��}���翼}�����/��/�C��WW>���<��/o�'M�;^kӐK�3�������x��n�����Ggn~�vL��8[������ut��n4G�,��GSV�m�P���^�ё������/Z"�tZ�i-�Z�ybJV��s *NP�X������G��fDM� s*j�l���=SBkǪk�V��B���z��� �@#Ĕ�F��\No�mf�¡ =�-s�B�K�0)5P�iK����B�<�8�Y��i�,>ي
�VoFI�(�MP
�rsL����i:�A"��B�D졨㛎�:���lQc�8|��uq��9����~�Y�q:�E�JRF�,yo6R��MֈV��ւY�epX��tKb�a��� ��*�!.Tz
F4�z(�`�G1-?�J'�6���YR���	�i[a�����LVb!)ȦNu#@�_-�@Y��՞��V��K4no/��F��d�`���|`�u^��&���AEH��\l:6�_
25HSQә;�8v	�U8խD����3�O�&�\x�_��9�����N�@�D����m�!F�����,��qL�뜃��9E+���h���SuNk1n���!��	N#GP�X���Y(���a�ā�é������S���F��\1�7H�iL&�    IDAT�mB-YB#�tS4=�m,�_�h��z��'Ո��d�k�B]q,���5gɪR�����'A�m�E��ҦB�)�N��������qBro��2˱��R�g9Hj)ȝE��1q&��LՒ���hG�e�S6�U���RJ�?$���ZFU�w�>��+d̨q�S����H��+�Ei�gj��-g��1ڢ��j)T�V-(�I�"(Wz
B�R��9�5�)~gŢ=�p�a��KG-R��%Ɓ�B5Rhfue��$K�$[Q#P:���љ�hS�4�U�>��Q�C��)�T�%��3w�W�UΟ���q"��=�2!H�-�()'$��r�IS15Y�&���SW�|�I�r��xNd��q���J�3�
5��0��覢V�+q�]ct&��Ⲯ�:z��Y���>!ν+D�u#�ؘn�޿��v�x��+��������C��������<�Sf_����뛗�\�܍��E�T��#��:F� [�Q�����7;w���w�1�7I�釫�>�L���=z�r���ΨGy��i���x�u�Q�n0�������G'�������|���}��{7���ظ1.�� ���������]=X?~��R�Wcm����x�����u�/�]�W];d�������fj�;�Vgs�@�Q�!snI�0��tL�d���z�Kt�0���"��j�D�t���m�E�/G��ͭ8��j�դZFSY��@�P��r�RB:�o�i�4U�1�pX-M290&�eoJԉ�,=pX=�X
��ȷ�9���72��U��SϪq�υ��W���l���DS�T{���\�)_u��ʔM�=��BFH�s-@��$�o�#�`�8�4�g�s�� �5��rDgêL�̩#�zC:���5IG:#kT�#�_E�Dx��&�Z��w B��8�Ј�1S>�T�tv���"$����G3�$R�tB��Z8L�]�"S�d� ��H�#Wb Bp�<K,���U�`�RL��[�X�P4N)RlBYF]�2�tjڰ�@u��q�	�ޚ�4j�8��hh�G#���3�����G}�@P�D_h�����yw=��g���*�mʇt8���kK��Zla=�P	�Ӛ�M�['5&�(��N�qOtu���`]��+�{�������>�sw������w��}d��^]�]�h�oS^��N��ꋛ��׷������|���~I����ū���Ǐ�W��W//��|����v������c�|���O�x�sՂ�����ݞ�����SB.���]���p��e�x0g�۱L����j���0>�5ڄm��Gh���\Sfo��dE:��P��V(d
�U{(���C�Gʍ�{�R��d����=���O����s�Fm�`�8N�:�Iʦ�kXzwL��o�t�i��ҥ��#h�τL;٤,K���}��Y���;����ؾ)$j�
��瘔1U_�z�o���6�X��J�
7erI��o�`̀	�%��'�Q�u&q�@4��@�TN�U1'�C���9��ҕ�|Q�B-��֭ބ�,�rF�8||�(_!#�B��ljtn8]U�;�u��,W��S�D�sw�	*�������f}�H'h��C$�^"��Ռ����-!mA�Z��P�|x�5О�	ajC���W.��7b2�S��?����%�p���p������6��?��s>��{�&_�B=S��63� !s��ԧ��3��pL['N l9r+�iӄ�h��VMK�!���7���׼D톯�Z��1o;돎��#O��|�ç�<9:ؼ���S��W�����ɽ������E���Ůn��yF�?~��������f��������o��_?����\{��������^�xD��w����O�:t͛��/������3�7�_?���>��9�q]��ޡ��v�o��Ƶ��|��37Q]���s�q�X��B����k��
ΐ6�2�^;Ю������.g���-b�I�IA�����"#2O�٢zp~&G��?����'@8Gn�r������*Z]����~u�u����CdLR��(�吚ͧ�DR��_W�|�4��Q���"���U$!��x�!�Ҭ���zEGnQ�d��� �h���1ٜmp��]J�f��������tj2q]�Ŕ�U�j�cjd���8U�,jF��3�4Hd�؎�tH!͹��t�#M\��I�KI��T{u(Z�F)tL2�,AN8��b�L���s�3a�q����@�3o݉��**����p"׃ߨ�PmC��E ���7��4S�-A
2��b�:VuH]ѱ" &��S��/��Ȁ��@A���P��e��y KXQ�R�;��19�hƺR��Q
˱Q��!4�
(��S�cʐm�B�,E���8I�����DӌOV�ߴ�B��p匓iZt������J�����^�p$VbWk{�ϷW�-�e	�$G">M!E��c5��ء�i�9�9rKQ.$A�� �8Y��i�
K����3dF��mE8ј�88:L�B1G���h��F>&e�\��F��4v6J�,a4��v���[<��J��*mԹ��<��!��G ���}��'B�V�TW�N��	o�N��HӸ�-�A�EC)�")�D&8NA�M婓S���s���]uj��,*Ş��խ�Ο�c� '2k!�Zc>����,}~��eEH�B�t�14�K1�1�s.��h�vVR��f6q�*N�P�쇓B��=Ӊ �6�_4يj`��p=W�_?�Ei�p"�r�HA���nC8	9�xj�R9ժ=�i�5�����X�y�T�f$�0YN?dh���S�Fy�qj�X�ъ�4]*�yԐ��ǱpOj�c���~��\w�="єn�P! MSUj&���5Ɓ[W͔��N�pF-A!]I7�jS~d#��ⴢ�4���K����T�4�T&��bB��r��_�J޸Kp*D[jq����� ,@ӿ���!�i�hꮁO\�]��uA"�����u������G';�������oqE��ը���]�U����~q��ng�5]��z?R7�v]o�sq}�s{���r����jo�1?�.��\��	�\Ht��͍�)���+��wB��s�4���}��\y����qѭ��4o��<8����+�w�y:���o�������_��_���\�L߅�+/J������wb��w5����o9mx����&�}�P��i��0�����ԡqb�u�Yo'C��`��1�
�5OE:�-�≘��.1���4'LS~77�Rr:ӈ����JC,P�h7%�j��FL��|�p/�Y�۲D�
�6Y|�D�|��4��R�u�a�%�����)�fJD��0�,WV�3����4�l@o�?�*B֋���`�Y�$"�o,ʱ]���R(�j~-a�d9p�RZ��O�*F�P��y �"k��e1Q�,5�
�[����wV��"%j�ݮ�p��"x��	��K�c�ks���� LbN͘���֣�B��(TK��9���Q�)�'���t[a*%$e`H`���T"A4���j���d|`)�{6`-�����Q� ��y�������+�d-�hk�t�Ƥ츐��~�����B���}�i�1��-OlR�;V�ϳ�Δ��z�M�ӉE��.]�,umaV�C]���,�6?��8�b�B����7v�hu8E\?`s����1�:W}�{|��?~��;<;��ػ����"�CD/���/V���~w��j�.�_ܜ��)������~����ŋ���W�G�ޣ\b�}p�z�~tt�:���\�x��4v�㱟�vf~�����}/
;�ǳLm{|��,�c�C;> ���
��$�>-�h�Vjl��q�"�� �+#�i�ɦٲWo�0��AC0�4;Q:	:����!��B޿ԉ�?�x�)��{��!c/��w:O�t�P�Bu�Z �s�N!2P	j���$g�QuL#�T����s���AhCp*m�[4g eV�,E.�Ճ(�9�"d�B�S6G{9�0�f ��GU�Qw�[ėF�t�����65f֥�4O27�ԁ3Տ�Q'��4U��8qL�p�Z��^�_M[�B��)��$Ҕ��Z�Ԇt|Scj�I\��M'GϥG0*-K�p��9@u��@ꤊ%�6Ȥd�T��������&f[�/*�ٻ�4�k�� Y�Ԑ�D���R��F&��V#��:!L�تxk�-��o	v�%���K!]����+�����wC�����#)d!]M�������i۸�Lk��1����[�oD#R�F�r�W-���_@Yvi"�^�-�2���7�Ǟ��_�g����7_�=8}�����]��y�;�>#��9�[O���o������x�{w��IϽ�����W>8������g{׏����=�я�W/^>�����������<|x��A�w�G�+G��˻��������W��q����gn'O����Ͽ~�����OO�6+?YⳫN�ծ��|f֎����9'���/[��4��J��Z_ȭ�9`O�'7Z��=df�Tavr� �%:�F��	��>$�_��iL�)��%FÜ� �d.�r�!�1�e��1~#����9���_��,9�"�*-ض�D�u-AE�-Mn�3s'9�i|©���D�L!�D��i
qocO��!�\Y�
soE��Ɣ���7�:ӥ�7��hD�g63K@f�u��`ҌS���F
��$X`�MM��%k�NJ
����L��?pܯ���c�
�>�}�t|�fŢh-��#�-R��!�YiSQ����N�3���!����S:��9M1�#�Y�hk�(A(��:�I�,��r��1��#�F#����c[�!�M����LA��Skl��#k�C����|�l���JR��6R�1�k��T�����1
�9� �iZ�tT��Dxd�h��4��ߍ�3m[�Z���!��ț{!��i->�~TW(��4����d��C��\��ω�e�5�ɱ{8g4kGV��8u,Rc�D$�(��1��)�� 8�Rß)5`*j��q�,$u	�̅�>��F:���v3r� 0��Lk������Y�qv++��s
I�T�9r�v����1D-:�2V��4[ �vu!���&�.�L�Y'jS��Fx�\ YHS>ΤUB�<�/��/�����D�����5��"L�[)g�\4�,f�����BI���	BG(r'[�A�:gf��M�Rhj��I���#�m
,�6�j���p�ID�����8Ir��HA�6��g:8�Tk�>�*ā�CGT�X���r�8�FK3N5ө7�dE�g��d��5fd@#Z��X&�(�D�|QN!�\�����ī���i��.�Z��<��+������!��8r�Z�W����A��kz��E���U[�,#ӪH�>�-v8⣥�4�C�r�� ]QYs��2H��U��������O�1"��@�i
Y��t��4��B��~4o����w��\�O)q��YT�;�b^"�(��}��E[�����?��(.����3��?�����c=i���(��ҥ�����x�T���u~s���ws��~u~�b���`�K�ϯИ�t��x>>�,�Cƾ�9�	�M�f���b�[��2|����}��/�x�u�]Q�?w������<8:|�w=~��x]�����۽���\��b��|5��ի�������ƫl.�{w{���^��۹;n/���9ih>O	b�oO�NTxGӮF��R���/�G����q�����n*ک���	@���I	�!JS�+��T����5�M�ǡI�&�s�@ӐȦUW����������8�8��T�^�S�äOf�@�t�� ���hߜT�C$F��cD��r��e-�D��mK"q:45W+ALV�l�2Bd��E��U%�GXQ��(S�V���}���Vd#CH�P馵�ǁ7B*�XQ4kL���a@4Q��h2&(�cʁO�8�i�s���Bh̋c0u��m~�֥�NvJg���w���O�hM��@���,-���Qb[�a�:�0�.�%2v��u��4Ł��U���h!t�nD���%�s3��t4gQ���T�3W!+M
3e�%8;���=A��k��E��c�tiTHݯ��ʫ��E���{UJx��|��Q7a6T O��
�zjTX����hݑ��x�tj��,��Ah�Ff��������l��e>�Zz�������޿pu��������_�s�٫����W'����>z��Ǯ�~�{���#v�^�x���}�����_�T�u��h��ო��w{k���L�ߤ��"�����.._�9��g/�<v�����_����ؐ#��7���Jk|����zFm����Ĳ�q���؜��6��sX�A��6m��͏�{���,�~
5�THE�@���w��>?�����z.������w@�>}�mp)�Lӹ��tjҍ���t˄��d�
��)o��jL��ղ�D�[Bx�˲."�ڢD�>�.�,�(�,GE"B�~�|S~��Rʢ̒2���4�-�`d����)2&G���c�z)��H�s�(X�QuRt�tЀJԕ�B4>��L���r�SQ�D��[`�j��dpS���8rE9΢aB�8�#�f�QT��[��$�B��E{�KDp�B!�Y�� �Q.R�Z���X�����B@��crb�⻓%�ǁO����hEU�Hٔ�l�4q���:�C�1�Z����FS8v����^f[Dʾ��'?񎦛�O-��ۭ�%�f���>Gt��k	�Mˢ3���Ą����|4fu�6-Z"hp4��{k�ȉ�;�v�Y���/~ag���qt�]���/K���s��O���w���/���V���24�k9)G����݅���N�ڧT��.�oW�T�����'w��G�G'�O=yq{�r��GG}tfsu����t����h�]�g�����G��]��]�_�����{?�����z����j�l��ć���y�ڻ����{��t<���^=m�u�]m��QN����H�I�!))t:phY�ڱ�o�9�U�D"�p��Nf)�P�(��cZ�Y(:C�_J4������%臕����.�oN[W��́�O�L����9�3kEN2������q���� ����,�zB ��	G:���i�M�md�?��h��˒�U	+?N��HYc!s��5-�N���r��Mb:c�Iy�xCh9������MV�TT���ENAt��f))G���$�W4��(�^QN�-hFI��t�R��4��U�T:Z]�B8-��"]
&��h��p����oD��
���r�8�&X��b8���9F����fL�O�fk$���v&�|L��!S��6�Q�`�8u��e���Q�)\��TB����G����A�3�Å���od��V9�
��>-�/�d��]����'��I7�V�~bҙ���"kDK�H�,R����O9��rL���2�~R��?�p����E�
QR\!�@�c-��>�?K����ϧ8�*=��?¨�TO��a)�pB�V��`,k��Z�]��5�qp��u��G#7.�gc�m*�D���-3�1��k!����������T���Yd�=όbq"�Z:���텘R�(�A���Z�h��F�.ј�89՝��t,&�C��;L�4�7��S��5,J�c�LYM~
!�|8��N8�c�؎�iu�ReB1���Q~i�R@�ND9Y�ͮ�E��.%�(0}Y8%��sE|{��ⴊh!F:��4D!�h~mT��=J$�,
�h��b#Z�E�?��@�'[�M;VK�h֒i�W7<��{��Y)B�
7����R"�sY�d��,
d���vW��[KL���|g]{��Z���)�TY5`GK&����ZR�y|8�����|C��TQ�ꬮ⛢A��kX���i��6�1�ڍb6��R��O#�*|SRF
��[�|�Y�n�)����;���3�T�@_c�[m|v��Y�
��I��UK/��Ey�s�>\�oD������ܲ;Iw��K{����������fp�
E>�{�G�,¥�<�����9>|H����/Q@    IDATF�|��_�
��Ʒ6]ػ�������v����\4Ϸ-}����{��a|�x�|�r�p{s���r�Wk�~��k;����3Ӆ�|^x�|�ǋ}��+���ý��'�N����O�^����\(i�Ή���oWw�6�_��Ћ��5�&��������<!߸��rf:�v�V۽FEX~'I#��i ļ��������+Y��w����,~7�y��.S��Ԗ=Os�5V�����B�(��Dj�D�L�$����)�fR�r���$+K�c�O����Ȳ��c����re!d89pQj�Ӷ���ƗB$�S�ڠ@�4�?�!�F�6"Ki-���f��%.1�t����j���-�Z��L�����L�g) @��m�Z;���gK�:��I�a#����B�f��R�&Z���
�b��h9L^��n���>�Հ��B	Y�B-��]��AP���ɌF���8�8Lz#2�2j@�ǔ�qMĴR�1�"<6'Sn�/����l	@
��J�̧]v@���lG&�(���(�a��k�#�mnjh�д�ɇ�e��m��C�����l4�^�6��;�u�����ӟ�t��޲�Mԥ���PLU�J��	�P-rD��qHC4g���9��S^R��}�=?*�J��޸G,o ,O'^�_]��3o���4����j��w�����f�����ߖ>�"��|��#���U��� =�� �k�9���K�/ov%�����Ѡ#u{��ե�^�ow�}�ǥ���� >24�e�rN ����pߜ�V�ؒ������:<B����3�I�Fh�!�u��o":���]�w_���w6���75)8KL]�Xȴ���3�wM�s��c�u��Z���R'}���~0�fL����@S)�'�nc
U%>�����4�!�(M��F�*r��pfÜz6)������産DӔ�Zo��0G.A���pd1��UP��o�CSo@��Ԫ����(@Z�,��Y!����LE[~!"�-�h;�ƨ�JW�'Pګ�Qu1,�#˘OE��Q{UoD�a�+*hlӤX��E�"Z�
5$�\�����+�D�Q��l���L)t,�%��J�&�á� gq����w���U�>�tSES���s��BV	A��q�YO���̯~�+����ҍ���k`i�ͽq�*-Z(P"�\�EM��ge�S~���R"/���+��LB�9��h�F�g�˿�Kww���)���U��<^��y�|�G>�������o=����~�q��篮|�t<���������<��닗�/.o����v������7�����ūo^<W]����������w����������ׯ<:y�to�J��o_��~�zuvu���+��_]���mM�	�3�냣����O6~<ħUW�w{gN�?:m-�����2��|0E0v{oi9�s�pYs'>���y�U:G(ĒS�s���v(k�G�SQ`x�b����(�f�w&�ج7[����[HK��*EU!"��ϊ� įz鐙�_�Ě7��U$���`#�� ƶ� ��'"�$BcK��l��O�6j2ec4|ʘu�$����U��o��Q���r%D�[�P۳��0�@#�d�ls�Ah�Ls;�i���mV��֤(��J��2��l&5>��l�U����¶�5P{UApz�Y)F�*�^�r��0Ӑ�j80e:@H)� �
q�h@>�i�9%��hJ���Q^"e�����_h�g���2�y= ���S�)�ɇ�+�_�,Lʹh�����G��fx"��Mw���9w�E���昆7
�4�8�㨕`U�8@Q>r|c��iƴ���mw8�iKE1Y4�\��]�C��69�aJY.Z�µ�p*�7ө��Z)1����Y�Z
��8�D~���Ǵ$�g�|��(�(
iZWpP��eVnʄ�-�!��c*��c(���ů4ڐ^n;F� �h���d��^ �4rt����Ɣ+-���2�&'���F GT�EB�ru[���r���H��TH:��ΐ[�Q�)��g[4>g�6�#7�J�,�6��;Ӄ8Z�F6����r�5#��p���E(�����p�(�`5)B`x�z��J��)Q���u���G����E+��/c���7�.���b��m&�ɍIJ��%���H/ʑ��ጂ)��[#�Om~{h�8+��7�[�%ت�8�Z|HS�BsK���q�[E�!%;!1�׀DA
�B8�ڈ�´*4w5P���Ȝڮ4���O�겚��8��n�
y:칶��D��E�3�#�F+o7ȇ�*�6<wnρ�FP@#n:{��M[i�2 ˇ#�m�����_	�T�)+�q\d�F���RY�m?}>�9뿏!�%No�����ȡ���$Z����u��i�c7Z��Zڳ��x+�>��hR���V����y�/D^]��s����b�'2�^!�lF+�ӞTv��n���q�w;^�]$}�qw��'�^��-Po�J���]�n<���N�$Le㪱��~VӋ!���^�@���*n��g�G&z�z/�8v恷%�ǫe�.����{ϣ�6nܷ7V����=_K��>�Y�/㻟㻭�
�>cl˼`��rI���[�q���r�iR����x��!�k�E{�@�|��H��Zvx�L5��h
�!8t*�W�sgB|`�q'���G��8JCj��19FdʢH��Ԍ@
5��i)|�L�V+���Me���*,��ڶdJ�e�U��r�<�ܥԨ�O��	�'$���WE
E�i���ږ�`�PHPHh�v+��Ox�:�r{e�b9�%X5q���$R��hM��]G�(&�TjCw	�#w�$��

85/Ŕ�R��C�v�h�1��vW��O��V'Xѹ(QV9'IS#Y�ZB�i!p�P˷(�v��<�R��?m�)p��EM�t`;f*KEMe�&U{Q�D�60M���-A.��*3k]6��)� GE��D1��Z���'8�&�$�`�5�5��|L���(A��R8����%:�SB�>�(�:y�����8��[<��x�W}�o���� ^�ah��⽰^Ch�6�ݚ3�S�Q�#�8�r�B@���c�d�67.����*ǃ��ok�0��k{����/�����~����O�]��>y��ёwAo7Ͽx~qu�����d�s��ۚ����|��ѱGǋ�����?�!�g�x������A�q����������WCwn��'�;�.�\|�r�o`��|�Y�p�G|'޲��b�i� #y�^H[a�f�цS�xdc�(�� h�Kplr�)�s�wnU��w�ux��91:���o�����]g��ĝ�����N��#Pv>�+Qm@����j
�P|-��u�R���'�)������������&�c9�)5���D��(�I��mTNh����!r��������2B�'��0-��XŁ�g�)D�a���gh4C��Hd��G��U�[4�)���x���_�F�DH�����X���jC{�(��t >_�S'|%]��g��pX�|��p���t�NN!Zk���	д5��c�ɺ52>�&�j�"Xc��v�`�V������,5! �s(S�t%�c�1��'��滉
��I��7��$س>�yҹD!}�2>��?���B8Mu�a��2�%�d��	i�V��oZ-:�#�Q"M��O8�����G}�M\��>ͪ��>{����N?���Ӈ�G����O��Σ������ݻ�����_��ܨ����{�/�^�l.�.��~��Ө�ǧ�N���֏���_<|r������k߱����ý�Ǐ������Ï��w7��_~����|��p�stx��{�����Ͽ�y�juv~�������[�v��_���"�N��>gk?�c؝�y��4�������Clځ.nC8�$�����m{h�A��0q��w� ��0�s��ʣ�,����`#p RL�r�
)�c�'ؙ��7M�S{h����0��4�	OJȴ�)L�vi8������\R�1!��L�� 9h��Ď�i�$�����tH��h	UO��V����-���(X��>ufŪ���qL�ʙ�@6����Y4d(��ϐS�JLf�M����L�Z�)����*���r|���t���\K�������U�q2`:��F]u,0�����r��n�,L�8����A��a6&K
��
iդ*Q��7-wrD�t�&J�(5��2~H�2S"|�����J�oE��3
�bZ�p|S���d4�� ~4~:��qZ�P)�9��Rf 3U"?)4w�F�§&.\���#�$r�S+C�SW|x��N ��Bj5~g�"<��FӢ|���m�q��McV�/�H�uѦ�8$�i����@��% 1锨sӐ�h�Y/)
Սf��G�3��2�cc&Ru�Y(_�gV�h�T��6D�5��:Z�,~�M�R������.�@��1����\C�p����?\zQL����8�t�r�ЌKpD#H��>�7�}����	ҡllu|N��f�&H�m�������($q�R�"�{zTR3|��9�c*�D��fHS���vi�?9���J�։��z62S��E���M(���F��1k���כ�N�N0���ۭ��n#@�*��3����e:�$�cJQB�_i B�Eg���N�3nw��\��VJ0Z=������㫛NdGJ���JX��
ί�@>�Y�d[Nj�+1����Hc�,"Rl,�f8���L+G<��U4��lg�L'�4ݨ�c�	֧*Bۚ3���6Aâ-�3����wn��{9�s=���A��-s6Po:��@LS���i�5J���F��o�X�))�D3���	UWWbSc�0Kȅ[#YO�)����՘tNdL��]-��B��&���3��&r�:?�9~�����o��~<���\5v\��;|(�\H��9]�u����kT�����=��z	w���(ޝ�٭�� ��յ�m U�cu>1�+%�.�}D�=6�=_���9|�l=yM�|��-zyXȲ��:|���	zw0�g�R�Xm���E�&8O�<���?����ǾuiQ�__���ϻW�wǮ<��w}{����r|�������م�'�}���ίw��b���$t����B�Q����DT'*z��:ʎfL�y12�/Z���@䱐�R�O綩�D4���$Wtl�bU!�8\�r�!F��FQ�4~-MY8N����C͈��K�#%G{n�4���8�ėH�*	
���AL�M��L+,Z��SH�t&G'pY)�!�s�B�NY|��օV�u�lE��/���=1U�1�fJ���A�1Y]����UBEUL�9��J4*d����J˅DV�z˂���ܛ��V� ��f�B^�l��ْ�%F����bğu���U"W���T�%�&�Zр9b�s�)59�P�0~�Ca�6d�*j��B"�-AJ��bjɺ�혐��� 0��D��de�4#r#����29�*]�4w����k�%ʊ���آ��NXd���S�BMHngcY��?��?��g?����h%޵rn��?AHϪ��hħkd��S*����,�9ȁ�b�LmQ[�\;�]��C�$���|}�;�g�|�������O/�N�և�/�.n7��/]�������_��哓���ww�r|y�2����������[;ww<�������م^������#����Ds>x8>:z�
���5O���U}��|�hy����]�h 8�!�F:Cm9� �FS:��AK�c�ڷ��E�A[v���X�pR��@����q�#��Υ@�i����<МQH�[�2i������
NE	J�U}���(0�&ጣ�D��B��>1�(���7ń4�.@���qTA�s�DN�D��LcUiZ��B5dI%�4}�ܸ��J�ɐ�dU��n�L	��yJ��Btl������TM�(G	#B�T��B�T�1×�x���H䔒�Q���� >�#Ř���s���-�2$&�T���U�:Z���ngR7�QKHM�Y��t(S豖�B��!߮�sʵ*�,�T'RBw�dc�EP�#�J��R��)d�Rcp�:�@�>�B�;y:���g8���`�/b��������������g�xoS��~�!���q����5Y��0�G3OA�\��&)�ijLjr�JS�R�Ĭ�JZ�i���rm)�^���r}vv���?x������7������yx��O��������_��g�ǿ���_��������꿸wU���E]��7-m��m��^~�yq�~�{t��zx���`탤'G.���?|���닇O�O������g�|��/�}}���{�~%z�op���i�u��S">����}<���ѕg��>�A��4�9n�����ٷ���؍vi��T���=2�;�<����"D���WR!��/��!#8q�
ۜ	����[,���tB��MہJ�@�VW�FU�����F�o�$b#�G��t�+mDh\4��	0�um)D��6�\~�:��iG_
?A|S>�`Y5� ,���5 ,������� r$g:<k��P4`�^��o{����̧� �rS
�c�O�*JIдu�l**�/�LE�:����fx� �,}� ��z�Ȋ�3e�Ec��rX�ɊS�d����Q�h�y�̟ȟ-��(5"��VQ�)�ٜp Y~Ѫ���"��T��5
�9��BG�F�P䦘�_ic�IV�3�r!��CD(P{R��u%EeE�V= KG��*E喂���å��tD#�rj���B���Á?��G㓲�B������q�,��,dJ�}�/](�lc*�ՃP4u�B��
R!~]����SX:���h��P��V�X�Eg�����y�8��Ա���aӑb�6�R��lJ�_oJ�v��1���hSS�����p��9��`ʐ3~}V�P#>g��Ԑ9@�����D365��d�f	��oo��o���Á`���4�������)�Jd�E#$�^)��nEk`v�I�#!���Ek��S�����+7�Ȧ5?s9��r�?5#�Bݫ�V=�y"�!&�~*�'2D��#��X�-�<BU�M3ǈ��Așc�3�Y�R/j씫R��e�"0QYQ�)�T�8)�g�,��J�����m���#A�q��|K����rPZ��eN���\H:���	� ��Xi~�UQ�;������BkL��*g�I-߈�9����v�N~�H=$k�B�F�)��<��i���"�5��1)�[�,Qd�"�r�+������q����>�U��)TQ��a�hME18U,Q�����
�J0���^��XO��^R��RqiRo^A�s��Xv��]h��m��Ls����㫜�y_yt�x��W|�r�b��>����͏��!�ڻ��^���b�����M��y��.�7ww��ك�}�����T���	2�%�}B���3_�,g\\�#�#�\�a�[���x�����f[͞�+�s(����?n1�n�$H�N��Z{�wB�<�����ט�q<�v��h7�i���jߗ���]�v�sr��Gj���|�s�w}㫮����v٭����ظ��'w��(wg�A�8����8���g� �C_t��ܨ�;p�B��,���7S)8������3�dA:��e1�8��42L4Z����܅������j��v�p)N���g�E6>�u�T���	������)EQdEрt�@��@�6^o@"j�f�85馲� 5_���[���q��U�� 7�B�Z�t83���N8�8|#3Տ�,���e5�	.���T+�X�Ѵ��MV.�1�'[SLx4KK.�P��W��5J';۫V��M�|���!U��,>C0VQ�r�d�v*��^,�gm`2�F%8)�u""Q�� ^{^~�$,�EA�AD�����*�I��m	���c�N�4q8@#\��B)�Mgە��|唖��,���p8L4�
�%�R����Gu|    IDATv}��HDhU�2J.7|�״��_�#{�
��������Ij�����vիR�u,Mrǩ�jWՖ��3&�E��1YS�����)����\\���=/?y�t����_}3}�/^~����ӯVG;��������_�>� y/�W)�<��ɃӇ��\���������G����/>z�����;i��Ȯ;�CD5����FZ/d�F�[~ n���B+��Bf4�D�L-�(�4��<W�*�r��H����\)Ȼ�u��sϽ��_D�{1<�K�����4�W{?|����W{��4���gw=<�o}q�v���l���Ի�Q��z��w8f��'Z'�/�����D�7����_6�E�Dl�^�VC�娇�k��Z�W��:l!�1&�C��uxKQ��F��4и�i>��c��2��6���~�ɧ��{�����u��1�����O�>�6!4�7�@�A����.�!P#ŮT4�aۏ�U���ɖ�:���a�YDܬ��9�┢b�	�ټ��%\Isj���&�)$�^��R�m���MMT`�p^k�9��*wP$��)�qZ"`���$����D��MV��dG�A̫���$eћ�8)@p��O��j0_�:p=[+�n�2<D/�t�)@
�
.����ƛS�!��B��h@�b�H���Z�fX��p6�&h�5����Z�jC��W<~�@x���,[
��Z=r�b�͡wS��~�������O=�[= 2��|뭷��Z�%��OJ�Y�tV�G x��t���adI����ק�Y�\���adGnq�3DT��cY1�4��t��"<���y��	:L�@a�8�������O?:���n����9y���˫�^^����+����zc��d�_��+��Q=��}���k�>������/��\=?s�����������~z��Փ��_��>��<y���o��{|.�g7{?\>�����'�7����/�����9+�!/�|�́i\�ё=�s�����譡۝��b���]Ԕ[�uhy[:�u��\��ֲ[Z+dx�V�Ia��熶����j�y�7l����0kHаDEU$�X.:���
㍐�<���N4m��!��������+@\���y+,��4�p��f*���	"��k(D=�fDc�����cP�W�>>\ޘ�g�'��\^)T���V9r��9��WO��Dp4���ij��LD,�^��y��.RI4�.Gaf&�,�1��,�'9�Yن�gTT�^�ƨ �yg��=ë'}U!ȫ1Z���,��/#2\�π�*�!�\�u���R���{��B��eTI��(}FU��\��@�qDx��	W����ǋ�%~ٓb7�G_Hʑc�y�E�T��jsX�\=@Q%���I�=W_+K=�+�DZO���U���X��3�+>͢� �3�3�5!j���3����(�75HIS6�h�\�O�(`���Ȕ�+�pV�X�EA7��5��%�0�D�b #p1���Ǭ�9A�uNMHӉÕ�!F`dW���"r�)�B2��@';5}\�)AdX4R�����D��P..�b�K79���,�0f���tj.Qj�sihb��Z�p5$�0d�iXm�����f�2�"��Q+\���Y �Ԅt���M*f��'�؉�@�Xk&�v^`%�\�&Ϋ ����pF10�JN�pQI��~�l�W�T�^�ո�z�V:�0.QLsl���@���Q ���s�\��FG��D[:F|L�c1k�KH
�8��'!M�j�HC-��t ;Y^�z`F�eAx�c�r_Bp��zQ�h���Az��HS���!UX���<���y3���^�DM��U[�l������)��<Kǥ��g���o����n"����ֈ 3:^����^�X4�¼s�Nu"J�M_T{�0Do:z��Y_`�A�C�-$}H��$�Q��O}�@���CPo+�H�:�`��y���S�Ѭ�@��\lYx�K��|q�^tWPu~uk�u-L�uG��MIߧz�Y�I�>R��#��r�t�H�>����R����x�������5X�GH�����썟 �X&��/�V��k�Ku���O=�����f�!�c^���֕X���;�.�(g9��NW��@��u�{|�s9)�[7���\�x�1>��9��J/���M�G~<�e#_}hR^����W���n��?ܜ��uu�{��OŸ<~��}Ph}m���.X;"��X��r�A��\��GP�*B� P���ُc�l<d�6ƫ��,�˷����1�4yE�!���B�eԗ�a�i5 �>Ð}�I9��\�xQBL�w���BЦl�P�@.�D(�n�C����֬!�8%2�$�R8�@���s�q�b�RN�qQf
�\Ea{D*PI)��J�
�Cc�58���k�'��ϕQ8fЬl���O_���ɥ�L|�a;;]cW�R����y%շ�pjlY��C�8�ؚ�XX^v�y�R��� 4S+p�%����K:g+��s��3�<��()��b؁�4��vG�gB\*���'�8.�\�8�Ypj���X�7��@�G_�6�-!EPȔe�r��:µ*���sɮ��N8����ĉL�� 4�4�xK
� *i�=�F�I�bk�.ʰ�Ơ��d`�ͱY�E_I�x!MǺ��n؝K6���+���kG}D�2��>�J��E�CM��^n�Z��44��%�|p*���9������0��rO�7�g������gϟ���{w_�{��b��}�޻{}s|���;�9ڻ�:����dt�/R\��%���^߽|v�����O�8zxxr~vy~����|�����_��9�_�z���%V�[w<���w��?�{��������/c�^���S��i�&q�7/����24.3�̎�7�\�e�/��UX��a��]?_ʫפ�oK9��=/MW,� 2@Ϳ����g�}��1;^��|��9�hW"�p��j?y�T-Rhd7��.3��G�x���.]���H:��ov�o�X�^

`�E���������)T$f+S�Դ��l"I�$"E��l-�f(/B6�>P�ұg����}�r|j�8�c
��F����io�5ّ&�!ġ&b��|eO0�a:��H�82������i2��U�Cؘ�*ǬH^��U�!��k�*lHGD�-�0�ˈ�!0�ٚX["��Q��NBS�:ͽ������dQ6r�5)e0��MS�s��}:@x5��
�@���� �h���R�X�_���h���J!K+`.M�Y�h��1E��U�lF6#[//��^�����n�y� 7���g*@c ����^�v6��r_S��r],�W��=�����_��g_~������������?��o����b���q����={���OJn�Vۛ����vl�k_|��3���������z���&���������w��_��:}��ɳ�W�/.ο\�۝'߼����O.��ݱ��v��G��1^zz�7��彨VS�۽�}��~��z�z�ΐeA^�hZ��i��ٲ�!���/��|��O�[�ʊ	�Gn�:)�"e�K:�tZG��!s���41����zR����1,$M.��]�%r���,W���z��;32(W[�\U�_Ul-{���&%�( "�B��K�zp��SU����4dܞZ�@�W��y���8#�>�䧯������@!�V����9�[CxI�g��@�f̲t��M��	��C!�	T�ae�e��
i��Ld6/ٹچl}������W82B���2�N`)�
!ŀ�;�K� ��\h��Z?��䚴4!=A����d��ӊ![�فS��v|˂����ĉl���H=&�fX�el����g����B�֋���K�.5�V�z|��B�%� ZRR3&��D�8!��	���b�2xat5QR5�>��8B�c�KH�����[1"������p®��;�pj�����S,�`�z�YR���)��q�!1�����KA!���F B���4L�	������D���$X��B�\"���� ��dķbJBP�^I���Sck�������$8}
��L��V)�!~kB�jI�V3�meCQh-�j��S�by���z�M6�4���[�6��--�TX�^�pv��$U���1�	]1l��R�B�\���~=�\e�/)W�#��p���a����ˮBR�Z�\�M��F�QΎ�f
�K�n�¯T:\�F��K�#��9g)/>&�)��\��b��V���Mm&Ť���
+�����7&ά!�$pUs�B�t2R��b[7��.�2��S�6{
1���\SA:ڹ���ʛ�$ÊO!Q�s�t�өN!i[�GB��O" �Z���d�-P6T0W^x�S�І�{�=���5A�&8
ZEi��_�S���ENG_�Ec��l�(�5��{��7��e/��$>Y�N��:]����i�Z�l!�k��pӏB��JӧG�����c�o8��~��� A2����9��$�5
T�]�~��&{����f}�ˊ.O}y��r3>��h�4��Q��/Y�m��������8�2�^\I�E���s������w�[8��Ȧ��c5� �-�����vܯ���θc���:5.������D7�/._/��ew�W>0��but��>�uI����G��Y�ʍ��d|=���z������γK��T�ۢ&�Gjܐ�eolƕo�S�\ZG���g{u�Vb;��0�BF�ˁ�4DK��}C�Ճ	�� q=0��#�!q�b�'zޞa)�{v#�)^��10Sf#�|�N3�J�] f.Lx�Dh��%5&!M=�~x��F����pB��lyє��+���i^<i� Rx A`Pы�� ���р��D�V1��+JvS@&�܄3��B�b��ld:h�b�K�-H^!�Wa���	!h�%n��]�m�)�M�畺�ri.�^H��h��!q�4ٮ�VLQQ�٬!P�H�&��,���, STu��dC���z	I(�]A�U,��(H����uS��"������0R֋��	��z���#�Rɖ���)�$��BL��A&H��:Ёg�Rhq�0��XJ�F�	��3 UR��� *5}� Q~.d
lFveS�_:���?�\U�[^�b��SQBe�[d!@�B�:�A�	�&��-���j���_ZXǈ�E~�wܙ?E�t樔ꐣ��ZW�"���s���#n����O�����p����yv�;dO��?����_o�vݽ񠽻wr���'�=pkr�wptptx���w�����@�_����O^���7�<���K��������_�u�;�=|0�K�w�?�����<�?~�z��h��=
�[|������������ʘ�ߍ��Rߔ�NGp�������9&�j�l6A�!�R�[��ld=�l!@E���kp"h\�N�m
h�\MJ�&��.]���>�k�M�N��x�5[U�8�|�����6�����̖k�n�'�
��¥�B�h8
�ۚvZsQ�X��,2�0�b3b�ea�y�zš6c_
�6�*�*�!)�,)3��#���5y��x!Փ�ry��'M��D�,o:�,Nx�*��1��G432/�A=>��*��b���+�+�!���	Q?�K�:�0��#f��c��F�-�^�ɮQC�&���
@���,S`�EU�f;���2�����C�Zѳ��!eCQt����B�Ԝ,-���D�µ@F���&�a�M�
��:�Rj�0pؼ���,��aG�ݸ����[�������	������uR�3���l|C���Y�#(�ژq"���M�!�V �X����D�M->;}^m�L�ɰ��C�h�N�k��=?'�������_��������o>���ևGwV_c�S�zgsv}�����������o=\����{��7{>z���lǷT�{�g���:<zmsu~x�}��[�����|���͕5o���?�������_�}���7�;O���Ov���T�����'W ���xk�W����{�_/��o`-u��e��K�V�*9R�����}�]���Ď��n�%|mdZ4{�����X�E�Y�/����E
��4\l} N!��b%�90�;CASXe$�GH�h��)�f��ĄTa�\��Y�s����=�������S����ĉFA� �5̘`�ʓ́`@�����5S �3{|ve�ƞ
�t"��ԣQV�2k@|���������O�u+�D��T4�zj[�@�Q8�A�YD(0�+�)�r�e���<C�,fզ�sWYx�4�j��l^�e�7� V��R�3�h门2x�N�\h���(.�h�������.���h1���F�|�W�,3�PI����Q@�s�+~q���@!q��75FU�WC�lC�h=H����*0�>�^C�L�\�
��Û�δ͚��� ��?��D3cR�2R�v|cVFS�Ɨ����lH)�����H ��#`ǅADcp1�"P�4D�� �K����Db�4���'��%bk2��"���Bؼ�Þ� Z�����z���U"��.He@��I�R� ��*�K�8�^�쥃��n�e-��ђe�-/���6�� ����K��1��j�3 1�C��"0��R :e��V|	od��8�G�f8t�A���Kl�B���
H��Ei,#>[�i�g"��Z��\!��0e�-__�?���E1f#(m��%HG�U�t���IMN̪bW0�f���&�ð������o�Ck�㗂&N8��ҁ��)_.|o"�t�s
��B�Y �\�jl�@�^j��PY"^n����O!��l���l!Ԫ?N�)�_jHu�1s5
����G ��n"l��hͅΞ�h߰t��Ne�e��lR������{�J���F�%}LY5����e��6������*��+\oc�]���t�E.xY����G��]sh.�I���pFv�<Fx!��2�Pz|��H5��~6�t&B��)ի{�1�8��@[tl��3����Ǟ������#����V���#?��iG�U���tU,�e�����|�r\SX����;g/|6��}�1�#����Q���)��+n.}����}���}����u�C�I��nV�V����	<P���{�,,���ƴfc�>Q��%c皦2��k�c�����.�a��{.�8v�f>�>�vv���ѽ����?������xƯ-���5�d)D
IW~
f,�=N�awM��-�����B~yJ�n��Q��6��`�������5H����CI�Xv ��
P""��!8�}n؊!8��^TF���۟\�H�\@��C*��T�ӭ\�	�,���Eo}◈-���(����s�tDE`�G�%�L�eR���6��U��qA"�T���M���@�d�]]!� ���&P�,z� 54"r1(��lx)��%C:�l������ ��ЩTD��@CMl� UQ�,VH��R���!74���c�R�B������[��M�l�(=25`S�P@Q�jK�X^�<��I�
K��&Y�.5S���h�a�����acJM�Wk%�j..�10�@~K$���Eq$��Wp)������OkC�wdZ�t-�QQ��٣��q,��Y�!��ġ��%]dF%l}�Tg���o��3�(U�����G��U�>���&C��o�����8+�rBr]RL�G�˟����i���d�U�Dd��s��<��1�h�v)�sƈ��\��|}~�}q�냙ko�q��GZ.��6;��ճ�{�e�������w���[o�UV�祣���_}��}��w��<ݼ�S����y�����<�\�&v7;g����j��i��Hv����]��$9��p\vt]��i&2vC��ʶ�khv���q,)�����ʐ2W����No!�=aC��o�p����6�����9����X��ND8}S0\���Al���D��]�z�#��+�;Z��E��߂Ȩ�Xje��C��-Vc�u�b��6
p-�(�    IDAT=~kX��!�LV3DN���k+ğ���+W�!��<�0�GM+#�rI�7}����e����31\^���I֐�P%�\)�#D�fUU=zy�N|��Po��Q��1�M #�!���
c�j�Ĩ�V�Њ�k��cI�yMP�k*�>�>|4���Qx(\\z)�*O���p$e��B58k4A��K�P.�E�)\�S���A߹i:�X+-���0p0�G�=���G�h�{=\{�������g�g��|��t	J}�Z"�%�kڭ����z:��5d=Dck�l��1�	�nY��@�mQ[%��5��(17ALQ6��y��͸��p��x�浙�����\\���c�ooǗ�m��������]���ݷ��|����2y��������8�<�����/���%�����q����5������������k�Ig����xg�?>��w'�|��g''��S�A�S������f|g�W�>������#�~u���w��<�l��5,�r��cᖅ՛&�rY����Pv�ճI<�C
A���uFv��l�2��4�Cv��\�A��X)Ƃ/gS.vǨR/6�ȼD��������ߞ�^�~=C%�PK"W+��\1��q���{�j��E�9�!�BH�B&�F�
%���k->�ߊO��͌Ŧ![H�˰p}!!j��9�f�ϛ1{�t�E/n8��튯�"4Q��\���e�_�
C�RT�4�>c�b�0�@H�鄗�M�z�٩2�1g%4�k���DR(*Z6/�e�L�g�Z|!��3pxy���MJcl�>p"M�pVb�PH9�d+����m�F+�2��o1Ӕz��x4���Lh���G�\�jnm�FO��ә�Z���'�~���n�E�D���z��&8k��9h�pM�#R�m�t����ĔB�y���!D�LN��b5�BL��ƞ����vB!�&��ZS�6dC�����S�N����j��H$&R�!��(�uc��S��G6Ĺ-��0�Z5 !l��-�_��(H��tk���J�S@������TY���s���5��Q8���>W� �d �!���?5YFI��E9YC���5H����LeÑr����Є7�*@`�)n�un(�QFLC=���og�̀k@-��t����2
!q���z���d���1�T�B��s5�@��׷,�6��U�o�iNg����[���%��;��T�T0����q�� L�p�`��1#Cү��VjSK��S9��%qM/��'T9�YC���v�-�4DV�y5�D��t�O��{��B�" h������ z�&]���X6jjȌ��i�����PT}����S�@C�^�y���}�^���hJ���:A�!z�^���=�A���0�B�`|�F�
��S��H��d˦�,*Y����]U��@�a�����^���C�u��;�U-�x���5�Q9��;��Y7���<��X�\}q��W�y!:^���7ݮ|~�OY���q��j��ӓ�ݍ��ޥ_��FJ�'?��2K��ݧ�G4W^y� �{��Z{K�7κƺ�zq�u��p����b'��.]m��t�Ք�s��u-8u��͇Cw�ٸ���H%*�Lwg������gƻ����w�l�o�=yꃞ{�Pڧˆ�P^��,ϕ�jm<�R�s|����`�f�僫7�K����
��^FY���r��@��E��i���[%/�!&D�c�zv�SU�K�&J���@!�%�9�m�R+�DT(Do�Qs�AN1�����#����2>e����@����{�s�u�1��jhz6P8[���g����5��Xg��B� &���y=���
��Y���i�"�ƫ�I��D���C��rQ�l}k�@��*�~R��XpQ�,��dA6��\l�3�H$����b�eO��BZ@����
������D���-#�d��d��=��z�.��h2d�Vv�WCe�����T /לl�t	׏�z�V-C٥���6���B�-�;���.^�Gk�4�ݫ$���j3�*'��6S.����(3���E'M.R�[C��Z=�t��,�3K #�2(X@}��M�!�ԏV��-W���D�k�C�;��"��ʼ� �Ss(�ejC��{�@cx*t"���{�Ï�x�+ϱ�'��^M�&S
ҧ�%����1[ [�\5LC����1qx�w\�%IE�ί/<���2�om���ټKf�}�{q~�|}�'���՝��xWۻ?y���Op����W��o�O�������/7/|M�8FN��xO���R�����������˯�3�p��������m�s�ۛ˝�?�)||Q���q�:M�C[�!&���&��tlAQ�r� �b��l��(ʪZމ�	��8@�i���G�.���Pܴ]�m���N�>��>�����N�p;D /�?���yʃ��W���Zy!)�EU���.������y+�ah��C�Ǒ�@����`Gƪ��>Da��\���&/D`�45��\%/�	/�&�P���&|m�C8W�
��Y��4ıt�@O�hB \RV	C:�ѐ)���!��(�ҡA�En.M�:ͨը0P e���q�W��l�E1$[i"���d�q�4�k�"�Q�����䕥���Bf�f�U�U� ��7k6}�cjRGf���AV��΅�6}��R� ��Ei��W-���!�D*�3�p:�8C��͝�RV��?��������"��������9C�G}�#D�*��գR���-{�֋Ň#�셣�6�,���
$�V^�l��'����hd��r��������붮�	9oLi�Zɫ�;�~s��+f�{�gWg����rl�~��?D�-�/�'+���2�R��w�죯n.~�D�{|����͓����]��G�=_|�v>>x������?�{�[v���'�\�����N?�^+:�{��y������ś��������]�}���@�g6/NN7�����[�9|LĬ�c&h}Z}k� ��{���8��T6��z��]a:�\V����(C�Q�暳�&4t���T���μZ�y������<����r��g8ʘR [^vò[��BP?��<3FӇHͮ	�x
�ԐB���3��T7*�"��@!��r����h�JZ`I��,��͕�
�+ o��S�D`��ZH��![y��F�gD+�1������n��WCH�\��s�д@�r�3�\lSKߤx��^=B��;�Z�R�Tv�Eͤ���^��*�,J�X��ѣ�AG+6�aL6o@����-Qv�2 �5S=H����\�^�� ʐ��%J+\jCZ��ST��#��v����4��d�5���# �y����S��ʘΐ[Z��)��5v̑��[|�5k�cʫ*?���/�CFS9W|`F.U5w.=�VHe�LP1��Z!��M_���4��;��
���j�JA`�"5����!y!U�V���Vm)JF��'K�ؼ�BĲ��2b�4�	Κ��a�g���k!2�RU��hM�H�e�#@�3eD^R
��8��K����>���>�q:�-�\�bÅ�YK�f`�S���Ė()^|+Øj����rj��AD��t�y�>��M��+	�\^�ʣ�[a�v/fQzC-�t��H r`�d����k���j.e�V�^l}j���!��i�y�MM��ϕN����p�f�B�!��ɮ�8�fʳ�������i�)�jL"i,j�~)ތ�Du.��G3M^�!���
Ǉ6��FP�!�����a���2d@����+J�ɘQiFNar������D�yg�$4/x^^á��m���
7Ě�~��^�B\h��@@�g%@C-\^�~.f���*���a')j�ԴV�!޵�V8[�_"�	t)��KS��3�!#0cV��ω���gp��Hޢd���_���j���ݯ.��s�ّ;�Wח�G��'J�oXnǏq�9��Z��t_�����nZ�x��[��������˽�͸bsdU��t9tw��]?��R����u*��\�.p�S#;�~�sw�h�{��w�[*w��>|puz��O���;v����u=��(���Ś�͊�� _K���������M��/|f�zs9,��q�h�l�>�m{�ȯ܇�`�ʍ�q"�,�W�G�{����j��᳞ג������^�W��㊴�s�,�^�:L�ˁ�xǮݢ���B.8��cNn�.���ԒZj���.
�'WvC���v��8�8�I
\�]�+
-e;��o	*of,��]�2M ��H�MYd6r���#$�cT�7�k�z�\���T�y��Y�\��5Q��Е
��N�˜]���W"yՃ�~��W
����YX�0}�l.�2Z
8Ӥ��B j�3��0��T*�FV�祣	��h��� ]շ,٥`Q�z�fPf�P���SP��T`��J���	�(W<5�G�\�U��2��1UC:4�!JƎ�:".CA�e��Ly�j�MI��@UA��U[5 1���p��i�,YH.vQ�3ksMT[-�K�`/�As�������歓�5��M�2�����8Z+���j�&�P^�"��8I14}��z�����E#Af���p�\��«�A�h�x!�G�%�\�� ��tkhRƱ��Y��t/�5mH��1��h+����=�q�e�n�͟�8���5L!�#3�*�&;��zÐ
RIRt\J&곙�X}�'�}?ffo9
7�W���G�w�߹<}�3W�g7~�y�����O|����⻯�����7^�����>������S�_p}z������;���4�D{�s��l����x���w������������u��#ߊ0V�}W+!�ɪ\��s�4����\�Y7D�Ƽ��X����X��K�:��m�� �ОpХ�����=��4v�3G�^k"���=��y�`8먩-� ��ﴬ$�Y-�a�x�._CC&(�)p��-�ؼ(��J�������̠Ps
�)#hU2��z�(����!M��p��m
F.�2�H�@̛2A����sk��^���� E�:�J������lF��z��K�CI3E�Հ6C`�ч�E���ͥ?ؒzx��h)DE�#�X��("�#��؞�T�餬6"�f�}8�7�J1j���ml��f.A����ͮ��咑o:����Uj�V��)ĄD����5.�N=��h�q�R[Cj-#Mo)|��"x�v.si����Af�tB��/���|?�_[$(0<}��Ws5���04��@�ZC^C�i�آ���t��d8B���\�cVq����e}�O>��×@hFVI��5�8�xt�������Q�������5k�����n�/S�V�'�<�NR/ެ���f�t���w�����'��gOn���}���ͻO����������o��'��y�]�K����z�Ӻ+�/"�g1/+מ�e��rg�%�WV�g�ݣ��/>����;.-�0Y}��v�^��۲X���8�=`'�,���Ax[R.�P,Y`�T/�?^q�LW�E�m�\��5Q�"�\�B$�R@CC*X=�ꊯL|"�S,P����g%�א3ҩ�p�(�V�=s�����J8�dټȊ��@���~��:�E^��!#p��k�Y.�������0W�[(C�,�T DKS��=��x+	�QH$Z�J���h��o��Y<����
��"�W�a�4Rk������L��F9q�އ����T��ʨԗh^�M,��t@�B2$�'�(��Ia�Bn���ϛl��)Tje ��U�o�[�b� l}ir���?eØ��Vs6��]�T1!�Ѧe�Ex���Lَl�lex�2���7�
�	
g��^� N.�hu"Tyӌ��P:��2���l��" sUpRzs��Y PKs�*�z��2z�U�
�!Dk5)}���{�b#r5̌*	���
gϙ&�/�����[��R�e႔�b�\	��-X�4�BA`k8E�"EC}���9��Y����	~9S�KP��DF+{5�,��C��@���XC.}�p/��4qvI�+Y��@�P��fJ��.��b�B4v�c�fʞޘtR��&���!�a����!ᥫf ��#2����Jv3�ySN'NʥH�]j�������/������v
�P8M�9�����=/�bDUFu�(MQ�$�U�؅2�d�+��B�%�oXކ8����<�y���գ������/j�G��xR�%J�(cf̀�(ҐaHA"M^�36�G�(-Μ~��\t��A�R��P1�/S�<�hpQ�h�txa�<�N+��y�D�X%�z��-��p=��e8�;@�f�U�k^v����/;�D�V8���d��aR�V��!E-���l�iv5L�Ԅ�ٲ����Za	gpi�B��)�d�R�E���ި��E/iez�_���"8�㳙��q��خ��)]i]�����I�l9R��y�>��K����<�S]W;�`YՑz�˶�pg�wI1�c߽|�s��Kc7G�v����cW^����+��Kw�����+d~���cWTV��/|=���;n��u����ޥ;�˃��F��qCE>�lim-�9�m�&Q[��Ӛ�^��^�Ƒp|}�սnE8h'��1�
�����,�������� ��m��Û+x�~���#�mஹ/�uAڍZ��%ԣ���Y��n�,]FE�;�m׎ ��Z��˚�hy����2:��,�>�K����{l=�]��U����*�)W�%b����@D^.=Z�D�R ��e[vC[��tݯy�=2��b��,Q+Ö���5���vUu�آ!dL��-��@\(�k�%5l�x����H�:!�T	\�LM������fU��7���]���Ԅ�O(����h�z���Y��CBA,2f��I���T�Xǂ��P�6j 8��3 ���p��,p�epE�a����NU	RjC"�ʢ��6N���ڷ�by�5������+�m
@:lR��q)FI\�K#ռx��ф��T��NA%��MM��4Y���׀�7�j��m�!p� UI�8Dh����Q [A렔�M���(^���P^�L)`v4=}�Br���G�%��D ��16�\�1)��;5�����_[��X.�-��?��'�'.��-��4��"���x�ŰE�U)�O��b-qCdհ*q��BK��*�t�V`ʢ暴�W������_΁�����ٽ���Go����G�⟽��[��>�awg}�Cۻ��ǳ�鋧��ݸ�����νG�?:�{����w����Gn��8?��5>��q�t�R��笏��W܌uG��rs���r}�ٿs���]?=޴ct�/�&e�Y�&�V�6��D �F�� a[��8�� ![��|��Davf����X[�f�3��N{Ws�_�����l���WJ��<Ȇß��z�+�i��Τ���(���n�LrWC�pd��YI�6�X^L�)0�J�-0��W%	�v�8�B̗�yŬ�U1�Դ��ĩXv=/|���4uv�zx�O\.�4!�[y�f
Ԫ\ߌ��]���3���/���BS��,)C�Tru��S�/A �E��Ðk�fk���&N�Kcx��F^��/J%���ޞ�l+�m�!�g.5j���eDhFV�!����D� f[z�A�M��z��3��2JJ���C�@Ao��s�)|��#�ڔš��;	��H�L��>�K
���G}�O�Ǐ�(Lv^
��5���B�� �C0B�zQy�9D��dg4k4�x���Ӥ�M-����64�7��3�'����4GU �Z�E��K�nc��`;ޙ:�l�=5N,������t�W�~I��ۍ�7[s	�N?��9��ޛ��O~��������őw�:��;����>�9���O��}���뫳���k_��?�W����    IDAT>�iǸU�,�VS��|����Y���������у㻧��ƛ^��̔[1��hf���1ML��z�Jo�����D�l.��^��>B�U߆a��#\�6<�
`k��4���3���B�w��f>D����	Bre�g#�+�,8�@xL���Uv��hًƘ`��D��G�x�2�d �;���a��"�up���I�m�����n ��lsdWXL=�~�)>זN
�4)���Ϫ%�� ~HӬB A#�m�!5:k��}2���#kRL�j�(�cB�3�����3�$�gTn��ƫ��[�B =m�j�p%R=����i�S�4�Ys"�#6��k)#0�5.:d��f��Y�j��$>�@}ٛi����"Q�p�9��G���F� ��z|�������7�Y8�ڦBxY�ӈY��cZ��R3ܰ�V���2j���IC������.ꐽ��*![
|6c��[�f!�0��� j����o7V��,C-����j JT�a$"��S^6�-�H������a!�����f��;I^3��2d�Px�z�*/v΂��,Τ%e)L������V�U3����4!eD��l��1ǌ�����b鰗b�Bie��K,5������~���Sn(v���1��Ҳ��q�Ɇ4M�V�הB\�h���Ҝ�B��N(Rm��E��B�eBjD�aN���83{FٓE�Y�'b��~�4�C�1���� D���`�>rj�b�p���I�!{F�1�۶K�x8�,)��4 ���![pq�adV�Qˠ��fu���P���&P��he
��#�e�n� �aʘ��3(����ې�%Rah3�9\xC.d�
`3���3ʁ��H��k�br���_����諧�8�$%��1�S�*mV+�p�^[�+h�����%B!͒B�1lA���p/0�<�B/S0t@�1��Os�(Xa�������7�9b
hZS��Q�e��@�����(�P�Ԛ����������b�f���G� {{,�&G��������t��8�h��N@�l�E�֤kCJG��eY���x�K�k��Oo���wJչ=��I�>�kg[�K�o��zܷt���������ˋ����S��>m��c+z)|��j��w|����P��w�e9(�e�yw����2f�!��;}������e���n�*~��ιW�>�y�W`�σ�߂�Z��d�k9NDGG�����y�5�V'�o�w�U��UI;j�買!�u���G�K�Bګ:W��Ɂ @x)4�L>\�j�ш��n�����N��?��?詹PV�v8�|��l[�����A_���UI�t�͔אWT��2�8�e1��k2��YP�\�����ŒeϤc�V:.:@'��\���єT���,�t����mxR�y��5�O�3 �U*��(��W?�Dh�*��� �lk����V�P��B�)�.��3R�2�V�rQklM�r��oe�m
@0$��%)�&��A�TL�����Z!%����)6���@��M��Ь���z�@��A".��\�T1�ٵ_�I0e��H���\�MP5 �v�W͘�l�*;e(���$�c�$k�9�p�]�.c��(���#�û[0�$�����d�T��M���j�kp��Û��o=�!�#d��BS���,o���O��[��A��#�M���$|��+�u��DyN�T���*t���O>�������ۿEc����;�c���FZY�c	�hT �0�`�{�`TP��c�3h��UO6/��t�cÁ�A�$t>��Ԟ��vg}u}��ur�����?8��x��ߺ&7�S�Ο��\nn�ߜ�={z��?^�==�������G��z�竵_J�:��88Zy��=�st����y�S3���s��6W;�/�]�~p���3��eǛ�4C/o��g��/1�M��������^=���E���_�n�,AR�h- �L15�]4F���]���δ0m���ƴ�0Kg�����CR^|�� �E��&q�hm9Q����d1ٵ��j�z%1�B�O</q�^�M���BGk8�_\���d+9��1���3ќl!R����!�y%jIiZg�V�%�e�+�F�Φp��r�[,5)x�Mr5k4^=�D	A�x��FA%3�e=ܓ\ /Y����R@(��es�Km���H���@:�z�B��� ��鴆ʨ��X=�*dk�T���*[OV�gV^
�����pL�z�R녫�me:^�f�.!�5�z����E�Py�tH���yŲM���|(�3b�	��4�����
�_K�R!��OM�����Mp���!�0R�ް�O<&�+>�zBp��K�e�:�l�fY
A��CV�&��R�`,�ZY=�����:��e��ʋު�۫�BJ�h��J�K/�.��s��+�ޜ�ؽ��̛m6�&��Ã��?y��7Ԝ�~p��~��Ͽ�ݷ�}������~|pus~�=��^�nW�^]����7����7�s�6�E������|}����;ߜ��i�^�-�j�DKj�-�!úY����Y)dØ{��[Ql�S�B�)�v8�e!X��Ѫ�0ACm���g��գG�����&��p��203�`���1��3ʂ#*&$q|Q�굘�ͤ�]���T���؆�.>�
s1jl�E5C`e �_ o����O����
�j1��ۜ�j��o�M}�_vR���_�*�Dc,cS�G�υ�UPHy۫��\���V�,�g#�dcָʒ��G j�\Z
��z:	���˨}��ƫ-b��3�,���S3TôO<�7�^"����U�>�Q��IH���6�>Y�fŀzvy�C!� ���l���I�D��t�'���Z�vܹ��k(p�BVa�p"�WoLSlHLCv�e7�\����.05�B�ڜ`d�ɯ`LH8�Z�ϩ�jф�,Q^O�a��Kdc��gƐ^� G@���'�b�U�U�7̛�^+E�� p w��a|�!Z�/��Ȥ*U�V�W B᳒R�'XW0q"��=��j�x��)@��4P��]X��ök!����@
l���g^�rU6�D�Q�!��\��8��̫7TU:µ\��X���t��hE�ͥ+6B��̳����B葹�o�T�!\��<_=�!e=����t���.#NC��~T'o��2�`5��i d׋e��Hm�2�ͫ�"��Z�l��
և�#ς#���y�o�D)Hg8�DhH�P�%R�֜�������̋<51����c�q:�*���ĩZȴ�
'�U�@Ql��U�~zL���*�a��XCO�l��>}���������J�|����I`���2�e$���+GH�0EAMǐ��0�~682)M�s��\����S=�[������w�"�U�T}�p"���7,��\�Iq��2P
C"�2ri@!��� �M�Vp���I�F6/��}����^��z��&B�uvz�﯏ϟ�2s4�x��W�������rx��z���5.E�4�
���f曣Ƌ�eC�s(/���\yq<��߼���Jv�A����1A��W�V��C��*w����������ڜ��_��Π�������b������5}�s��$co;�-5p)�٭���&�GG��#7I��Vm�7�/�.�|���D흝��l�㻗l��p�giLa�0�\��K�˥6�W;��#1�P��i�T�:��:w�gI��fX��5����J!2o��e4�쌥�q<D�!�_������{�-��N�}�����Ԅh\^�3��%.;�ٱ;�^-8`T+�SOY=�(v��.iV�[�6�ؘɺ�U11�.\�N
���5P"���1�WˋL����w����n51z<�tS�N��Q!�pH��*�� ���H-jV��	@W�p�ց2�v.m�B���h�MGT�d1�x5N�e����3<Đ��P�ՐZm!��

#��k8
�K�
��A�wƿ����������I
���gR3�,M�����Հ�U�leac�`fs�E��t�hC��@L�m�a:��]����Sy�B��x4����Zm�D��Gl��-]�t�������V���|��3�E�[4%e4�	�.\�
Ȩ�)$�jF�[��!�"���/v%-5$MF5�����=���(m>b��M��8�̴�EP����� 6�uS���O_8�('�������"���B�j;�"DnB���X��Q�@�Bhj���7��O0
]���;b�.�\�Œ����O?;�{�W?{oy��v>z|����{�<z�5?�w��٭�Ջ�͕�t玳b����S�G_|�ͽGW.P�����';����Sk����>�x��]����ÝgϾ����b{sי�`���W�E�D���O
֛Z�0���sαa����C��p}C�6�#��6��)���͛�����������9����h���a��@S���z�*���,M�H��0+��lqW�&�a�B�@�hֲd(>C?��# �g��5��g����Z�^3���5��6���v�!P�aa��!B��/�F$)8N����<�&�A��p!!��Bܱfxe+R���Rj35#B{3�tj&������	-}�\1���6��O�&� h�j���㚾CF����]�E��"����P�l�{�@��P���,ܳά�H!騇��ԣ�V �B�j���I�D�A"^��U�����P�-��������2Z�B��y�������G�!
F��l��@���e�8e�Za|��z���5Ű���h��0$�f}4������9@��^��9�\@�X&�C�i��c�+êj�cmᦆIV��S��mP�����(���x�utp�%�7����v��6��ƻE�����bg|c���������v�͖י��<T
G@�(B��V(:BR����Y~m����P�V��ZgP������x\��X��g=ke�<�����}..?���g���;<<y����O���;o��}x�����_���>zq�s��}����ƭ�#���&�C�۟����Oh��?��3'����F5�m'��\w�����ԄYa��Y�ׇfɽ~q9	{�[�"0Z4�ƅ�&��Ƥ�!ۺ�h쎔s56=��V���[�:���C��#Gc�K��$��ӐB8C��^��b ��D�yç�#��Ѧ��/2c8l��U��< |D��"Mj��訶"!t����TL����w	���V;!��7�յ�)��S/�b���^80�J2,]�b!ڮ��%µD_������^�\����˦��\S�CN�pR���@��ǀ+@O'�h%�k����������B��������M�Y ��� ��O�#2�Ŧ�A�&�h�tJĨuN(<;|�&[���\=p��e�0��2�cUMI�omD��/M ;�>\.:z����ϰY�l�`�(��(P_ޢ��i�R�d��i��YU��L��reLvH��h�e|c�B�,�\����[^Ml�Oa��[���	ǧ�`���§N��@��'Dʕ`�@L�46��ʮ�x}
�/D��MKH�q �Mo��;=�0��8S<}�V��(�
v��+x�f�S����l^H6����Z�^+
a�l8YL��z�>f!
�!�C��V�U=4;���ȼ�qJ
����T�a��!C� Db(
�[��'����2���V���	�����cR@����b��2�1�p��SL� \��ā�b!I�<��q�8�h%��d��Im����#�9z-C��1�e����D�5���z�UY`�\��o�l8� �ml.�I�����6qLQc��?{�E��[��\�75�c�U���@}uV�\�՚�yeW!�*dkՐk�^�*d�ŕ͐��솕o(P���!ҡ��.A6άdKW�\����!�dSfC���Bc�y��(�K�.C����ͫ3�l0伹��Ee
e��P�&�k��j
�!n6C��l�劙]ϫ)U���0�g#�������>�w����υ_y��2|�\�S��j����+���Q�����'f�7��Yu�զ�,����WM��#��Ҩ����汬nOn� �c�v���
�F�,W�X)���"��PX�"��k�}���y���{�{�.^^���/����x�j���1P7J�y��x=֭P����ZG�r��u��U�U�3޿��{�/�Z�������վ�]��5��WG��{�wx���)ˤn=�v{��IzL��<�U�V�j���.�O�V�����4-^G����9Yx��NP3L��ؐ���_D���Է�"����4������ƒ���" M����s!�KF"[]��q�3��ھ[�६I!uv)��9B��S�!.C�춫kY#tِ�\��I�B��>�Dn��,_�&�V�{�B�O>����@�c=6�
�W3P��a�h\l����L�k�m�ë�k�6M=n}
T0M=�?����������ҡ�畔T!�p��6"�������-bu��-�x��8�C�W�W�j�D�	g�����m�����~�dwՆ��^%&��e��ݚ�Z��B�����h����X(��o�4��,��nWx�ZIw�[�}w��QK���A�E����;Y`7���{UHa����i.	�����!4�!������E��}�|��L�le�.DÙml�&֔����F/_�ފ���\�
}�GS�[�k5�Q�2�jʘ�@�^�)�ji�ʧ�@�2���ۄ�6�W�	���G���ԓ�o��nn޽z���~��'��w�=}�����ܜ���_�{���ݫ��S��>t��ӳ�#���On?���^y����W�w��_\_zö�<���س���^|��k��vJv�#o��6���t��9�&�lS�g7e�)7�-Ē�7�VU?���I�"�b��\�_?�h���H���]��q�����͏N����['�g�
�!va�ih�ؠvǝ`�c8�z.4�����W*���6Dh���c"�h��!P6��v6�"�`F8�� ��lR}� lb�ˆk���".WR\��`;��p"���dҤ�@��qio�+u),Ð^��b&��#}!Uo�:��7�L�*�1�Rh�z��hb!%b���6�� �3~�%U)�
���\\�R�
D�si��bB��%%U���*t,���V,�7Rl[�P^������A��2�V��84sA�Y^�k�j^�����P����#��z�e�i�&��IA�d\�-)���駟z�������G�f�f�:ϨrI�n�p4F}G����23�ĩ��MiI�
pi@�)��`ʥ�,&����jżdܮc# �L�WË�����Yb�'����������rp{�������>u��_�:v�7�����]��믞^}��Ğ�Ø�����I��WW�/�=��偿�������Q�������S�~e�Owl���<=@͇�nj���~������p�Q����Y�~k�*��ӭ����a;�n�3��X�VIH�
��BY���G�Һ!��������2�C�
ގ����.o�LRaCn�U�p=D�����#�6;L�����Igz���cT00�f�-�m��>�đ��0�����bȋ��gW	okȕ�2��8Ֆ8W����('����!�*�)�p�V�����T�F��s�ؼRH��Q D�<4��W.) �8C�5�hbj�l 6^x}�C��F�h�:|��A����&�A���E +
S�[ ��G8���!Y`:#��e^%��i��؊�,5��Qn፣/Q��jÙ�D)v§���ժ\�V�"фLb��К&B�j0�����hi��]����u��*{Z�(p�б���3dc�"�NlC��Ȩu,�u�CH����^xE�C�fU�<+Yj��)2M��g3#�pv��T���l�R��ښ��B+;�f�\vCᘑ)Cأ�=�@v��|�!��C.�f�i�=���7��q�2&j��m�    IDAT(�W����S���?�7�`qz�f���\�ƢI����0C��k�z���¨�]{��~S���1�
����
N__�݌b��*�W��ݒ�����]�!�
Ԫ|4�����q)J_٤� �����C?\�B='[��ɦ��!c1��V,��@��r�z�%�۲��%g#w�0L䛜pKAd�l8D+���w�D�}���Y^I��R��0�Ʋ�����0�3�b�Υ�+�:��@j�'n?�mS�Y��-CK��\p��Ѥ``jd� h�3hj��Ԁm0�Av��X
`�K��O�!�b����:|���a8�]
x!	굍��mL�';U�{u}��|��f�GJa�)�h�m�q^�N�=�i�4���Ɖ?^��j�s�%"R��-�P�u�ΐ��4M"�阬���gV&DF�\uw����ѵ��>:�%�\st~z��_���6e�i]��*Y�n�����<��3��V���1�-�좭����gN�'^|9����'ܻ����������ѳw�=�y��������;_4��#�f|!�n��NO.�=��ۖk����*`�R���?�~��Y�Z��?�O�(c��饺����ˋ��)�?$�#��k�x�V�E��C느)lK���ɾ]�����W��,Zsw-�6TP���ᰅ-�7��K`x!z�цbKb"I�=��5L_A��?�s�w|_��� �O$R�3���t�j��F��6؊�I'e�M5CW��« Mv�u�f�V���mE����^�W���\^�l�!P0�X�	4k«�j��(��k8�eM����D�s��_��H�H��A��;_F�F�)+�,��u���R�KhC���Av���b)�2,oQ�p}Ӭ���
N� f}L��@�lR��@'=_5��B�
�����9�].�����!R��O� Z�G!�.�x��� g���&sG�fq�wo݈�\����Q��t�ݪ�l۩ީ�������D���PV3&�(��A�jŦ��h8�F��	
XR��еq�8&�,���ܵR����}�KC�bEeX!����̗�G}���OJA�:�v��*&-mյ����.u��k�\Z���j�8�� 0AY���ϩl=�2���<^+n7��{v|v��t��/��>������sz�z�y<F�l��_��zv�j���w���uC��ѹgƻ��t�N�;��μ����œ����������t�]�>?>x�������g�oy��>��s�9��U�jMmU�m�y��A��zC!MS!/Doer�B��YO��7ϊ5L0Đ'2C#�_�*� �+�T�]�U�5
W:;��X��!)��S%��륶}���C��f!�lU5�Ѐ啂�5�U���y�\A"рͮΆ�QC{OF�yU �F�pA�(�)��%Z"=)L��P�a3J�0�W�ld.H��fh��m1\�ټt�p�bC�@�V��������Qӛ]�w�Д���1+�YpY|�ư��F�}��2��"A3;.�]jgF�0xs�`�	n���p�8�*a�E֔���!2Ľ|u�2�.���W�����4�n��p4C�z�!�8�"8e�I���i*/6���Vf�R�֪��`�?��O|�ڏP�_�>��7��iГ��+A3TC�5C &��s#�o`����	�@xG�DqƎ�Vdy������rSc@bv,l��ǧ`�X^Ɛ;�.�l5��Z�´QN��>zx�����cz�'������ɳg7W��=x|��`ޝܺ;�w|�Q6W/�.���y�ܥؿ�:<��0�����s�{�&⻚���ngzK���4���c">t9��aB&�,����Z�۵'MJ3Yͤ}ÙZ+FG��&6���m3���",��Я��F���W�Yg�f���F�l�E�~�*�Ta�����D ���e�5�~��3!�h�ҵbū�h#2��!�r!��e˰�S�pmaCxE�I���s1�赥Sk���HQ#9!\%�*W8���Soe�@=����V� 8����BD��@mw�)W�-5��9V*���脋Ҧ��3e���)�J�6vQ��zv�2�X��ȫO��6N:����D@M1�W�>�X��/��w���RI�����ᚹ��,�8��Pv-��p�P%C����!
�R�t�2ʋ3:@�ᰇ�H�a���l�!%mȖtd���7Me0*�������h�p��!��d�hM*\U��lF�S�fTv
�p��Z
p�̚� 2o!�&X�3�S(V��a���!�FV�j�c'���D�6=���N����Ȑ]\���g7$-D�zI�,)ZU1�!�hY���<�g	��@���q/������*;)�95���KOP��?��X%x�zH=<٪�s�ҟ��rY��OS�oʆ�1�3^�X��\��E�>2&��2BJ
���Z�������(@J!{� 1�=��UB�B�0����f��i���@��0*5B"�l�Ѹ�����1����z���/�>#}�\��rM�d�wנoؒv8p �1h�24d�͗�WȮA�`[t�m�d=�D�!iN
|���4�!c����U8�p!���vk�T����Y!�������m7����8D���lm�
4d�5�X��Ԛ�MΥ�G^o��зr�0Ҝa
�eD��h���SHy��b2�Gm�D��7$��r^v��������YR8z��q^ńh��a�1!�ٝ�3\��*�,>�	1d�+�!��%��&���	Q����k�
��hM<Z��S]k�R��s�g&/.Wv��o|��J��w�w��*�a#p䎟�v�<��@�F��c��Lb=�v� �s�<��=D)�j�|�ӟ��mNZ'w���z���R���z �Cw�<'��˷�O�~��K_��5Euy��g��[�D�3M��L����m����7������.�e�=��m
_��tp�깏�&���}���G�^�����нV��͛�wA�]��3�^R��g_���ώ�t	��հ��ڭ��dl�edhʋ��q�]k;R�.L9���<���mJ�/
�ߏ���q�.�ҴJ��]�������ZRh�eQC[��F"�h�_��8�'H!������&Wo
�?c7*r���G�a٧x_,s��o��o-�5�{e��.Q]jKV�uȞU�c�4�٭ۮ���EU@�B�JZ��d5�l�@���T�^��V���{]��lKD&,�!��>ﴪ5���6���f!��s!�@����X�Z��3����0�!�:ى�����Ǥ��0�M4ʣð:�'��H!k�n�!�w,��?Pp/�=,?����G����ư��w@;(��QǑ1��Js�c�Fk�E�`��d2NU���b�)���R���m3�p��d��Nh�7e��@GO��L�`hv
�W�ڄƲ�hI\��g{�5�M�k�x���'|6qL|�)K�z��MʰY�y�=����5j^�/�.�9;�����w������7�/ώN���B�/�={��?}������(.U������;x�����+J�=x���#;⫻WR�>�[�s����W�����&�����<��g��g��֢{���f��o�G�6}�P�jf4��!b��&d�-�(H*���-6�ݪ�j�ү�!}^K*�mtP\�wd����q��q���S��\�x;���2��*�ϙ�7D�\l�Ɔ`J*���� 0���b�-~�7M�����M���H� L��6��&*�ȚmOD,D�ɦ�	�2��p�!e�2،2"P�H ���ZeD�E�������p�`8|�)H�2[���4_�@��j�r�T�G`��ZI1E��'On�C��6�V��(��F��d����j������S.kUF�Ԉ;�ɥ!��I��A�P6��\I8�Uem���(8/+=5C^.��&�r=��N�84
Q��fH䆮�o�a^\~AA�wA�h�r��V�榦ؤ���5w�B4j=[v���[�!B!z6��`k�5��&#5�,/~j����J(�����;
��ᛸř�,�����*R������?��o��\�������G�[�ۿu�=g���?/==<���ؿ��8��~ħ���>��R�3�	���U����'�z�t��1=�9��?:�A���Ci׏j�~� ���lZ�F��\o�~e}�۶��_�|�+�&�+Ҟl.��Ub�-����'� �{�M8��>�Z%ŰCZO^�Z��ӶDc K��1Z�h�B�Ϥ�Z���1�v�lmZz ���GKG���S��C���F.ܼ�2 z�B����i�&�	��W��Ŷ��R�X�8�"�J�b�Kb痺�@��m/љt�z�"m���BCS#H��!�~��,Qފ�%{"S�ʷI��y\� w8�%���O-}�R�qځ�l�l���ҙ�@}���2,���\p`^G�"�T�Adl��S��ʈ�Uyz��->�M��}�$�U�C�@�gȫ�<�����-#�,�)��P����(��GcX8oHFQ��ټ�bktd��fQ��!�R�����ց(
�P�����<�.Sm�ia��#�&\�`�4�j�Ƈ���%�ݼR(J������ց�(�xFsbj��$^�c� �2*۰B"Pg��@�&JI������d㰓�m�	6��-D)W�%Հ�IQ�2�$yW��f)*fE����교�z4󅧙Q�&����.��D�����ix'i!�V��������E%���B���M�_�q \��z�����G?�l!�T/��=F�*�2�G>��En�����a�N͆4�.�^aq�
2v
��<}���z%Y�4�&����Zs��ȫ�(cC���p�X�.��!B��Jज़�C�\�AV�����M��� +PK�PT
q����Dƌ_X�8@�ː�,>�u��o�*G���SO4U���Y�k�談T�뫪^ȔMVaB1��� ͽb�-�UVj�-���dSH����B��x`�p ~C�V�rU ���7l�-��N�Lir!S�0ȄpiE�R�>N��jf�r��J"W'{fB'D��/��"�`�`�j�tn�0�W:&UF�F�g�\B|�.��*�Φ�V��	)��P��bpeSf��˻b}���G�o���A�o"�֊��Yw�\�t�ї�3��3��<���.��]�k�6��m7!�P��և{��HWmx=CV*�(}�������|������尕�����������_�\�Z��Ύ}��|����'W�����������ۓ�_�X?�r��v}��0�z�\��\���&����b)}n�ސj;_Y|��
vc���ߞ����Z���//��6wG��fo�=<�����_!{��s���G���ܓq;a�[�j������yٚ��vxK��������N�%2���7G?�ޱ�����Wh|)��o��Bk�[mf�����V�B�഼�2���R�~�î�]�];�QjCF�D�1�f�M|\٘��z.���3��k�^P2Z.�l�-n�g�z׶َ|�B����5k���qv��]dvA�*�?�8�1v�viى�}��Sm;����4�EF䛂�!���폑q�]�=٣M'o������'�D��׈ш�E��4�C�i��}w�YZs9גj#����DN��y 8_^�)�_�l'�ޘ0ѐyъ*f^:ڔQ�z�f!V���4]yΞ2KjR���14����K8]�V���o�x�%�ԑǐz��uתǣ"�^�Ζ	. B�hi��@��A�5H��q
��N?R�� �\�>m+ಯ���Aާ/n/�n�O^z����ѩ7��ӻ�ޛ�>���~��;+�����S֗/�z�կ?��_��sO���w~������o��y��_�8�=yus��<��Ϗ����w����q�W����ً���S��Mj;X�',c�Ì�[oFM6o���q�����C��M�F����]��F\z:�41�
p*��1����3;�-��'#�[�GfC�� �����Qc7}�tz�&\Is��K�W M���f�d�`d�1MAH�3��]�ps�SkA���M
��˰p�dp�eT��W
6C/0����3�4pҟ
#W@�Ƚ�
�V)@�=���p�5!\)3R0t.�(k��Ey�X]��7�zM6&���)Ds!�M�F�� �*I�2N��,�>5M�:����1T�@��DA� l:ĉ��TFƪlk����|!3�08�C�e(J"���3r�!�j�Vv8��1�Z �����]��y��4�){�PM^|�_T���7�^leK�O(2e�"�6X4CF��V���~ք���Gf�QK*W�gɠɞ���)�)�2
��E��)���7�Y"'.Y����oр��g�{�{w�Z0�'�������'O�~�#�W��NN�����;o������O���?����'�~��sh������#�z����>���uv��G�zk��ǿ����kg�����q��7�(�����������W7����p֭Mo�҈�=8��"~0�(�97YvͰ֞1��&5��\��-�@���0Ak���1d3:�-2Z�	G�R�����w��/��ٰpHC�14^-a]�p}RU[RH�tRf[�� z��3C��o��4�>�!X��nX�1�۟-c���LAx+�+^�H���t4��TjSH$>��f�����"8��%А~��:9p��ʕZ)rU>C�-ϰ�D1�M*��d��`���ր�URGo�߸8�4���Fc��JQR���j�M�Y1`y;�����R�0*,�Ъ|r�p��[���J��W^82Fj����ȼ	���d��.�aġlX�U�����K_T�i�qR` �*5r:�ǅV�M-��	��csQk:t��ňV1z�]ee {���T^|=0&��"��@��@mJbs����L��ak�VҊ�i:�1) Q32Pc/W
lxe��n��UUIMj:C|vxC8P�����p�A(�6,�-�׫QTx���"s�ŔQ�5Y�+K�EaR@ح�S�I'�&�&A �D8PT�~re�#T�^H�!8��2r��%V_R�&��"��Bv�%�C����إ�k�Ų�����6ox��#׬��Ԫ�]�p���[|%�R$�j�6�}'<|�]����L��X0"i��]�d`"c7/C8�����t��W3f|�f*�dqR3
����R�1�ȦP1�!��M,>M��*M�����Ҁh�F-)�B|6�dDUO�q���r�YGOm7���n͆
n��c�K�<�z�z|�-{�b7Gl��i������oH��(�f�������o�a�N�v.PÉ"ˮB}�%B��+�B���|���E.W|��x¥�Av"�Ѥ�L�g""r����m�y'�YnAk�����=�»H�~���ŧ`
��D� "a7S�.J��[8Z��D5k��>5!���r�#mWH*�Y�,�߳�;��Hw|t�ǫ�}�4/�����?�5�m<��ceݺ[��Ѯ;g�[ϟ��+���n��ݾ�yp,n	.��W.�\^�]�����[�~��ٹ?���翾�|�TOu=��{����e�%�����ܾ}�~�J�o����/��"�����ዛ��Ϯ<~�3����z}���.� g �"�������ٳ[�6���>U����n���n��owP�ȋ��~)�]L?B���������kҏ|�t�̧�=}��;��둳�n���/ظ	��җY�/:)f��Z��u:)�12q�c�dwe��/!Ee�r���=��[D�DO���IG^4�p�����mi(0ML�� �*Qy�Z`�>o��!��0w�#�������k�]�T�0�]/{��3|��c��ɵ�(��.E��v��-�]N���=����    IDAT1���a2J�k����F�І9F���'p@[ח5.��P��+�p����P��qL{ް�z�@�"�^e�˞C���ӡ���(�)h8�R5��#�� �E�'��LG�n?j�;?Tg��3VR`%ѩ�-��u��N�C R1
k5�l5PH9[o�,N�nq$ը!���a�8l��Qxdh�@�+CS�!����c�4	jМʜ��پn�'�\�u�ׅPM^��7��T�l>*$�d�tB��b)�p��A�rI��n�i
��qU�D5s4���#�@H$��(���;8�@�{�?���� �v��������ɣw�p�yJ��Ve�����O?����<���|筷{�K��'�}�/.����?e��x��^y0���{��wON�/���7��s���O�.��������b*W�oRن�+�Ł# ��@ؖ=�KC� ����"�
O�M�W_A�=���f��3�p�^�]�Tn��4/u��t���d�v��[�*ÿ�
�i�,��S%44����3��6_Xyf���ǁ�Kc�Գq�\Ie!	«ʤ؅��2��	�:;���գ���f*�W.xK�q6o5�ze�-��khVIj!l��!��P0�]1
�#�\�WX��^��#�l��R�z Ŭ*�51���O�Ӯ@��քȂ�&�����4S�����EJ��R�P'/�dy�_
�	��b�d�O"5C��QrQ�,)����I� � &\3#85�NY���T0��X�*,/fu��Ȏ��E�>2ċ�>�>��3L����wGЋW�V�m��^�m%5
�ؼ^��wħ9E"TOou6�"�-��M�/�a+9\c��7�Y�hB�5��"ėNYk�U�D�5wd \���u������-y��:�^���/.�:��&�����������޷�}|������_}�ܧ�ǏN܍�E�ۓ�Gg��.�=���?��އ����_���~�����_���~�٣ ���4h;�0y�/CO���nk�D�Tv����=��/^��SSv�4��7��f�`Y� ���1���;���V���5���"���m	7��؉S���ՆV:}B�0h�y�`�h�	�,�fsaÅ@�`��]<e!q�c���@��Ѱى])�� Qޭ�8~����8ü�Hޙ 2�K�i�3F��!$���!z��r���	�(�Dh�e�
2�Nm��"M^�N.��:"�*��8�"3fH�><��I���.i
Bh���Z���(�9�@�2R��+�m.�3��B��v�����U(|�8\l�x`��²i^B�DC�W^!��q�#���3�҉�k��N^}!�
.����ed"d'�&���n!&��\y��d�#@�{���)
atZ�tx#l_�ń����F*[�֧Ԙh.�(^�p��f�B�fͨ!3��B�;"�l�
��jH'>B�b@���әt����B0���ΕTQ�M1E�\ͥ�h���
�,:z4��8E5l������j؝K��"C4�nj_I����)����[N��ÆD���H�v����*���L:dvZFjl-�y�'h1ͱp���3�xLC���Z�٫���23� �R^�C����F_���l!!���{QT@%�%�r���� �	2���"P��Y!W5'��w�� ��W|R85�n��P�>ox��Ҝ�2���EиR���N3�i�,��2�Ga���"���e�ޮ(/\���^�����8��q����Q�a�M<�E�th���s�A�Q�p��&��[FL�pޖk��t"l��W�����Ȥ��V�-�	�Soh��0��4+5q
Eq�ut��+2�Ʌ�A"ď ���-��C 5�����U5yG�@ä��0���cBF�ݤ�ٹ��NS�ϼ>����?��5o���
�f�P,N�5�K_H�L.���r��
�k�q��K6e�/Y�z:hp`�d4����]�[�3�B�c��by��Nj��\�-�7.[����.�)�cd����]�L�g�G�Olo�A�J�Q]�˪��6A��|�uO�����~!e���_輹�����OϞ�x��m{����Ww�N}���`۹����p#����长�=<^Ļ��+�s����{Tt�H���Y����'c��)�������'��֖P��`LR�_�4S�v�J�~#����e�/.Ś�����W&r�����Ƀ��'�t^����n���n�}��I���J�+�n����2n5�g[g[Q�����І1AWY���j���1�txM`�)���W�l^�(◥(ʣ3�.8!�஍�;ܵ��2"Vf|��G$c��=��a��hߜf�p׈<��ZY_�_�p�n��U��0�C�H�jM�Q�o�4sM�d�pr���#O���{\
W�!��ZFd��&$]���A_�p#�5%���YX�ݨ��c5Y�r!�N���{��Ȉ�K����AF>���bj�S����&\"=N�	�rC3�K�HY��j�\4kѼUusN8e�y�g3��_R.�?�C�v�y�2��fhM3�R�3�V9Z�Y+���ɠI$�p�h�A6�g�����^^
��,�~�[�Jݻ*)���S�M�z�oj�q��������9��-P��'Ĥ�I� �hp}�T�as�tCU�ŋB��/��L�Di�h2ΐ׿X����}������u\���[��7�����cל�n�.��x����yq��/~���/��}������G��><=;?>wLn�����{���O�_�ݼ<������(�Y��^�C��;�0�f�a
�	�B�S����7_!lm\ҵ�vs���2�϶V���B��i�\hB��ֿ� �@���.�eӻ#�]�����B�<������J�tz��6�@�l>=>�v0)ӄ���Bʮ/���q 1k�@ʚ
���E`3������KY�z:ց+��h��!��
FV�,B�tTh=w�����d���b�B$�H!��^�q I@���0���8Xp6>C"�2TH��٢��Q�"����%5�g3H�ى�ek�LP
��ٓ�2���F*2�d5�m�����Y8|z�R݊�(��Ł��g�Z�z�+^^�]>P���,��<4����&c��lm�y�	I�K��2�֫D/�ٙ�	�5\���e��x@�W6�N����y$j��c^�⢈�R�S��+z���է�|���E!�7;=�xL.�\��c�1� �UU������/
�[I+~�3�fݼ��{�E���z:f��c��Y�U�O�^c}<k������ͣs{z��Ͽ���/-݃��˗ONO=zuy}{~t�'��ֻ~዗7W�^>yu����?��[���������n���w8W�'~+�#}����C'�I�.����������.��'��;�~��gΣ��s�����r;�,��x�jjʹM��bZ^��]7kd�\-����{:�������D��敫�\�o�j�k"
��JU�6
l���=0$!K����!N`U��ƈ�O.ߐA'�X�#�Nj�Ԥ�b���5ʓeW�� �lyE�Է���)[��qWx�# D�b'bH_c ��΍��*���Ð��lȀ[vF!j&(�,z��dk�S��b�ђ�oXR�F?e��d!M9N�e7����MAlIM/
��tЇ��!C�T3D�w�r"���ZƦ�^;�z������4�[��� T�.���%��Q���F��1J7���J�w��aM��e�͋K=�@�0���2�U��~
 �'��~]yR�8C"�r�Q�h���WU:�jA��9�s��f}Y�8o��C�%(�(��ˎ_az=�W��BjpjqBv5�����2���p4E6��}�Lͤس��lF��UYx!z�b:֘�SF3w�Ъp8�p�]�L���#4�&�p�a��:Cr�oy�Y"�V?�+Z:�c�?S�rslMR��9e��8�!�S��'o�����-K;�`�B�d�'Ș���Z:ٻ�J�@46q8�&"*�B
���h"z�^��7�I���=���#��>��;���s�S8o6C:.-NŌZ�'���@�Plu��k:Ȓޚ(�-c��!�	d@�E�㷞��F�H��!7_��DC>Ð �ݺ1$��[�e�Ɔϫ�]K�����sc)�@m�٭X!�◥��l�ǟ"����DDD	�XH�6�3�04RB�5tb����g��,�,�i�ؽ`6>/eF����B���d��l�!B�#�#[��K�Cc$"�K�U��w������������N��&;cSZ�T��M�}l��s�VpՀܞ$�njb���<�1J/X.�\�3|P��aR�pH�^��6�a#��ʋ'����Z�L�Z
fmʾ�ݹG��d����������UKt��c�d�Μ��o._��ؖ�pƶY��g�����Iׯj��]zP��ܮ�����G.�<�����.�^����q�ʸz�l}"�����n��H{��Q��	�����W_ݭ�)��|�ң����<��6�T�:ո���9��qV�W��͕{���wW�xݶ]�U���ۛ�u��e<��`�&�SONOn]�[�����WgW�~����oi�����[?���5�h�Mzs����W�Y�k+�-��J=[c[#N����؊��{p}U��`���>^��g�z! w��攝�I���n%���!��	�Fd:����
3�Õ��<">!�4�QHmz4�ÉB�£�p.w��fm	�&O>�7D\i�۱+�fPf�lI�
�w���T[��,<)��"
/ﮫ�1�L\�
�@�f�gˢᴑF��W�tݵ\�)0l]�0�jFvD���N��t5ҵ���:8�C_���NѤ��l���&� �����6�Dp �2�4/�� �$�%��I�jK�a����æ����	ѳ������0��	��f���ؤ��]����(T0�M���)�T_m���VT�d��*�6d
vp�yk��g�)\�f�񊥃sleT�>~�W.�Q�Nbnx����O>��N�ƣ���p�����d� ��v6�O#�GM��t�d� V���P}��߲�%Zu䒷@����>�x=��O^��������o����[c�wz�;LgG�{{��^���/�x���;�}rv����/^>{�ۗ���_]?����v�}����}��_��O�>������'Ϟ�����{���������7�����gvMMIj�U�{ܿxB��G eX�u@fs9�h�C�A���`X�hz.x�*ؐ�W���)�!^6���ﲾ<N􆮧�'���`�x'���~f��Rn��>���2����
�]c�)h^���h��z�v���
é�ȓXk����
��))[�hj�hM��aAIN��4^4�14�\�)4e�4�p�9����z�O�������F!��m%q#5d�������6⎔�p�^�^.�p���:G�Pߔ�GV��2J��xk�8���X��uZ[�SF�@N��¤4���+�\ei�����%BƩ :P�,�D��B��z-$B!
nS��R�,ᆘ^S�.q}6�p^���q7��aHdez��T��r.e��I�>�;ym "R#�Q�����%դ���z�9���fԒb@�eH�6 N�pMU�d᭧�RE��gZS��¦V&h(�M�Y8.�ւ8˽����/����=�˫W>��r��Z^<y���s/�W�gy�������Ň��/�?:�}�d-��/�;x��ۧg��}��~��O�����y�ww��)�>�g>�9�>�\_����({���xI�͟����/�c;��yN��yR�޿�2���P�ּ�O�>@��� #rKm}:�h����=���[7����a�EO-�]����#2�;�\�+/|j`�ʛ��D�8k�DA��O�i��p�h�#p5q�JT.xGA.�8�\l����W?j�]Z�:�
�iXv�R'�5���:y[����ڔ-
XπW���%����Z�x�FdR0J$���~v �ae��v#N�楯Vf�n8����*�&�����<0<&M|6�ԀPv�ٌ8� �7}� 4�12�Y��H�zC���Hqip`F�	�� o�5Q�\\��'�ajE�d�.0>�����#\�V�x�����hM0��(&A+o��m���R�z�
�bĲS&�HDI�z-����g$X�]��չ��w!ôIAܮ���q��,6\�l̲C��X�DRC�����02f4H�!l��~I��Ȁ�-S#dkM������oSȕ�����0q����jP�S=l�p�Ɗ�s,�����pW��˨/J8�a}2����A��A�փ���P��auꑳ�K!�>A"v��(�eW[�A.��K!*;o�#�jE�#��i���:��%9"@�B�5����J�wpލ�^�����//!/�B��A�D��+F��_J8���$�"�i(B5�5L8�����K���\Z44Q8�FF�[lM�y�Ӑ�<�-��"�D,MF��sE�%�b�ad�w�P
CFh���A4���^b�ƕ>������[O���ST��S"��7��!���J|�\�7�5C|��.����씣��W|�^��"C���d�.�7#|�o�$"[l���|��f��A�I?Z�h�24�e�N�}��G�2p4R�B+�����8����V����kY�)[v�ENj�����W��ah���8�
`+�gv�JJ�%-��=D�&�ƅ_��lCd)�+�yU���A�R�t0�kR����\��o���1\A���������ŗ7�-����t���+�����s�ں�璌/D�t��ԥWoaR^�����Ƚ뛋�g�
:<�����s�]����[׌�ݱ���w�%~��������4��\Y����Evv��٬�G_�tW��f���j�H��]R�G��[���.�m�m3��. �%::xu���n������{'���n����5���냫��/�}��=R�q��\�[���j����zq�q���D�z�y����J9�F��#�Md�U���ہ���4��kB�OeP�����ʰ%�q�w-�@4.�;\�eSۢ�&dP�V�4���w���&6��˛��Z�X�W{X�TQ�8�&��0C��nGd�q��bkB�1\�p��Y%�hZ7+�Y��_%tx�fdW�Z4/��B�󮭾�B!5�Ls\��&�&Vc
�C!;��l���&P8|jfS�շU�ԳmB�%�()�f*Ď�駟���o�y����Y:������+��qR� p��) ��eWj�W!Ϊc[(}!��&({w����7�EV�^U�W�J4�B�Z��TŅ\ylxԣ)�QR���&�Far!�
����b��w7d��[.!��,�R ���EG�.
"���;��yqz8D+�a�9��ly56�Ld�3�U����+`�t��Gpų��#[��\���Dʣ�&�?��?�ot��	x���us/�� ��f��V�!��\�
�����ky���4��4����+O�v��[�y��ӏ���w�~��[�><9:}������|����~��ã�?;9?{�Ջ�_\}���k�}�*�����|�}9��O�_~�����/B�i��O����˚�џ����W��BS�!ႛ>PmZ�F\L�i�E��A���a�	�f(o
�y�B^x=�Wkyr����&�w6qC�*�������J��&�ucX.����k�fjH��R"��*�W[�m�^��Wf+Y1�@MTdH�-�Dd�]��+7�jh�pF��e� 4��"A�S�w_"32q�_�)� k�ȼZ�(�zT.��罶�[j���j�)D���S�!�T���Z1SU�T�����e���С?�!Ze#O`����LA��x["A:ٲhQz+c�`��*C�X�F�C���S�Y^!�L���Bx��!���J����#3d���    IDATZLQ8��Է���:ReQ�5ᴋ4�7�6����[:^����x-���obk[�{k�%I�"t���:B���c4��\�05C��P�2V��F6�IG8��b(J/�(��:@v�jSI���фh7G��*��9"3�y����k}xk����m�tv���[#���v~�ß6����D�h��м:x����w����'7Ϟ������_�\������N�o���?����'{w'��i_z���5���m)V[O�Y/�J�
�1������5�=�S//d���$�5Sl
+vk�k���'I��i��	��J�z�y�y�%wO;Le� X%!p6�l�y�t�l.Qf2��j!��-d����=����8�p6#d�G!���
S{U��+!��6��"o�?�[�j֘�Q#��0�E�<�H|e ��T��������)�`��o"1�f�wDf�8b+L�|q4��:.`ޔ���\��Bb�W
vQz���xC�ƅن�6ddc�ڵ+^`F�,)�\��>��W6�Wa�R4 Zyӏ�L��,(�_�ȩavD�gK!
G+*[��MI�eh��V�]��Y%S6d�b�M�ՆH2���	����2�f8:�DR3�a��l��v{��7k��N.D�A�����K'y���f�k1�y����Y�V	ΫQ�&v�̀��7��Ψ�ʢ�(�O��j�j(d7�D��Z��a
�F0�r�(PTGa�� �(
%�d��a8�9
�cJ��;j�S��5xM�J
̥ߝ,M��TR��#7�h����7�0���;)Dl�z�VI8\��ry�R@�������b��`������$���h��"j��7T�Tn8:�p���VO@�+���%l����k��X�΅,�Ԝ��N���$�`�Cҩl̲4��!$�lI'u��S�o��22d��-�A��"W'5FFI���P~��f)�٣i��p�DHM,��hl��P/0.�>��TOI�b'(D�SX|Gd7{���T`uZ
H}5�c6;��^x��4c��]��@=��7MgW���4T	��c�E��������g.�ٓwԈ��B�Ǧ�Q�³1	B��z̐-hm��t��@���1x�P�d����LG�a^!��D�C����?���O\���3�Z�˕,㍂�M�mq� K�`=ܿ���hI�B��(c"X�jSp�F����L-�bvt���Ԉ�wF��)9>Y�V D����V�-����\A���5c7�D�,V��<X���պ�PD�IćPN}�SA7nN����{�k���I�4:=>:�3�΋n��9K���Z�����c_�\s�;�~��Sq�x���\t���$���g1oI�ݝ�_�ǹ��>׳��m��o<ʲ���y�����[��kݽu4|u��gA��_��W�9��_�4�<��p������u撬_�|u��C78�./�|����������y���]^����ʨu\?\s���e�;2�-�˵e�����{k�������=ra�uX)k���l8��O��o	��j\�q%�׵\�	u	�0AE"7Գ@��5 e=\C0��@W$��؟8�&����H�P���I�-.p�o��Q
xk^o����e��A�%V����~�� p[\'�P�G?���,�,P���`��Jg��(�"����~v�bf(5�U>��D�֊�W"d:![�n�kmM|*��'NDo���X��p|�ù4C"�*� �,.+#��u�p��K�ld�\�T*��⦛D�q�~):@��a��zl��s���{-�:Q��isK�d�6�mĆ��&�ys�\0`�B;�-H�E.�GْE��:t��C~��w��Rc�xꩧj���=��lS&�\E���/�a�hj�Yr}
��ò��#��4���)ߪ�D�尘�����Fj�24���H�� G��-Q�c8�L��]�G�F��c�d�5���
�DH�i�$XR���||QLQSKJck�=����i���V~��A�Xod�LuuK�"��Q��)��wy� BL�d�k�&H�1uM��(إw�}׎��3	:�<v�C��L�c���!�GQҢj;��@�3��U7|d���.r���C%nZonSrO���G������<9?~��>���|���F��_��������_<����WY�Ȥ|���o�����7�����={�ݏ>��ū������٧����=ݬ%�5�l_�Y5��[�΅�!|��ҡ�3�9ko��@ ?P�C�r��6�._
?'�t	m�
�ߢ����眨��H:��Â�*���_��_��:�VR:�H9����бc|:���(�#��������Y"z�I���"�� �b��q�"�Ŕ��,��2�1SјS�&������\!x:�%����Y��c�Z8nyJ����<_��N�h]ij̏a�TV��F�ZuEhd�CM����d��(d��
��D�+��A�1BR�4O�X�6�Ta���H	Y���AҌĖ�͇ �Xn�����&J���AF�� ��aS�9cueins�(A������!ӿ�΍n�D��	RH��5�@��v���
1�~m� Q��G�I��կ����R��8|&b��p�@>����2�\W�Mz%��̑"Ĥ���4-M!��cB\>�')g~�p�����-�9�m���{��t��{/�h{	wrt��O�_]�\<}rx�g�N��x��׾�ַ��N��������Ӄ���ͯ�����ཋ��/~��{?��+�������7O��ߓ�49>?��M7��7H�k,�����������������9���7��ClQ�4v\�݊� �6��j'�r�+��̎&�	$��$��9�	�ܖ" #t��o��� 1K���ɉ�Z��&�B�qƙZI1S�k�A�R�}8�J�h�)D6���~z;١�ߺ�9�L"ɮ>~gdƉfL!����Y����΄V�Hg8|YpH��th�s��"a���M���b�?Y%�ش��iI��B��¯JFHg��=��iM.�ئ�јĚ�4�)E�E[���\ME��OQ��A�1�(T�/Z��
Y�1�B!B�)�4�v�k�R�#���+� �&�'�l)��>�xU�<�C����I�,1媧O��}�Vߛ���4&k����m���d9���f�3��9�|��I_5��و&
������@{eN3�Ud�rjL��) @�R�`�# �Mo�V�S��Ȗ����k�N�W�D##Xq�@���кjXTa%?6���Կ)q�ZB��h��l�p2�	���RL�(���!!��G�B��S)dG�Z���IqL+ȁ]h���\Nj:��_J=�ƍ8�K���;��n)������Sf�GY
&#�`-G��B&U3�6�u��$���Qh:�98M�P`�%�)Lo��CJI����l��8Ԍ���V��Q�P��ں����JE���*�&��QT�*N'|'@���1!>�Dc��{�0���%^Eg�����ÔˈwPR+ߔ55�PF�Q鍜89@
��H"9� ��~��O= �p�!ܴf�d����z����r�р,߈���VO�,��Ԅh.�퐙�6 ���zF� �h�)a�GHjtL��W�I1�B|�,dD��1É���7�c�B���8�J�&��B*rR�,�I�	I�kؿ��>{�̋>�M��_�~�s(����SrM�,G�R�m�B�l'�L�t�;�r~�]+y�AI�UH��ȇt?o4�L����W�ވZ �_<R�������X�{�Ӗ뻀֊���=ռ����G�����=��(���%A���'��B�[;�]�=\W�#-��Zɑ/0ھ��C�^z���������t.�:=\��gaE�;'�(�^��<�#||z��'篟��>�E���/B��Պ�����|��2��H9��W�
�\#��۽�9����u��z�J}������ڴ��>��	%����|su{}���nϟ��͵
�1��[S+=�����ݕS�����T�/�-��u���V��E�õO���ݙ�N���m��ﮝ-kc�_�u����ȱ�w!�z#M�v7�n�7=�.|�᭷��y��8.�~ .�ZM�UQ�!�%�YQS�N3!UL'���La+�p��'nLP��f�L��@酀Ȥ��T(Y��`9��b?��"�������qD�L���n�������ʁhC־�r�R�c�@�B�	�F���(�gS��V��bh���lJǡ�V���VK:C�%��9���H� �2�FkW¾��5�-u��1�V��x�.��9#�K�ᘒ�)��S�E���!6G�)`�/���>Kp�;1�8����F�r�E����H�M J�[#���0�@��S[��')���q����.A	��o����˖�~,M
��
��|ki� [��]9S�8p�Ʌ����mi�dQ=��Ӭx��42�m*d�,�\A�BU��Q�����e�Jsm�M�܃s'X+r�Yi{�.�ʴ#	5	B-Ք�n2���b:H��CY��b,�x~�&k��m�|Y�L�2�%m���B���_>;���o����3�7�o~���}~�Iw��p������/��g�҂[_���3����/]X����}#����eW	�����[����(-i��D��i9-aȉ�V��n���5�R���b���W��qT�&"1�-�?#S6��Tڔ��p�:�0���޽�����~�}9�]��?�Sg´d���^Kkd�Jp h���l�����3
n�#�%�i!���Q(Ydf��!�D�8����'<ͪؖI�+4j�� �ꓦQ�5���mr�G��D[�D��1��wr�����;�F�qM
a�TEcƌ�բ�!�BD�q0[��9#��
B�jՌB�SZ�$��Qi��8"@d���T���Jߔ��g����1N�Y��_!@eun7 -�f���K1��(��'U���H�;�#���t8�M�O/��
i�c$ވ�񻩿t��@���^[oo[�~,S�s�ٟ���>�)��X:������}����Ǎ�e�G�*t��$[4q�d�.jj�U�<mXQ��)Qz�������6z�+
q�'�%K��h
a�����W�/�U{��ߌ�Z�����ۓ��מ��'��姟��_?9}��������^�����K/�8�����W�>�?^���/����<o�7S��N�K�ӳ��e)�/u[�σ:�ۯ}����b��d��cD6u7vuo�6�᥈(�K���aN�NK�N<�
�����~�c��Bۄ�)���
W����є�sJ)$�t�U���,˔��*@t%�r$��+��)J����*T:���_��%�u0��6>$r���QF��ڈ<���%�¯��>YR��6�f ��Q�
E�����*m���
m�W-ߴ�+e:L!f�~c��(�V��Җ��2�'\�*�Nې���i	���[i#�!G RP�M�Pd �t7���Ho��(�J
�S��O9�IǙ�F��L>���RK�Qbь����0%�8�!�Nxc�QBM�t%��h]�M��AK�Hy�$�'��CSRΊv�_()>G��ƜI��Q�#���-�ag4�	Ue���)���f�9�Ҍ��K��qS]4��2���jIH?F�����_T�ё1M�D����8��5i���pN&JJT�Ь�iHE�R�s&�T	cG���@�n,
'U?�����_���i''��a�h,߈)Z��
�����LD�P颦CP7��O9Gn@\㝇#����(ԏ鴄���Wq��MG����4�����E�(�L�Bp`����Y;��c|���
�8Y��9jÙ�CK����G��P���9٘�i��ꐮ}�.g|>��hSc����CG!#�\d�6�D~R�MA.�)m֨�
��@;☬**���O�Dx�dŜ�!�$ȯRE��gued�HW��'q��?�D3�h�t�'�|���x�AnK�eq�j�)�ʹ!��%:!�1�N�'�	��D���t��h�sLhJ�8dsV����q�4��1BL�B�eq����#�5`�a|�FS�1N�c�J�{��մ�~������7E��l�Zg�f��-�sL���%w�#Lc��B��U!Suۇ��S݋,�n��o�Nj�2ҡ�ɦ��q:�q ^��Gz�fL���/ǚ}�*�U��ɠ�@���'6���]A��>e��`��6�߳������ds<*�aKb��s�V׳��ݡw��6NQw��퓠��g��}����S9]��o�X��ĕ��_�3.��;�޾����]�xu������^����c���g>�y�rw��,m��Vck����gu�nGA;���>�k�Q�	_���wW����ړMf�y��������cX�����Ͷ�����������7/w'�����~wp|�����~u}�<p����2qݨ�z��hg�����h��/=2���:YF�ő҉���cz�K�[��@�^�wk�r�x�#�tc�t�� t��L�)� ��N"�D?&CC��t���|!`�FYF��a��ճ���L�tOPK�����R�^U�~0mq+B�7�"��N�NE��E�x
e��k��FY���i�ϡٍh����� �����5U��l����!1��$%'�r8����j��t�Vg��ړ�B4&W	fߤ�RU�)��b�D��'�#a������<�� ����;Wr�TX�JPsv�p���j��td�&��@����A������5/D�O�\Rx]���R &�^��#!1�e���~�m�C*!�{w>Q���s�Q����{�[�ʡq<�tEqtbi����5�(�m~Mj��(�DQ��T;ОK�U�t>���8��@8�@��\L��-�Z*���GU�4�72�jt�>��7������ʙAp���������r�;��*'��6�R����T���'�q�߶>�)K�_��##��Q���i�gw���ǧ~B=�◟|��������s�ׯ���uy�������ݥ��y'g���?~�D���:x�k�_��Bg>��34>sx�'���l�+�گO>��}�c��/ץhE:Q���R��u�d�ȩg#���T.�	%�~����˵�d
os��<}~����������i�qi��э��"H�����������!��9IT�q&(�lk�:=����|Nj���.�F�.��^�|�Z��R͈��8�ө��QƔ���ь���Cp��1}��=A���&���8�	_T"'���r�@��Z>�B|[�¡殺�����h:��G���E&��%.ZW�i֛1Qd:�������I�ί�U[��9F�j��0��6�m9�7�2$0��)�օ	�C��
�31)�����=����5�#d�l��z�'R�U�YR�S݊�ҍu(����V
�$CF nT�X���U;��I�
a�eR���뷅SSK�{�_s��	��n%j�QT�4��Ԍ�%e�8�y����*�4 ��*��T��v�djDN2u�"��4��;�D;� �}����O�מ~�!�x�m�����~��ίo/�|G�����o?���7>V�����/Ϟ���~���<�>���������y��>�yutp������������>n_�sp|���y�y�L�ˀVe��Z�=�4�� [�5�o��h�tbD��Q]
YYԈHlǜ<���b�CAz
��Y�P��IQ��4��P4�@~�
/7fcU��4�OGhE�T��F�R�u�L4!�*50ecR8BF������U!�ܩ����J75��f��9j�pcj�Rq �R)5^�uE�X*�a�|��BM�JO_T	��ttp��"���b���;���%$�$�s+"��EI�h~Q�~�Qb���h��i���M���@>'q��8�!4ѩ�q��L�g�>�z�T�I�,����	꧍�+js�#2����5�	Gn���/��&�M9�X�    IDATr+���tD�2�͏��3)����)�G�C8s�����8��L���:�$UEQLk���#w�������C���/K�*�V�Th�d`��P:���@+��V��%� I��	��؈��O<�f�W�#�f$r���F��BӤ���Z�*dL�Qb��9��2���,�
��sX�m�Ģ� �*���N:2n��)8RF0NN����z�Ý��2'�C���O:F���Ʃt0f�˭��'�m�h�QN��oK�&X�@�X�i���sL��fB��ۜR�R�PR_���:ibDl>�A��ߊ���J�1V���-�!�T"<p�L�GN6��\��ЊBF!�@dƏ�):�p��JbH!�vF�h�I�VȔæ��!UV|�Vg,%�8mį"\Õ@Ќ���4M�-
M�UG O'��hmHa8�_4��g%�+jC�X'&dD������J˚(�_-���LT'��J�؍�p9���X�8El��VZ(fP`��碦)�3k��I����}�^�H�����C-!$%d*K�U�T�y�.T����
_b�Q�*u[�����d� ��OS����Ǜ�4�9eY���=��lD�*���yxy�[�N<S\y�n'?d���խ7q|Vҹ������И~��d�C�>o	��C�>|������uA��'��D��2G���w3w����y��|���tO5}�t}1�����z��٨o�%{|�>�\���~}Q�ϔ�Ch�{p׍�GS�W��&����m�S�)履z�+�r}~��_��u��>拐���.��뛃�������S9ke�.���������D�������5�f^���^@��_)�N�z?]_k��}~m�vu�L��f�)��6i;��5=����w�@4��Z�j~;�pgH��)5S��弓��ݻ��g�rx攈����߹ġɼ+҇��{���%:��	W��Kc��5��@�������m�uEG�R�}�]�vٔq2)�Ѻ����ũ
�; qQ�����3Yt03 MKȼ��{�@0'	)��j�#���Ϩ�hƲ�WT��|ǔEn:+2�d�R
!g@����#C��qbJL�~��h!"��р#U�hB@#��zh��u˱'6���`X:�7��'��q�KG��,B�&f*
�-M��q���nc��Q]-�٫��6�\�h�$V�o�|�}0kq�t;���U����.Eᦪ�'��N|��U��~��w�y��&�[Kn��/����'�(Y:��d�S~�,<ȑ�pD)�XSN=�X ��Bk-��N�Hm��QcD�mS���#���+7k��d�3Ӷ�FľA(���A'���{��]����ܘi�����ZT�oIDհ���GĲE�)�l��v�ĩ�Qg�	G��B��1������?��������{���0�������_���r=�{�6K�/���%Bj������ao"�+^����������Z��!��?ІGw�~����UWj1!m�.�m�W��a��8F4�t4m4����Y8��+������RH|Q�Ʀ!�Lu�9��b?�z�[�)�ӟ���C��pb���_�����ߺ�A����	�X�O�i@u]9�8p��<��gYp:J�$b�i�hB���ii"�46���e8|��7R��RB��(4�N
�+���)2���"��������@�G��k�(�H��i�|�@���7m3uy��"�Q�ȷ�ri�5���A�98�L�ZFd�hG����*���#J$�}&�Ñ)��h!����$[��V&�>Pb=�\:$�$e�~�d1 D�z���8v������mE��B]q��KC�n	��Et!@����]��C��T�ݓ˟��碕���t3���gG���Bpׯ�|��w��7}J��ê[`�9�N �i���Hg�Cb������g�,G4�q_�&}�FYQ ����Qh*�'�SǪ�vbC8~���A�oB8^۟�����o��
�����ۛ���}�oq�]��?�O���������+/瞜߿:����7�����«��W/��������<��l�\�����0q���������P{탠믈���ϯ{�y�*��k�,��i�V�CԤ��phB���^���NKQ+-�H��S�6D��%q8e8gͪ�,�v^"5)�}�H��V���"H��9	�H�X+�2P49�s�9,����ZZ��r�_Q��QƇ����gZc��ɑ̤<����\���mo9#�	5B��	� ��et��%M
qx"	n��0Y|�Y�D�1U$tYU�2Db�eE+�DR������	?�rS2x��Ԇ�,Տ�B�f�8U��p��!R��JA(]4ߴUp�۔/75Z���c6"̞T�1Z`飓80��bZ5$5�I���-ZV��d��Г�$.wRL	��EGA�j-SVH��κ���?�;�x��7e�D�G3�*��� �-��B�(���v�Y�h�tx�+y�$�˯4Ǿi�-J�dZ
�R����7/��+����h�p�؏V窸P�>�ND�B�<����#��-��N��QA�tL���p��;�RH�/��H��	�#(ͦ��h��YȘH���2!�\{��/����d1���Uc|
��K�G���)j�T�eB�����pc��5oZ����؏,�� e%[K|�F#�~�@�hٔNP��_	����DYB|�?H��BK�����R�(�N��%"w�Z"1���~J�*�
ȡ�99Yp�i��:�����oںD!	:V�c��!<>�,�ߺBLK4N�њ�U4)�@$�'����zH���ì7<#\z�­������P�T�A�ȇӬ�����J|�[d��v#5)�!�b*�	iLܘS(f�1���z�@�Z{e����iZz:B����Y�4��>K��d�����[2-%�:o�A��ħ�#2Y�S��d�%�Z-ũ
�7�w{���
ݠ��ř�мe�Jg�;�a�S�%��G��Vt7�4���1��B88V*�*���}�^UUBQ�~+W#M>����L#��J�D�xq�p��wk]���c�_Z�& C@��ݮn��px��&���K�@�v��ո��[�\{�;`}�����2}�l;f���ũ��G(]'����X�>y�Oe�t'A�����t�z>�{U��b�q�|����ޑ����*�=��7g'�;ռ�;>8�]_����n�n}����f��ds}?��ן�t��W�G��%�1'RΑ��6}s[�zt���x�z�rw�������f]ޟ��z}叀�v��>#zt�Īw�z��!�u��m��n�/��������H����(�:@|u����o���Y���7�'M)�v�;�I�W���	r�U�Z�舚J��G��ë{b�F�%���!x�������\:ޡbԜ~��?l�L�sS]y{_�ei	�o�4Eֹ�@Qo���c#q�����!&��dDtK�,�Pˑ+����g͈Ni��,�@#_K���w�|���tD�#`J4M�G+�GВ��"Z:D���!�pXʢ�v�,��D!&���d� �@Y���&2!x>G�(�8\"Ĕ�M(¤p���G�U��
ql��5@��XNoQ:Ӽc�|PNB�D��@JՑ9d���Di�>��y+���� ~�N3:p�B��p;��ф���"ep~�J�[�u]e	�i��]�އԃ�]n�>8�u�ag��d]M���ܴ��n���6�-��/*��s�U�&��i��Q�a�N�#
OV�T.M>�@8F�
�c� G�ˁ���%�Ur�fh�3
��t�˓`�")�!b?-��m&K�h��������J��TL�*L�@���D�@O���Yn4S�F)��\`�a����ʅ0E������ђ/`�9ӿ���q�����%FN�j1KЌ�ڨ�pg�k ���~�3#�M���ٳgn�~mB����4�	�7=�uC8ȭE���)�_�ۆ���"KA�t�tLcK����A��N�V���ݰv��N#�sENA'�[o��K,�!'����!)ʉ�:�j�~jO�US��V�N'�E�^��z��0��J�15"Kd��6�՘������t7C��b2�"��բ����`�+���$"��(���]Ml��$�dM��!�%��
a�X����Gp�LZ2�qD%Zq�a���r��8�||>�F�pVB�@NV3r9���P�EM�E�Y�K�yX�&��/�\W�x~�z,�zc�\������*F���roYU�з��Q����[�>�4)4��,��K�_J�DP�,��VX��,���CA]w<ם��^�r���@
������p��'ı�nznnJ��1gu|S%D�BL'��h���W�_bN�su[)!))���YC�:���܎WmTZT.�hg�jy� G���S��WV稙2���#��^%�na��.��Z ����_����{��;�~���_����ۻ��?�~�͛���^��~���o~��[�7���ӷ����֫�~��~�淾���Ջ���w�/��[K�9���t]����=�!X[�:�ȯUGS?F�e�6�D�E����Q?7�4�E��F��Ǚ҅�Cn��,�	II6ܨV>�*�H!k4E��\V:���K񳤖覓c��U#Ө���BƢ�ZR�Ä���@~�j	"�JW���Y�)'Q��X��m`= �(ꈐ�^KU7�.��l�<A!�cu(B��R�Hَ9�G05#�%��P
K�(D+�յW�}��M[W��=�D
duh���V��f�Z�SW�n�F�~L9ģU�,�49�}s�q��I6)#C(��a���W���1#pܵ0Ӝ��Ǭ���<U�S���$��DS�):N{+Z����Ѭ�������@�%2Q�)�<S"�����QK�NB����Q�ݠ �Ĝ�v�K5q!:8@jS�Cd�ގK�
1|YY�[H��ؘT�"�_Q`��8ʵi�攒�a&�͈R�y��b�n�^?�t���#��F٬~��pY�8)�7��dE#�K�
,Z�"�� �D !1KƱ��d[����Hq�Z��g5���T�H��CY�i�VŘ@V�3�[�(}>P:���$(��5�ə>!��.�8NW`�C�Հ��5`OLs�8��m,�@��)�*N	��
u9�N!YpSR������p�ET��Lǔ��D��0)�� r1���!X�A��($
��F!pV禣�A��&�3>��$�
��*-����Rj	
�V�D�3r2K�	��Ǭ�d������D�
��,�tR�(1q�ik�E�N=g�WK�b��*K8�i��+��J���D�L��8��ȗ,� ?N��B��q5���o*����r�rV�^���m��5I�e<h>&�1��_��hE�6���h��I0)d�l�
<?�T�1A�Z���RB-)�'ȧ���}�/��/�^�v��Qz�bJW�U� Dp�ו�B5��7��5�,�,�5-�Z�RXm@����dH5,
!kZ
Y�)���Iوo�8_���<��_�\O4�Q��>�9��/��;X���B�s��G�����T��m^�y{�Ӛ'�z9�<	��3n����t~��D�`ԳFO ���[���J]�7�zѲ�����r��K��������4t֛��������o��$tr��m�2�#�|��g��:���zζ��kZ�ZfW����B2���}J�G��ko}a������|��Zd�B��'>����ۃ��t��1s��^���Y�׬��yr� o�aQKX�A�;:+��]5Gj�o'�(��e�����}o�{WGT:�7"��5�5;�����3�wY-�w
kQ۪+�\]�g;I�뽋�)w9���H���G}�b�}��|%��aT�MdL:����j[����m%��8�*-��kt�Z M�������{��d�#��;>A|"����c���&]���%ݓ$OA��C�`�%B$�Z�er4��H׭o"�3��84�($<Ĩ�8h��ش�����o!e���p�AH�Z"�B�L�"p(�'|�4E٦�ձ.�I,}�����)i�b���+j�W�?�w�D�2�y��F���y�h::NL������t}:��eU�w��cvFա��a���N�I�
A��(MR��a�6%R��SW��o�K�&8�D5��v�i��q�^�Q��cD2%n��1&��!�EzQ!jȔ��)�B84�u(A�,S�:^�1}�BPH�l
��XR�v ~Q#Y� �ڰoU�UW8�ZNKPڞ;����fLSsX!��rG��t?AX�ik��N�ʫ*9�H`��Q�m��2lڅ�(��Q	���p�q�j����!4uT�d��.�J�(�g���w�������1�O����IY �B�U���D;w1�>BjR��}��LSL�qb���c�F��1�F�$���c*D!R��S�E+o�шs���+7�86���F��B�ҏ�V���rM���?4�b]ì*��.�2{��R�4�>M�Y�R]�NT��%�9]��[)�f����f�#�ЁH��ZV$ĄX��f#���@V�M����d-��ʲj� #�R4Z!��b��C�V�EAx�H�F���ܤt��&�宁��!S�/K94��NAȁ�e�52��:�1K׃�Zz6"� DS4�)_���r�rE����4Z�ߓ�?
�LFӚ��Ϟ-����V�oc9��Z�I�O�=	ו���D䢉��Uh�i��m��z@��m�5RV��m��Z�h]�����?��?���'?�id�i��ק�׏v����t�Z|��| GT]#�����;P�i�DbZ2\.'�,>ǘ�x�L| ��9�Ui!��O3�2|N���5�V�r�nk|!|N���tu+�ฎ(���Q�F���������U�ko|�[��������o^��ޟ�ϧ7����������[_�~��o���������W��/�~�ͯ��o�������/����o~�?����:��_��'?y[�������^���'������޽�>�hm���m�
YE�0�߈�d����L����8g�%CX!�ZBFw~�DR������
��w�!�:i�b�(d�o!Bu�A>���LEӪ��紖���D%��1�B��~"��p#��)�لD�F��C�{N݊�b��4+M�S�����G�����R�s�Q��g��4����S�c&��q�h}�I}n��!���60��[�N0+
��M|�+N�ˊ �Ǵغ2��^M��Z"��F:�ήV�-����cG�Sw�%4���L�0
�SQ��>����J4���0
F��ڔ�D���0#_�T��L?IA��;@M�^z�OѢ��ū�`�8DJ�T��X"�Dc:�8���H:��[V:��+4!H�栵��B��NdŁȥP{U4V��t%K�|)�F)�IS:>g�i:rs�D�BSd�.v!�D JO���-�}X%��4����`9P!x|�hH�F_ێ�/E03�6�rM�1-��	O<B�CZD�Z֞B�P:��X�}H�f���H�i���j���N?j��4+M��)2�6�4����R:�ң��f���B�3�� &��A!��E��a�̬��r�� �"L�YѬZ@4��m�#���Q^c3��DqC��v5M�,^i��5�k���HS�~�j-6���˅ ��7�-@����ՀYt�Z:��1���A�9�vD[�Q��8�c�g�y���ӥ�,�&!S=rj|k!(�`Kk]�c��/����N���:O�3N����ү#5
�1)L����r�֮(r�*�Ǐi-��3�  #�+
42�|&��(+>G����VWp���#$GR�ҁ��6Vw�em0�s S�1��7�1q���ҍpK0U7Z��N��&A05BZ�rƘ�4�R�c�RȬ�v�f����=��p���Xc�B�(�D�88^�v��?�uA,6fc�WZ3�pʐ*�����LI��pdS�h)INS�(�������z��Su�~ԛѫ�u��� h��$u�!�6=����cC����ᱢޠѪ�q�=�,    IDAT]_�xzq�kZ�^��\?;8�g�.�G���+[ڡ����V���Ֆ/����g�W�^��s��}I��k���*����>�x�b=DC�ysur|q�]�S��\�ӗ��9畨���|��vwt|�+jO�{(��:"�N?\���8���^�.�N_��*�+�|/;cuk��ڧDo?��������C��ۗ>�y���tاF�vy�E���������C��2@s-}{suU��ױ�NH�S/ɽ���%�W�}����5�H�z|�7��_ERB��LA�,��1$��vG��w9d}����u��@hR��J�Gc�Ԅ�9����-Ad�v��ߺ���o�t���ժ������u�ސ�
d�R�8޲x뭷�p
��yT�	�C"I�u�]�pS!H�4%8��&A�a�#����4m��*«�t�(��o�P��O8fxU��[�5&[��p��m�uI��ƚ$��R3JT҈֊$��BJ1:�Γ�M;��,.�!����t����r�0G��NgA��u�ꤟ 1U�{��d�[V's;�Q�s��NSi�V�l�R�Z�t�]�%Ŕ�+N�t4�"Y����o8���KA0�3d���*"�X��ADeq�ȉ�������%L���P-k�bMV.��M�d��4�de)Qn��u(�����)�\!�M���R�nzo��q�w=�Cr_��H�
�H`�H@�u��P���-C+��5$nIp�BFʤ��,��0!L�}L�y��.	�M�|��5+�OΙ���ӱ:��|�
!K�$�j?>�͍�ّ)�UA3�1U�sS�*�8����H1�dYp��i}BXY�W�]�(�G(}�	�[!S⢍��9�i�4j Y?��"D/`���$��`��y&�`�EV�~{K�>�i�aB�i:(t�����j)Fj�Q4}`A��9��i���v&�($qc��|�B�a���3��u9}#2���@����4��ye>��ҢR8M��7}�������m*J�%O��c�nM�C:F���)QbD&�VTTK��íR-��)8�H��b��T������	"�2D.�\�B| ���l��+*�N8���#� DQY�7�(e���S�H�(�)͔�i��ũ�����.��?����+)�`B�E��n����}��g!VAS
�谲�RQ�#t��[B�l��B�B��i��@k���!h�+�T�F����(G.�2d���%��l]���0��X��_M:���l��m��D�N��C�3F�2u[�2ÔN�[�/�=�ܽ��Ï��������?�������?;=z�_�����߾��Ϟ������1��ۋO>����.>�_`����7ߴ������s���>zv��>���GW�u�Y�]Q�������V��V�aS�l�u��DV�|�aj9���WF|R}��}'���Hb(t5P8t�p`��J��/�C���7�`2Յ"�|��F&^��.�D �gR�1Y��m���2�8|����Z8E�pp��!d~✦�����`:4�뜏ϟu�AଢF������%���YȨ�j�(�pc6���6⏈(2�T�H�\✐�A&�H����T��b�2H��\4�rb�F0gjq��4�6��*8:T�T:��zȷW]w�L�Xz�J��ҕ݆�I*_����#D��� hi@Ӗ�Xk��&��i�4�Z�M�l�j��h
�~�f�;�#�r�{��*�N`RF���z�t�.Y_�G��#� �����Yi=��22�越vR�(Q�h�@���`T�H*>���(�����{SK"3e���+a�g�B�tRU�`鵁�a�O�91ӯ�p��[[Q�p┧�%�1��F�B�����2q0��d��nL������(?���(ڈOA�T�e"C�
�OMil-s��%��hR(�����&�Ʀb�������;֥�I����7�J�ƇKa4��OB2LMLQ`�#���Ԍ9�@�j����8B�xE���CN$$M�i���i	"���8$��%IS����I���M���MY��B��Y�j����$A)#B�̡O�iYN-Sb��a[!�?QNj�8cr�2�An`4�h��B|��i
�0}�E�4���8D�R;o#!���d�˪�U��(OW�� �K�{)Y>��Ȑ��%&.ʱ�W=H�8�F���`rJ䫞�������356|N�ġ��W�V�jb:��;ل\�9�S��&�a�Y��>n*�T��:L�����)��# k	a��&��r�O�^�9ЎD�2?���JWQ�hd��8�-״N0�t�狢A�V��Ԫ�)��m5>ܔ��7����Y#��wH�]�N�C�s�>ɸ�+����j�on�;�?r�d=��ݯ�����v�����^��/t�B���������D�����n{�@��W����S��t9SY�J}�������8ӂ=�\���W�޿�䌚�V�/�\�?/��˓�'>��Y_q����p���V䷠UZ5�G���nv>�٩
q�eo�@u-���������x��۵L������S��<>p{�ng����9s��ƣͼt�hv}���=̓��밪a��P[�q �l�����-�ܚ���	Go��I��\4��,�ۛ?tY�Z�8�u�R�#�N��2��d��},��4Ei��ӣQ�j�ʈ/��KK�{&|�Oe�F�@/�ԕ�����z%E�����@�V����t��h�r�֭�a����#�L)W��z�2Up�XS����:j�k�S{1�m���q���6ÉfL�rEK�'�&��ٯn�6�1M�I/8�c����t�b;���eA�C"瓒�g��t��HϢu��iv(���;4)@��\qGٳ!��#T�,'��X'���I!�|Y�@1e�N�hm�)�D���Дāw�V]��ĻRЬǕRu�V�b�$Jq�&�ł�
NȝN�#�N4#2��J�C)�\����JT'.����z�e\��7� ��Hԡi�E�bODSFmt{�_�l�*��A`O�>��{hE=ڤs�]`��	�vi=@�[	69B:c5ԨK����_:Z�+FP��RJ4l��J4�eT��>��mY`O���ߗ[��[9�r5IJ3hp�t�B�bR㸹� 3r��k��� ;�Z)�h�MѤ�.Z�i�ik�L+�d�H�H��U�:�)�2�I�A��h����?\l�����a�%��OP��	vɛ���}�]���#O���wb�O_[�W�S��0���a�a��t,�]<[����B����b|8�Q����g���4��V�W]"�Z�
���T���S���J9���|#&5�h6Ӷ�^:1�1�R6�3�VR��(T�F0��c����s�:4��j@E)�)�@�8�u���C#���\|�(&Y�B��t��!���k��&P��ݩ�`zcDk�5��Ln�qB
�"�M��Ҧ����1e�i� 5��S�f��E�G�c��z���p�P�-�QT'm�=��ٳg�"�\���D%l�~FA-L�s��nPV�FM�'):�)G���p7l�M��h�r�r�BKn�G`)��|��H�I�-�,�)0�)
���J�X��s[�W�׈fd)��ڔs8��L	&��>u��w>����~�_����2���+��W�������E��YJD��'��w^4>���Q�����υ{|��h}���O^{�o��y꼻�^�T��F{����q�3zsڋ�EZ-����j�����7:)�Ѥ����mq��k�N��|[5�#kvd���%��tXY�,)EC�E��Д�OS��#4��F8B~C'=�	�'�"Bm�؀*����I3���|�蒬D+Łj�|j��C��8��p�J��=C6K�8k�i��	��u��5唘�G�+gd��N:)�LA�?�m�i&��=��P;��#�T��c����(�
5�4��h-%�4���J���a�0���׉�^��������D+J�oڙ�	јD�od�	����DS0�1S0�|H4���Ee�[`N�1�,)��0GS	;IҢ�7B"�~ c)M�WB��ϑ�O�M��)!���eq�*�&2R��� ����U�N>�r B�THK34�h�%��Z ����M�d�t i.��A��Xۍ�Z�g�I��4�t&w���h��mW���ny�ݪ[N�qB���SԈ@B��B�8R�*�/��6��E�,Nk\�{[':F��t"�(W�c�+�!uUԽˡ�� D-N)|_��16ݯ�op$�C��.��C�i�D�t����E�n�Gn��ArЌ|6ќ8p:h@��$��-�?S��G���%����1*���i��,�L]A"75��3"8��䇤Y'�l�.r�@Y�Ȣ~XЩ�Dm
Gk�!��B�K��V< &}�8Eۜ�Hgj� ��*rf3Ec)�'��Y+�F!
��K1%ň+g��72��X>�1g��G�.}B�+Z��PF~�Ux��Ws���/9#%}�S�Pd"�*�9dB�
1
�4�y��B����V���B�[����;+��B��e8Ʀ��@Y��O
b�b�3�*�Y! �\���*:k12��6�����[�EN��v�qL-J:�X����!�CDz#�S4Gh�t�l^G4M��t�J|�40dJמ�0���ԭ��>� g^�9�k���%�:sn��	>���y��{�z����]b]����T:v��n<T�C��T��>Q����f��<��d���G��Mu������8}U�v�Qq�-%oO�N�G������w�f�ܼ������ӻ/^�3�^�̨&H��������n}�Թ��Om�����?�̎�'n�����z���i#�Ο>����+O�w�W��W�~����v{��L}��߽['�:Gn^y>��������.w뤺���Ձ�v/��. �v�:��NV''�1YRʚ��Ǣ�2�D!}�S�;W���*���7M;��H��� F������z�3
�*��"C�����u(E	/iU���;0>4E�BZ;���o����d�Gi���SoA+WE+eR,�H���!Bu['|����p�p�$r&a����'>#�6RH͈���%8R����p�DHd�� �Ԥ*IA���SiӔ9%��w�(�^"�\r��`:E!eO��I1d�F8Y�ϯA������D�h��l��Nf�|��!O]馢qrv�6�ajbd]�@L�8)>��фR���!���"r�C�(�s���|��E�GoޯuQ�Lǔ��JD��҅ ����p4/�QnWV+�C�|K��9u������JAÇ��C^��~)���0�. ��<�~�X���ޘs�ު��/���������u[��G[��G�c��P���Dh[u�KZ{Q�,��J�o��f8eS��Ӧ�;SYubBDdY�ƪ�1���EUg:����D�ٲL�H@�6dq������~��I!�I��
m�M�jd1�(��H�Hc!�}Z&q~+�d%�c�O�~)��U�*�J�R���L�]��Y���k�6��N�);�]Dh�љ��,u-���p�)�!ȝ%C��M��A]Lu�E��g8p4
p�$"����ld�p�h��ZF��f�шp�F �Ȫ��N��3R6aە�w�m�5l��JH�`*e�e��y4̖@V)�öC�o��Idm�J�VᦪT�L�@���mZc�#��� �H��.���Y��I�5�@m�rNN���\#~7u�cB�ҭ�Z��(K]4���#�o以Jd���fl�Mg����G:���_S"FQx7^��@A�X��e�ٙw�y�X�#�=�>vzx�is�W׎	�I~����?����(Yj�zC��,�Ĭ����7�r��$"1�K8D�M�J쇪b�~F<���v��`��Hh�hjq�I��nE!��	����ﯯ���<>={r���9���J�=�}��W����"�}�K������Ro_?�;s|��{����v�a7v���Z���ɣ�pЭ�ft�1����FY�vg2N|#ki@��	�NNܫg`�����*j�*�#���떟ID��*Q��07��+���8�4�HG�,Z����V9�g� mHY�Ԍ���?)�g�JM���3R)�A(�p8���Q9�Y�P��m����O��%�¡�L�b��1��6��)�Z=@��⧹�6�1�3$|J�Hiɣ0S�4�~���1�α�j!�A������(�1�΁r[`|�(e�4e�̆4�(�c,w����:�Z�d����R�:1�0�B6��!�hY�tD����Ú��~K���	�)QV���L"|.+~]E�
~���
���G׽�H�eU773DdVC7H���Ȅ$ F�)�o��	BB0@HUR�cЈ�*UeF�?��w��}��{C��g�����k��캙sF�c�����Zj*+���l�P��;v|6�Q0��B*]�P4NӖ���Pk�8�3�iV��RXE�G���D�!Z~�}
$0�Sic!���>�S����D�#XQ�Rࢥ���s22Em�pF��,�mWu�T�I�h�X�IS�Z@F�t��@$
E*jL6�)M�8rC�l��&qR����GMH'�1&|���K���KpRʚ�D�����
�H45����/X��6���1�Gmr�Ԥ�/7��C���?f�|�_��&�����9C�6ڨp��M�%
�ڋ�X-c�@̺-���D ��tH�L���P�#��&D.e`W$��7Z�S�ŧ9#���S"e���)U	`U��hkڈ�I����!F)p�U7����9BI�
���p�WO���d�I'_T�T�#4
��S���LK�����L9�S72Q�50���r�jj���T�1~"h@c�*]�)D���bj�t!�%���	��0)�cV�i�@��J����@s�ᛢ�R�-om)�Ùf�L�iJa��|��*���~�9�X���%��Me�Ek)�T����+h������k)���p�FSc �7���ȋP��bդD���V�f���F�G3հQ������(��-�h9~�RE5�_�9K���ר���\$Y{�~ e]��׿]Td��/��������g�`H)�Y�֢���)P/�}�m���Z�&0�/^��ޜ������__�o�O�ki}������%��h�\͝�>ys��_����w�޹w�/��},�r���(O�8�`�\F���II�>X�r�,p���[x�/��n�^���~���?����G�8{�N�������p^?⹾D˯���f�!�V�i��g�ب���_�w��Ѵ�U�hmEGʈ��St������C:��l�Ǉ�:!9�H�I99�pD�xۧ�*Fg�r��9s��_�h��A@sFyKJ�6�3��Y#��Z�_��_��S7��@��M>>Uo�)�sU��Sfxm��c��ʍ��u�6e\Q�D�8�
���*���E!5'8��56}E3ULkC�18{�5�O��8�Ư�|�$rTa��Ƭ�c�FN�ڔV�ߔB��Q��BF>���>m���r�`�L?sD�� I-Z�B�M������C�iu��6�%"�ґ�)�_�Z���!�r���-��r�s�{�wG�M)�L���ޛ��CY��AJ�G��c�x׳Zm�t�1K�i��#ۨĴ7�KY!��|)FS��tE�� M��*rL)�!D\XҜB@Q"@��hj��H�+��Iڄ�}�{t\R��J�6���_B��G��i߶��ť幀�d�iT*�H��G�Mm�Z�͍,wփP�B�Sp �#� ��R�l��,= Y"��F�FL#54�����9S���1ml���BU�S������ �҉Q!=Wwk��_u��	��!>2e�V���h��4���r�BU1e��c$U� �%G�n���U�F��zsrzB��Z���i��I����Ϝ-���� ��AP1�=WԎQk�-�֒6X��=Q:��R�Ԛ�@"�C�ht�?� Z�t�p!6jӼ�0RF�3��mc�5�����    IDAT���0��8��S�t,< �DHGt��O=���&��T�UQc|���8F;��@�A�s6�5Țn�1���6M��IvZ�3��G"PEx>��@�Չބ�Ľb�R�N����!2���(������ZJ�f4O��Z��Bʥ�i�d�v�/��D-(�S;fj!V�T�<��U�6H�g�h�\U:���o�磥E��a��&m�Ǧ*R�jC?�s��{�2�|�:�**a�bd�!E�b�o�
B��ZZ�	��r�tT�t��h���/=�z�b�l�ѥ�z�[�����.]���c�$�(�M-:S­ǓWtG�z�����x����m7O~���߶�/7�����oln\�|����z���ky�|�@��\=��?�O��E`�1F��M5i4i����(QL����������yg���q�Ǵ	@�`��Q.㝺m���P���B�7���53|)���B��+Ԉ�aV:�_�������S ��ɏO9X����V�CQ��BB�q�*��c�Գ�\�$�+�)::���M-3��$"4�
���IQ��r����p#�\���n:k���N(ܔ񍢲�KVk�6RW��=7���7��f,dd��p��#�`R�2qY@��``c���c�<A!�	��+Ԕ�1N=�X�h��t:ALK���Ǆ����#�C0mQ!e�?�-��P��}�����%�>j{�(9�t+u�k 5#>0�d��)�fu�~=�S>���@j#��՞�|I�BX4xK4�ԚR�\��g#���6�H�Ȥ@5H���_E#������Z�R	#+�c	��#eO�[�^-�Z�)H��7~��B�1�9� ��M�&+���R������� �,���m{�<!���۱�'��O
'��3!�iW0N�Q�JCl)�'elڊL��'�~X;,�C��k�i�=^����҅�'8�B����H�k`���H|cʥ�қ�0�\B�7B&e@��n[H�ٴ@L��H]��)'����A�c$eT�(Y���-}L�!��b:\����ҍ!�s2��GN*�ٱ)�:��	���#"e
����FĔcEt[�s隆�B��*T]�S"��K}ӇG6�1:��Mu�,?q��ȅ�F4)S���3?��J�E;�� ���)�Vq�ӕQ|�,�!ȂGgI���A쏱t|&qj��@mt���hl-`�q�.DH�h�� ,��L��@��F����8���4�ՠ4;|Qoh�����eI?�)\z�BxL!�tXi�&T
_	Y�@>-�t�p#5b"���m{k�4B��Z��+j,DĿ�����떃��o�Չ[�[��5���.�%��^]��nU_7��"��R���W����ڏ������S�~�r[�IK���|t�ӟ��o�u3r��}i�}ț������+g/����8�?���kg���gg��������'�h����v}m��v�Xu����y��<ׇ=�k��;l�>
���ڍm��>Y�#�F�z�����B��_����.O�won�O�붪��}���_}E���ݹ냣OO2��<O��'�[�|u�r���Ys��r&�,�ۤ���qĽ��r�1��Bz��qW��$.�Q��f�:p3L�}�N3������n�����}c�w	L�6oU��>��.%e��M��گ����J��&5�v��U�Cmz�2��Y�)[Mo'y@~!��j�q��L�][����i�/�c�9�1�0x���[��i,�"��\��מS����cV~E1G_��*4�ĄC�D�tL�FÙ��F"p�6��Li�fYU�zc{�/���WHbH����\jF��
UȐMCj�Wȴ,Ӎ�+��OGE�)��X�|N��g5,B�����U�,��z�r�:Qe���Ǧ)C�r���P� HK��x�TK��B�N3�pU �����i�n�R��JPv���B�J(�SȬe��4��}�,�/�n9�T.��h�8���F���K�taA��"�F|�;�Z�����?�X�!�����DIHn�HÆX�(_%S5�C�M�)�����1my~4!S��B�M�ZR���{�^����#��}m4�P!��"�C>�^S��p�@R�����8��f�:ZS�CD���J��.)p�t|�
5�O�����D��-%2!S�i`�1#�Xu=l����jElE{�A�7�,�nL�hvF�~�����Y�'9�G&�K����v���UL>Pz)���fL#Pp��4�K�`J�[)g��Yx%p���)H�`�I���t�Z��\WMр�B�@�f4~�8�ǚ��B"}"NW��m��Ǉoy�_�d�Ǩ�U��=i�Mm~�J����kc�:V?�{�%ԡhk	�\���c�zn!���Vq��Ƈq**d�D�NEW��th���'+��Od�D8��u�AŊ���Z��O;�K'Aa����n&Du.D�&  ]C�m�,2D�,5|L��3у�i`"H�-4�-B
�C�����":BUo[�p���b�[]��%JG����F~���(�!<5cLcm@Ц"�B�,��r�8)DNĞt���Q6-)��)�Ub��T��Z�������z�9�~��p��2��3��P�
�t��������h3�k?,B�Kƛ�����^yN }p��;������Y��ji[���z�;�h6'�5ֳq����t_D�Y���%eng�4��W����DLS�Ԓt�����D#p�
�cdBiMU� �+�;
�M�Y����|4�[۝3��f�`�Q42GQx���.7��
Y��G ��hu����	���Q�T�K��,�BI�̇K,�r4�|�D�q �˯(�45)q�|s���4��S"gߏiF�;���������V!����n�aVor�dBe2���t�M�i
UAp�LbUH�����L)sA���ï�RQ��h�l�BBG{���s�D��9B-s�B@N2�q�Ogd9*E��'�BʂW�a���E��3D4�#Toq�M���8��<?��>rLS��_'�����'�Z�d�t�K���p����(Q7$�αR��|c��IhZ([��Zq:[*��\Q�C��8���c D@�����s >��`�%�9�ė�3
1!�A��Ѥ�r�*1E�!M���v�h\�0M��t�0�ȦV�hĩA�:2��H9�SQ�#�nM�D�V��N���'F�2��a�#�4x��L�7�3m�PV�h5ϗ�8�p4�ˢ0�)aJ�ӚB( t�8�k[bYJ��B��5BdA�2��_t�S�ԒX����K+�VE9�L�Ө\m� K):U��J'��4�=h
�O�O����BPT��a::m �s0�)L�i~]�g���|�B���QqV7�7
1���'X�he�U#���H�il{���d�m�3��D�6=ԕhL�i�����"�t�%���"�"H�hҁ9���!����rc|�:rL�Vp�0C5���R��N����	
M��s��Sk��U��/q���.���)�OA{B|)�RS��r���L�?P˂TEb�)s41�J@��r:X���5�M�Z�#h
�Uј����G�@�TT�rc�E)H!2�D�h����n��o!J�#txz�*s��sGs�ji}G�������!W{�><����f�|q��32��"�Q듖O�{������"�B��]����Ϯ�4��j�~�� x��)�����N�x�����wni�=*���>��w����罻�~~�O�\���EO_�X�9Ո�^�+��ͣ��<��5�2�I� =^NzX��Q�f�޵
����{z��1Q���w�|��/��z����~�G�<���Ý���%���ᝏ�zA�����|u����g[��g=�3���%Q[m��c�T�̼�∬�z����ܻ.�����G�gr��Z���:e�?��"��DZ���E�K��"A�Q	�߇���W���] 7�m�3OF��ea��}JY����^o=!�MHch5��T�ޗ@6�')�9��DhZ�Fm�3������!��|Lc[a�@QU0�djO�66��j#��9B��A��MC��~":���q�!8��$k4����B�6�P.�~LqZfjd˭��������D#��	MG���u%%5�p:�4�a�L9��?)pMg��@4��j!L�&����8u���0�V�O��vEK
s�XC�s��� 1�R�N�d!>���v��*�TG3zDx z�y@�-�?��%�ۼ��qǯ�DS&������t1�����U��q���K����{�܈L�o�6�
�%���Ł��b���!h��ՙ��E��i
!ng�]�05	!��{yD~���nQ�)����m��Q�������U%Z���5_�47�(VB{�T�t|��]sm������/7r|��h	nd��v�@:���~�}�P���B"��&A��z��r��Ƨ���H�M�˽;�n���F��]�Чf����i�#�"K7��r��8�a�����8>�-��zjJ��ʕ���-��
�4���4C�iK{z���_|a�<��+�6�&wz�@K�n�������O���Ąw�(�;��L"Z��X���jb�(r`���p Ǩ�Mu"%A��0Ј�CˆT7G��Fm4�J,HJ!d�@���	�]F�әO_{h)�����!B.�9��r%�,�(��Ǌ�8�_��q�r���V��kE93��1%+��q��\�[����)��CL~�"|͈��^�](2��iS�7���U��Y�)�X�6��T�X�Ȭ�/ZW56~��%W^���0;X�4]�|�,YW$m���-BF�G�����,}��챼����+Y�Bӡ(Ĵ���q����[N|�i���0s�ZZ���d�Ѫ�b�J�T823e�dK�E�����5�8��W�(�3���,%�)���[�T��=z�d�|ύ�B+y���P�7?�,Z�����
��zݐ���8�
߾��+����g�Zk�V9��6G����K�m�M��c�Pk���DH�=׉g7Wo��,4�L��KwR@&�j�C\5 ��1�vy!1�b�|�( C�(�V�Q����T�cS8C�X_��m�moZ?�{���\� �-���Ĕ���~����b5PԔCD9~��e��q���rc-��k���E4]]�>*m���P &���R -��_�ĔcM5il��Z"L��	a�%KK�P�5I$f-�lө�_��OLњQN����
�&���8�ȩ�a|�VQ�ǯ.~Eei �M��Q	a��)��a���f��ǟ��2E�ޤ�Z�)ͪ�f���0Sc����
em��zJWGhL�Τ/��őU9`
�'5~Rdk�/Z9Ӑ=�\H�j!W4�A]'��5�� 4�8�^�G��V�_{FѪ�dt���^�s�jX�D��M�MB �B8��|�P�	�B&��T�\�m�'�BEӄ�eҕ�8���8�^.�=��⇘2"@>�GpN�Y2:@�/+fG_hV!��YVR�ь�'\3�##D�Վ��.Z�ɕG]�P�6�,�J'� s0M�8Q���M0})3My�(3
q��5mϓ5����$�9U�CG(�Y�>K�Y>M&T���Ԁ�49�8v�=ĄO�G:�+��_t���;��R��Tt�='b� d�ⷷm�iՁ���Ս�N�)[��{�B��߈IP�#����-�_oi6ͯ���bD#k���4��8ҫN�c_.a����XӜ�}4�����SŚ\Bە�>/���%�oR�κ�����gz��F Z�����#qb�V�(eJ�V"G
���Gf��堑*�4d�Ht�+��oY��[�$�oo��D��8"�SN�_���9���!��,Լ���rtRc��G�$)�� �I�h�/��bĤ@�&�L�^�k,Y�����|S���L�Q����N��8n"�ڷG�I�7������ÃǕ}zrK�B�k!d|ݐ����/|
�m�ӵ�Լ�t�r�т.~�����w����o[ʴ�K8]���·���~�iJ?����w�����������-M���nz�^�׺>\��|����}��*����e���������\��w=�|����&�|���[u�돏��(�4��M��M�Ս���O�s�V��z��O���/��
7'�����~����t{w��V_ʴǇ��ݸ�ۓߤ�n�xs�į�(y�����q,�a�xy/�Tc���d|�������g��ӻ���{�}lN'���n�\9��1eަ6�*�Ӄ�����22*�o❄:M�����Ϊt~z�H���xd��z���X:��� �|�j΁	�)d���d��Q��Ԙ8GJ�q,�)5E9h�*�MY>����7|8�B9pN��9�p�C����FVif�SPa�i����Bۙ!��P`E�BYH���M���n|�u��B�BN�)�_:�ρ+AnLv8�N�e�ld6�,~�҉Gh���ǉ��D�o�;`����)2�i�������CQ�4�h�H�p ���Dҽak�t4! 2M�&K������2�][�y��w�<�GzU�#e!�t��@!S=��e'��t�GӭQ����Jl��$����Ԋߵ��~�ҩy�����\�D��ȕ���G����{�������U��lYm��K��V���}+�Z��G����u�F����0�R��'Y>)#����w둸;�|Q��v�rD����Ǟ'�4�����g�g�o� ��p�,�s�g�}�]`=|�嗝g5���۴p��iu��Q+)1�J�cD�H#ā��b4e8�L����C$n���~r�!B�H�L����>�F/YU�BN#۫���r���F8�}[j�l��������()�Fu9dф�=�ф�ag�:��Y�j��CD��ΤXHQ�1%�P�`�h%��5���#�լ�rE�
�C�B|NU"Y:d���!�M��0:ٚR`5c�9	�DB$Y"�zCⴱ!p}v�H����ɨ��{�8hr)0��s��ȕ#nR����j��D�ǬB5CS3��JA�����!���Z�U��x�R3[kk��J���%[H{@�d�U��#Ԋ��E��iC&=������¢(ZE�]�R�Zk!.ݟY��s_���8�E��65QMbB�9S�'�lfJYԘ��9B��(
���4��I6��J$�S���E˪�F_j�I�b�7Y�BôR��������_�7�dc�B=.�LgE�U4B
� �l�U�&s@����QS#�}���/��I�L��5�?>ݞ�R��B��(
ɀ�m�C�4F&�AC�T��il����v�hN	!��ҷ(�yY����4�%��h�rՍV?85�j�~:)���Sz����������«�\>r��,G��`4#D�t*��-+�4)�#+�� |�Vn�!:B�h8��p�	E.:��Pp���&��*�� �C"�Bү��+7#'r)�XYD���=R����#�3Yd`b)�un���+ms�J	�)W�/]!~�I�2!�z�VBǈyI�GM?p�Ќ�F!Ɓ6��L��L!��G ���-mj������1M��h�*�i�)�1�58�U�[���9΢8�:�oT:	m�>1A�$(J$>�����V!�*�2!
�|&ݸJnE�9��RӍ�rJD� ��0�r�>�����TB"�I\]�VKʦ��Ω�:��4�MNp�L��FF܈�l$hu���8�(�N�0?5#��m��
?A~�US&e���i����*�vL�#:���L�H�i,�i���d�f�>�D��Bp�~�h'XmtX���*�-_:_r���������A(Y����kCDq�M�� �ƒ5�g�i�`-i������Mo��.
ID�&����1E��#��4�Q�������ȡ`�i�?iB:Xg]��4�9�a�,r|c�ƚ'5�k�q�G���#���&��ȅ��T>uKTz�^K��Z��p�0�4��A�N벓��fJvhp��,LYSȘ.7&�cj�1�'�F3�B����ƆO    IDAT��&X"?~cS>�_���8REE�C�X��1S��1M1q���qJl41qR(i���Z% p)���(0!Gb"��Ȳ�ZFY�MUߔ�Y�逛�Zrd
N�!�^W|�,���4)��p�L�B�N�*F0*ڵ��d>$5
����W�T'L
>AL!���*4]	�1��YW�)Hd�]��Fo�q�d1g�ҥMk'\!dcxu�ȅR��Zޝ���?_��7w���=��85�Yq�-���77�ۭć+�����;?�)�xX�OnD�����^�ۣOdN�7��v��{�x��-�������4^�?�_�j{s}���o��������Oo|��p8?<]�}~���G-/�t���^؁X_W{����yU������|�;����Hn���3�nj���Úk�k�]�\N<�D��S���o߯���̉�	���'�q�W�"�ֽY7Jon{�p8�};?�|�?޿��ه�ӣ{�t��2��;A���}���(��r���F���	��z�wt��;�~T��r �:�6oݭ��;�g�S��S��r���	9:�hĽ���<��'�����A�&�;O�)�\)F>���Jx���A�_��A�B�U)~"C��lIۑ۞;ʕ���ϑ8�d�����kXV�P�f���B�t�'ȏ�"�ьĜ������OTb�������W�6�Z/�W7��JPb!:� �úe���v���`!�	�7������'�X����_�1�^��pZ'~;��O�B|��׮
��YN�M�Z�hꑅ��-�R��B�q��G��)�]J!�j��Q��i�Pu)@�0$��
�V���F!d���� �& �l�hVatY�$"��"�e�����zkK�Y�h�����,)�f��7��yKP��N��w*����wt���]6��ﳍ~�����nu�|^��z�֪��L �b���?i|!�8�h-Bj��ė���Bj�HLPb*�~4
�XL���K�`Un�9N�޼�cB��~T�b�kn�v�O��O~��~�yf�*Z{|�h��UW���HJ���9�H��0�ۄ�L���uEȁ38˩hY*��S��cB��'�P'e:U��o����ҿ���3:Kl��J����i�D������~��?��_��_v��JM�\���T�.�1��Ɓ(�>��ۚ�(�o,�7�E|�L.�Qu=���r�|�,�)K����!ASg�Ҧղ�����E��U��	id!:���(�jx��s ����~�k����F�eW+��9p���h�*�(��iWņ0���hu�rZ�DY��p��D�V�`
�'�I��+M��2[��~�r]��-����S� �C���8k�Q�(]��tdm�
���1%2�#�o!Mq FF�kKݖk�hZ���QT�B�y��|�Dg�(A�t�B�z�SoVW�����XuG��p�r�T}����F�,|&����D
�h	
a6jF��4}�4��/�Zc��Q��t��SB�廂��[D*���CBM��%�/��Z`�n��I�����=1�|�BD��|Y/N���H_��6�E��(��Ԉ�y�h���e-�v��"GT
����������=��@T�bj[*Y��� ۱ZU(�iEE9��(�2�΋FʙR��Mp�j�(�a�;�-v�1e|Q��drGYA��RL���D��T������R����l8|kp���T˸e�!��ͩ��hU$����V9�1C��W��&]4�����f(EQ��-a"bD6�h�7�k��fa;�� Z
8����M�V-J�t~4�(r��(Nju�%���P��l�l�U�Τ�U:�/�Cj#��׃P4HL��Gp�,�,YQ��~�G4M���R*ʏ.��ZL�΁�3[�^�;.B���J$�a��C�K��@�үm"�hI��QiQ�1Mٴ�B�V޾��Q+��!���(�~9�U�?ѩ�cEk����h��ȅ�@�TȔ!E�lZ�O!_�>9ɦ̇fSݦ\{@��1jF�����1'�
QP��(�,'�ZhF�ɼӦ8�5���4��E.dT"���1M�bD�6��5����#TAV~�u�O9�8C�PS4��ld�9lB|�u%�g�3F�\ۢ���5>m��M�E��k;��mj	��i:SK(D:�0�bZ1��:�p>���C��C6<^3uDs��w>p�Cο����	&'5>e�����FLqV�R�S�(�(|u�Y�E�Tap�t�u���+��DU$r�*�5��M[x̖��X�BhF'+��Be�88g:����¡od	r ��| �:l	Ӊ����XV�%�L�)�J!'�*�����!��z����s�`�>$NN
Bq�ܐRLF9�ή&"*T]c����_�>�i�)�C�BƔ��L4����)t�����ȑR�l5�&a9�D0{e�W�($�`H��*Z�D��
MujR��|OX�r��G
Ĉ'�JC��j���S�,P�\�,�3�)�nů�L�[(����w~^4�WS6��MM�ok�0��g� ���mq/�>��3��Y�K;gI�>���^<���;KZ�-��t|vˑ�׾��x{���H_Q{�z������ ����Փ{��_���������[��K�����3��Ǉ��>�yn?������)R����f}����%χ��={��t�}	��uZ�/���n��`�i���{�+0���Z�uoTl�*�1.�7n���\������S/��E�����tsq�֢��\7g7@o���:�~��S����t���i]�}���/и�#��N�u�Vg���}���h�y���E�ވ��?�ӿ����˿�K4!�w����mX:VM��������/���X\�ѹ�ֳ�+��� �;d�+�����r��NP���
u�%ha�v���N-:�N�B�^,p����-���89FV:NS#N��:Q7��JZj���qB�NYB�0)*}z�(��9
�ۦ)�=1�&�^��4�2M� ��ϙB�Y4�ү.sBe�Ʃ���Pu���D�R��d�A�����^�WW��$�*�&�+a�O�r�jq��8r맑rj��6$f��
!R��+��ԅ����0�2�	M�
�krV�����j�s�n�x��!�A큟�D�ՠ�H�ј� ���&�ʃ����t~�e�2�\�$�H�s\%���žg�!HM�lQ������#s���F+��Tn�F��J7rݣ�bH�rܧRY�8폷�]�*��M�`	6v���~�7���P���d����t]��*�2Z�t�rp>bT�(=�:fEE�SȂ�aZ�6t�eU�R�=�D�CԀ��k��}g��$e��	�Y΃�R�4������U����F��nڎ�eʪˁ�-�3[$��Ɵ} �_:�t�c�8�|765"���%�g���+�T�J�w�}o�����q�p�n�����d����F�X���]m]�I�>���ڮ�8����~i�����=�4D
�M~)kT�X��75�K�r��M����IE�I7v�b���RZE��!�-{/�Hyu�~��U���n�1S[m�z��� m��֫����k��M)�2"sE�u2�m�8p&��p�@Z#?�_Byj��DhB��Z/'�Q�(j��r�%e�B,Y�!6��5_\��N͏T�4�Cɉ/�Z%��QN�I�Y�}ӹ\S"B�B]��r�D���f�JGJ���?��o8�;!kIn���v��8&K���Ճ�,>��lPL������(2d��O!�h���r95(��_3E��`��L�zK�����W�����1�����Ƕ���!�˅f�*"Ad).B�y���?��o�J�P������ۋ8��a���]��v�C`��::v8�=�B���dN�ьC��?z�d�j�JH�A�u5��w��-����R� �9#���'WV�5���S��C�p1E��p
5-� 5���:���-�4&W
���Rf*!4@�S�1��&��d�j�e�ӧ(<2~�)��M'E!��0�!�⯒�Ç�O��� #<��p�fbjfO�lN��k,0��(�C���vL!>ٔM�P��|S)��S��_�t8@N��(�AZ��L-)!��6�D�.c��6�&�fJi	u�����Id��������U�D#é+LH#��t+į7~�r�C3-=�}阑��S�Ui[D�K���(���\V������I1e1���l��Z~LcR�!C�/�B� ��o�h����4
5JWH���,H
�\W�� �LVg���J#�����B��0Y����D�4��^��!�B�/Z��V�"�R3JaC�����d�Z��p�B�d�x!�Օ��t��IAJ�����u�4�hmW!2!�b��q�z��p"K7BАG���@><�D�D��0�)����[�FSR.�Mi>rg�Kb����)p�����a`��-�8|Q8�1_�EA�j9u�<���Mh�Ӡ�^))@jƔ,�W�f��4�Y
>G���L�a�<G��%��i!�r�"�R��Y{ed��S�Ҧ�!e�!0�h=�ME\�����U�ʧ��t+��J��S0m+���r6`���t���C�V���݃ME9k]T�z R�&��9MGĔ/��3٩�c��6�D6���L��8�2��N�6͙,T-ю f G�	g[� ��Է#�ߴ,�Y�w;Ï�6N
&)�k9*�D�� �o�k?���9��9���4�?mO�8���aڨ
BE��봞m��M���%�)/�P�h��t�͟*���8�
��֪kL:'��h��I̚$�`��\����6&D��Eǜ+~ ���U]��X�/�����u�y��������̫֝���n�Z��󃟱t+��3}N���㛻{�A��'o]��W��a��=�2��z\}���wɺ�����{���A���z����'?}�ɻ�_}��㜾~�����޽��~��}P��]y�������|c�����Y?j9ʹ�z�ݵ�a�Oj�ӵ?����!�������[_�ֱv��������_����r�V���S;E�����`o߸�{�j�Й=�w��>�����\� ����z����z�2�B{՝��}�{d%�><�uԺm�Miߒ�S��ޥ�Ճ�R�k*k�=?���#+��	�����W��M �u�_��4�{��t�J�Sx��G��Kj�&���b��v�A턄�h��)G3�U�(�>��X�M�(��ѯ����IB��aJ�Dko�z3V�ä�����aL�\'�뿋Lk��\JR!!���Z� !pH�jŬG�S�~������Cy�Q�u�B�]�D$r�t%jGT"���!B�1#p�̱9p`�g����J?�J{�Di~){N��I!?G��rM�N�_�uqbr؜�S�&'���=do��s�p��l�;/�JD���֨%Rdǝ����L�O���H��Io<��i��Ǿ�>�g�}��䵒�^���u�}��^7_�<D�-�CA9�V�()�E1EK�ɟsS���)�2L`ozS�,
��C�X�W�n��X74���1���pvy������UU���(�Q[N�Vbh$dU9�v!PI!>���E�o!Y�lRDUO-��1s`S�eth��k9�є��o٤�0dQd ��1��o��ow���:�� ۖ���1ȆG Y���Y���(�q�v[-�|���	�	,+PE`m��a&�~�+GYTE�mQ��d�<�z�@�ǡ����n���,���;ѧ�K"u��"�c�nc�Mq*]�pH��̔��Ө5��Q��,�,�+m���m�,K�&�g����0&Db�E�,4�*BX)8�Η�����g�t%�SU��h�� M�(���EG�Z�D YN�L�2�N'r�e�k$��\~}�OM��D�"�)3E0�9�x��!N6���e��?BD���K���IY�5,���oi-��'�n�
Q��8Ԣ��kۈ a�~�4�1u�����H\�V!4����G�f��@�T�T˔�@���DI׀V=i��d�p���N�SZE�49v9M(�/dʴ���L��pb��磉V%�ZJ�Z�8�b@��'����8p�Zd��
g����G�˅;����<�X�Jđ�f�KT�y�pS���l��e�]]!���:(�k)�~4�`!$BP!cG�_��n+W�B��Vk���!������64���|���Yc� �f�յ�����/�_R FHc��M��`>��e�p~�q�����RWn�eq4�4ah%R�0NQj�4�O	�ꖒlm$(+��4�IM?��t/�iJоuP u^�)bDc�t�ۙ�~m�fT�V�rh4�~B����)�.���(�0�(��T����Mc�ED���M���c�i��B���Ԥ��hJ�C+�Hm��©�|SF�B�4bZ]�������*�&���ê��:aZ;�I�W-Q%��q���"��߷a*K:'B
�:4�d��fʧ�c���өU��YHzuU�TȈ��	�q�kJ'�RV�F��J��(ge����D�E��m��kU(Z�B�S��E�o�ܡ��'Q�ǯS�o�3��x�Z�g�s�MX��"�R��G��!1e�ӿ��!�q��B2LΌ�����2uC098�����(�g!L�����@~&ĩ
ܔEH9YLW�u-��)�T���HS�r!���@c����l�FaG�N�ȢL�X��L�0�@"s�@C��B��r��B�8��Us��s:��"��(��A�|�f�)��i�E�	�Ԟh`]�i��� D6�bL�P�!R�l�4C���u� )�xS>GK�M��pS׍��'�" 9K��^���>�,�XQ�@��M�jI�I��4Bf�)'�?�y�-�����!��&e�7��D���;�����L�$%0�4�%H�@֢HM�p�ԃ�To��Rp�!l�|9+��%z9 �<���|���J�W"GQ����T�T����%B�,`��.���Z��B���gi�@Ȭ��i)w�M��*jRo�b���T��0�����&p�\8)##�d�Ҝ
����[B��f!d'yj�%2�&[$N�����Nv���)C�c����K]���|M�wкy��S}���u��dI]֒e=|��i��v}v��@������.-qw@���>飖n,n��O�7ww�~�O`�/�o}�Ư]��}O'�ɏU��>���}g���������'�No�|pC�����֪��0�짷�_~�7>O�ھi���܊^�׋��\-��Ϻ�\�\���O���>:�̷̮;�n����ѻ�o�~����߈���Z��.�u�����N?�y{<ݝo������/��?������\���|�:���:|��G�9�{u��g�}�<\��G�qm��\�X�j��p�O
_�f�<ā�����ڿ������w��xWAAV9������R���o�������������[���%���,��e���C��Rb�ޞ:�Y+m*W֦��Ml!R�F4����3:�IM:G�Ȥ�D&NS(ΐ%Y��#�QV��s�ɶ:��Z�i#3%(j�	���
��S�O�Ô�� ��Hm�3~�ƙ�B8�=� P�X�q ���!$J�$��D�nDF0�Y�8��T��~9d����e�R�B�ф����T4�h�
��,���=)i�2!�z��J�P`�n�y�����2%��؛�|!R�J �"�����dnoy�2j��+ˣ���~����E�K
�+5��u"�[�ڦ\�r�ּ���%+�0�L-S8���2B�,&���K�Ékl=�m[��ַ&q\0��ʱ{�����i�q������B\���!۝*$�Ϻ�A���1�1�3��XЙ,�h���� 1m�9@
r���8ɖ��!(o�L9�]bzj�?��4ו�s�)t��2�uU�����3����78�4�KJ��SJ>�v�g��C�� +:YRA�,!S8��3��Û���JJ�S+'2�a��R�o�n�q�t    IDAT=�9����*��d'�@>�#đ��jd�)Q'L
8N1vⶱȖ��+m0QS4�Lϭ��Z_
���Q0��5L*�>k��%Q%DuȇpLK�����࢔!�S�b|%��DS���d
����h�(����9ԭ\H�8t��>M�����X��g�tD9��bqXݢM;�WԸ����R./�B��e|L���%H�˙(H��Cn�D�S㓕��*m-q��+T]Y	�0f=�>�,��h�R�t�Ϣ(�%��r�z�鍡1R�Q:BF�#�3�4��d�*�(ǒ� �$��a�
�G�j�L�,���o���t��oG��9�jL�@�_H!��6�T�h,Eh����ɢ�#�p��T]u|�8��M��W����&K(r|�*�i�<��:Fh�ğ�xґn�_|�gb|�\��a�Ig
A�H'd�\�2x=@�@P�qOJŤFpZ�D-1�t�9I<�ScȣL�C �:$�sN��a�{�E5�ъ�>��
��5�)Y��f��Sz!|�L6���p:C�GH��B�bY�DM0|�'�΍k4&Z��S�\
�Wq�@U�[/�QcE�R��V��p
%����,��0��)�/��7�G &���)��'ܴ�8pL`�5Pn�S����i�8eM.�h��F��Js��C�n���|Hʘ�� ��%��_"Y:���mu�՚N�5qR�nJ�� [���M���B�%TRݦ���Ȗ˩sQ�19�de�Dj))����-~QӲ��\N�XѦh�8�7E(e*�&��e���(HO�/^i�i�\�J4�R�R�����CV�i#�U���`Jgz��0�@4�U	�m�(|d戛2|mpZ���-Z�^�zK�YD'Ïl�f�`�S×����fYCVB�&I����fV�cN8G眲8
�
a��ܴZB�
Q�)0��fi9F��	� G
b�R�#Lp;,TB��|L�5օ�(Y�HY�o	
)�	��P҃i��(�,7�s~�R��#1�(��� s��+�AK�!7�<L���4f�C$�R
�Kٷ$E-65�*���V��aֳ)Y��t��̩��8�q |���#Z�t�F '��|�Cv�P�i�e���ẻP���p|:v��鯔@�4	������B��S���\-N�8	��KL������b̩�BFS����	"��0���$B�-?)rK����7ӔN�����J����P�4)��~4ܿF�Ӊ<��_b��Z��r8�����KG�^9#Ш�}������mo���,ӽ��,�PQ�L>��6�ﵿ-�e~Mⴄ:��:izj���
�%���NՅ��4�Hi�U�N��9�%;}F3唎?�p|u������l��;���q�=��7Ⱥ����Dyw�<?�������F������x}:���s���}x�����z�}s�c�>"�&�ɽã?�}��.�^7����x�wa������w�}h�ͧ��+��8;<^�]��@��]������p�/�U�����O��??ޟ�}{�br�S���8�����~��}ڋ/�ջ6֕���~t�p�h��nz`� �xv{��F���{�|Yo�=�K���nݥ<����o�/���\|!�ۻ����'�����Kл�l�şB�}�+��A�%���d]�;�!G�)��v�)��ޓ�^��+�up�2AQ�қ?>J��^�{�i������Tn-z;s�!��{K��W4}��8����w���
oP($�& hFQ�C8"���T�hZ�ꦓ��K͈� d�p���t8,N:�5�z��q�ОF�&d��Ww(��Οi����hM�Xc�������}.Z�88����E��j&'�h�9�F�j�Li��>���P�7�:��L[rY��p��e{��:��\Sx�Ao*}�e��Qi��ޖ���B4&w�.*D���C��f�	��nN��Y�Vp�?�wW��0t��������o.���'��p\F,��9#&�գV!�>��;�\+�hF4�)���/tzqMp�Bp�X85�t�ֆ4�j�ͳU`�e5-g��Ւ���h�8.nݑՌ����H�a@d�b��t��*�v�ί�Uy�ܒ�#���VL�k�{Z�,Ԅ��N|8��(��Ȃ��4�;Sdx��r��DFä�7�D(��8��F�o�����1Ee9�H[ �͹��"�Q|�j�_6T�l�3�� ����)_�� F��8�ʅ�Y8f�!~�ŷ����
�-��*9��N�u�Ƒ[V�T�SȦ9�pGV�`�|����k7:dYo�C�~��.��G?j��P�y;�4~HX��5b:�DՉ>�A��J�jO�J�S�m�Q9;�GS������`4�QKF���H�4B�g餜��
��+*�#��G ���Tg�l�4@�9"�hm�(?�fB!�o�}Y8|֣[:�u�q��E!)��r�(i�����[�6��@Ĕ�Á;XIe�|
B�Y)�#�V�"=&q��������� �J�$պ$գ (Q-�|U�F�!v��1#���} �A�����.���B�I1�i�|Q�RVx[�{����$ܟ�hr�c����,FY������b߹Qb�)��-����8�2����O]B�����B��d#�I���G��Ԁ�T{|� 7r�uX!�j�m5�s[�9����[#'_	��2����|!
b-��r2 s��������@GA��
�:��v��C֝u�vWϾ�WB�T�E�`wUÏ��~��0�X�H` �6�g���g�θ^@kƌ���gg��w���ߢ�������fj���Bݫ�y�<͈��T{j�Ѓ�|���Ml�,&G
f[���8l]���,1|vXo�'�4&���~|S�|�-GԴQ._�%��L`�.� f�r�J1L%Z��V�֧<�����/�I�����NG�����m�Σ�zN��<$���@X%�I��l=�&4����S��.��ᰆi��C-�\'�M9Qgr� �E�́��+S���7�<U"ԉdAZ���1��t��*r��a�A9������!���m>� N-[�D ��Q��K�-��iʹ�����Yx�ʊi ��GK�\)m��|V(;�게h,�����:�k�D�|��d D@���(T��ώ��� �l۫��tJ��b���
�i̞ [B��㗕&�R� rx �=!�gg-J���y5�w�4#5Y��
�*�"�0�9M9u�1��lTh��p6�M9S��O�TrLH��E����T=`G'&0Z�]�I�U(���T�B�Q�U�����1%(�>+�#�G�x��h���X4#M?����
�.R����\>>0�8��M��m���p4`��L\h�JG�x����!�J�ꄃF���>"��D��Y���R��\�n�d����A�!`�.?R��T�@
~ĤӺ��4(�������E�%��n%Y�m>��R�I�r\g�FM�QK83�|vM�Y������z<�bK�Ӟ�Z;�3�,�**�&�R^}<V�f�t��;^�rEG9���EYG�����(ew��� � �n��1
�i$+�8����8��4r8��b�-�'�A�1dډ$�&�1%�1Ly҇,�ҥD5�:L$q�h&�f �V7�I����1�����O<鳽���7�ڄ*����L��9�Q��u�
���G>J��M���ub�>��'���2a���~x�R3���`��i��4����r֟�>��v}W�O�u_�#���!���?qp��f}Ѧ}��?9ڗ�rqwptx�L�)��i���o�/����>�{v���	n4��w|����ӳ���7��ҭH_�y{}��_�<\7Aώ���._�]��{ ԓ�����p^^����|T�>��[�����9��0nW�oͼ��~��{c��7,�r|��:������]�j�*,xt�L�h7o���n.=ٺ��=wgӽճ'�t;�woj�+�N�,\W�#{;>k��)�z�����_�(���$���<�1�Mp�k��[��!�71||�����~��GY�FѼ��jL��#�X8o�����,|o_{�_Ew/zk�)�����t�X��jXT��>�zf'�_b��N#�qm��h�l��9����@Vb�^'u"�]-��L.$0Y��#ņk8��d�B񭱽-��?���V�t����T����}�V��8�h�A8;/ʗ^�mL���u�aBM�b1C0M�G��MfYє�)G�8��pL���r�*�(�8�h��I!2"ф�OiY��r�m�~�G�7F0)�P4Q���#�ssg�,/Lo}{=�y듃PW8^�IA�(1м��5ޏ$�@QdL�
m�7��i���~�3)��������w7T��P�~��_�� סU8��kL�8DD9�b�g
^:Bjz�1LE_�v��U	�s�B6e]Ӫ"Q]U4fj	�W9%��S�c�6�&,����\Mˤ�W��e,��&��u��0\�V}��m�A)�9Z�%���cY�D��/K�M�ԕ(��YE���DF�"�����������}�_��_��#R��qZ�tC4�*��]0f�h�f$�P7�s��m�h>�(7�p�BKk[�nkxR�[�8^H@G����@���wn8Wz7���|D������t"Q]���[9QV��D9�4x��ꎚ��k��i�L;^�Z�������+��U"1˂OGH3�Sd��Pi�h��r~��s���T����!e��}K�dKD�L����k�F4�D�FNj� ���Qb�i��B�>�#�D�a!��jKf�֞��jiې(�SKҍ@LNd�́{u�^U�c��v�5L�Y��n�q1���V�.a��ŴUP��b��C�B8�XKC�)���v��&}!�/Yh��VJ"���^}8^�^��a?����!D�L�J1�S���1�O���w�}W�j��|V���8@:��B�Bh��؞K5���u�K��)Qh�^F(q>rNS�4���#�!�p�?�zs�� ���"Պ8_���$"�S:!��)��K��6�wp��(jZE>�ZL~
8��>2k*�V'�w�˲RѤ��H=WG��^,h~Kp<}�Z⋚:!��h>[�|[*+���U"�Q"�ڴ��Z/��g	N�ї%ZcE�%��J����r�1�����r�s�����T�9B%FY�P�)��A0��^(э�@+M�r#OW�w�%&�T��r;�vw>m#-�aSN�5���e�H��Knp*$w��^��B�hJ'K��ne�;�q����R�ʤL�r�؝�5�UTz)l	�d�� ��� >KS���5�s �(
1�pNYj�D#�чCR�e*��.��&��LŪL"B��2�j�����k���Y%�w��	q�̖V�Դ�'b�5E�-?�(q�S.�m�)�Y����Dv�c���������@�!D���Z�R�,�P�a
� ��:�C���V�'R:YSVbpv���!Y�)�&w�ɲ�0�r�_���ІCG"Z�-d�s�̗npb|^�@S�|LѺ5M��RXx���^W�-����џ�K��g�W��i�˩"Z�9�r"�'>R�1T�Ԁ#��(�C�&g�r0�U|���MY����A�����p��r������B8[��S�Y�PCcM�4	fM+">�eM�
��|��Xd�1�b�YLx����B�B@"�O�8�p6~���e�C4B���h�U�R�o�� ��gDR�U3�kq������Y͔�c���?�)�J�/Z�ffCH�:U���FC0%k::9>_J4��R�F��X�ʘ|���"L3�(�겊N�r�T]
�T�Th�Ʌ#�l����Cdô:���#B��9[�*d�L|!x��8�Y����l�#@��%��1�[���AdH�z;d�.ڢU���_hMk�pJ�5�9II�;�����%)��#Hǧ ĉ T4?)dCHz�$�XUR��U�d��F=@0�Z��0����Ȟ9<9���tQ׾��f������������;����s��x��@�����Bz|`�z=|i��Gǟ�D9���z����g�ޞM���{��wW�/��>=y���^\<{������������ˋS�z�hX�]��_�#O��������cᎤ;��z��N����=�U���>,����һ�.=>�v��K�w��[�k��n���*����GP��j�>���{��O_;�=��/=��x��#����V��:<�y��;�5=ʩ荀��\/�r�����۷�M݆#��;4�k*
7d�z@����w��?���Ty3��=z�~��m����vo�x�ǣ#6�����>ĒS����цw	zG�y�'�m%�������t�p �|b	�m)����͘t��,j���;�����ǁ?dQ2���]?�j�����In��)4S�$�R�7D���ɦ�̦�[�[�WJ@F3��n-m�� _�U��;�������Jaj��Tmr5-*%�]�j���Y�D<��Ac#.�M�ȣ1m9��"QYM9�ߨm�e!���a7Q�贜���K�O���%�4�Vs���*�����%Q����o���H�W��+�E��^��W�WYi��O��BK�	^榵�+�,q1q�Ӌ��Uſo�o��?���+�b�A@����
��6Ƅ��L��w�A:��׾<��&E�����UX���[���+��u'˭\O�[&.��lIu`ئ��X}��l4�����
�
�\!%XQjQ%Z<eSN�A350���U��t8e�/٦�p�Ja!J���2 ���&�Q������]�6��j@!��)6���5����d6��o՜�RT�7UTJ���K1�r�1ͱdRѤ����6D��I��Tg��/KA��q�hɖ�"Q�(Q
��T��\�h��B��^�R��)�6�Q�1!�q��K�iu�HC�tv�%�����JLe>Ш�Ș5/�i�Y)Ms��91�~p�q�g�4S�d;V'�z�4j�B�nQh|�t>���o�+1��.4Q[�4�B�4�VD�I��yN����/���/P�!@Co��p���Bm(T����TJ�l�~���{^���_ES�,� �py�^� -a��iX��M-ӎi礵C��(�L�P��\��&�,?�4_35І�iCHQ?).J~2)�'���[R~Q�(�T� ^�^�^�^�B�R4Y?`[��$"�m����� �񍤚�[u����[�lY�K���9�G@�	�$[ʮ_T�mA�K��'���,ў������^>�zs�M9���:D��8ǨQ|E�2�բ���|�To� �b�#���H�Qz�-B�����*'�,��@�FÊ�]�Y���4���'H��U����RsY�s�5_m;~SV!ѡ��@QSRj�KL*VE; �dK��$ȩ�~�p`�l!�H���(��HS��i��J2Q�Q��M���!������[�1��R�t������ w7���f=�儛�B�yĩn��ɚ�Z�Zz��!f)5fQS���^�����S��zC� ��c�쮑����³85:S7��E��ѧ�� �8�M�)��_T1E�U�(�1JW��r4|!�B!�Y�d9h��rU�YV|�B0i�PZ=p�c%F+Ddv.�U�-%¯DY��c`��#M�)�rp�h�!	S� ��^�)��P�v&��B�H��"��j5�����@�T.eQU*]����s~+��1(`�:�T���G-~Q �>��)߈Á�I*�D���5J���U���X`��)#g��� ����nZ��UD��U���ω�JIJ�V��R�#7��ҫ!e�>[)9�,>�p��J�e�r�*�Ek#<�M��-m)�iQR��I�NDMGj���p�)�o�6�8�#�lO���R����1DM��C#�S�-������Q� R��ܔ&>�S��Zcx����B����Eu�S������Pn�"kϧҪ    IDAT�y%�J7JķV	�ت@�\�i"�������DS��*��ۀe�SoJ�H���T���"�����*���h)�RH�D`�D~�#��m�|�6
-&����&�
o{¯�&�F)I�B��}/Xo�a���H�(+d� kB��F��7�'��=:R��]�S�(�5t��vNZ�)�_H-d~kg�L7�/�h�9u;�bvic=D囪5�MU����8�l�i;��B�[ �;E@���!~]�f�/�Ŵ8�tC���'+3Q�����	NSM�Q�^�:�!k:���Yc@4S�����e9p4'���1������8><rW�#�W�w�I��{~7���z]֮}T�r�mw%���?�uC��×Gn�����vN�\�^{�q��E��=���=Ľw2{��\�߸�x�w�r����7��{Gn%�ｼ���=���~)]_Vr|���ٰv|������~��_��/o�/}��Ozwp|�r~f�}���݉�4-�P-O�:���g��u}wsx|�r=����M�t��w|Z�G3ݯu�����͠�'{7/��]+��m�_?�h���X������qf;�+�:{�G���x������v=������74��8�F�i@����wBo�x;�G6����z7)���o{jӛ�R~�ӟ���?��*�:��P��Z!t����Ɨ�{�������Ս���ѹ������;{��'3y/��[o��������7�%���/���(d�\(K_{�8 +�x�o̵�N�p��<\���� ķ^�.Q��T!�?�8��%&,�4[9���YW��p���)7A
Ѫ�6�a�M��b5����F;���k ��gkx�|q�JG���J7�� �ڙJ�u�[n�[�T���8� 0)��1�D�d5 �\յ'9��FSeJԼPQ)BՂL.�?�)�����Y�,���m �>��*�'_T
����7M�J�9Bz�h�c+��>���'g����aׇ�ON�} �o�`�⺳�J�K�34{�x����o|������!������G[�w��	۾�XQW
�]y�{P���w��ρ���⒢�ۄ��o3-����2)d**��4�[T+]W��d� ��S��Tem���B�)���M�X�p�ts���sO���YD�����{���uC�Sͯ���R��-�5e�K�1��KD:k�b�eS}�^S3�0��iK�e*�J�����5�0E�A q`
��Cl��B�A6p0m����Җ��nZ�98B� �Ƭ���F�CE
|��"�Q֮���*Q�#������Q�a�@�Y�Z�L��`?z�8:�";&d�l}4��������s�0�mG8N�uv��'e��4���BhD���IJ"��+�3_h�%vn�|���N�T���A��QBH
fR�Q"
1�3J�ij��rp��!ā��pQ!)�-�2Ш����'&Z�H-q4�GH���	嘒�(>S����Ҟa�4��B�&1�"��p������S@3*�iu��([�_
hr��wy���-��c��X��E�����)5֠�J��i�8NN)B�3�%��U��3J!� �4e�����tAS�O��>�H	w��N]Ё>pտ�!��rӃ�T��� �o���԰M�_�ǿJa���[�i�-��h3M��Vk�V @�B,�H�I!B��!D��%˅ȒU7�R�p�L��l�]2%�f['j
씞� ��+jj�q��I'��
Y��5�C���D�
���:=$*�
�~djC��E�tŶ'����jC���[�K�Q���jC��9u�e�����Z��;P�Y>�3`���Z��־lG*��U�����P�Q�a{�l��ʄ�W�f�d�85�	Mc�#�/=�y��+���i�)��C
,�=���FKb�?>����M�}�K���D3ҁt� Q���C3�5��htr�ڟME�;7*�@��T�Nؑ�����-咍4�9�U�䠱k�l�{�ԛ<B�Ec�N��@?�'���_:�~8�\�.��p�j�����$:�j	^9SN��N<��s�C�P6���|8>Y����Ґ�A6����6��2�0m�v��c��A�����Zr���c��a���>�)�,>�T �@3�����m��z41�HE�g�!,�r�tY��v�g��͡4�g�F��t� ΖHJ4�uU�Tz���K!Z�Dx:���B@!�`����ƶ"?����J� ȂO.��BR�bEq8F��Xۈ_����k�CR�)�Y��F����d�
Ub,�DX r�r�M{�Ɯ*9��lu�lK �O���_�[����&�N�
%ϩ�!��($�h��t�8�g��>�i[)
!u�"UuvJ��7Z~��؄8,����ܮ����jIhV�_o�!��i��Be-��iS��ĥ���rf��P�Ȫ��o�Օ��ަ������Kc6M��WtlS����i�JBx= u�
��XC���L�J�M�[2����L�i!�,��C�EAd�kZ"�@Q�ő���5M�!Z	�8�gB6fN��m?�i��l�f!6ST�~M�rɲ�>)c6p*�κ�%�z�ćH1�h��`SұC3p��"�3'�h!�M|��N�i�_4�ĳE�JH�%r��c�<@N�X�.��}�vh�t�S!V��=g:�tj@?D.�t��-��"a�oќ��+a���V�7����/#B�=9���u��n�W?ޯ���FJ/+1�	OC�t�=M�!{�.�z�=O�,k�_Rc?��wP���+W�"<wDo�	��>��͙�<��'4�mBW���������'�����kA�Nt�wwr&�طWz��d�)������_�)q�F���m�xf˝ڻ��a!��GQݻu��=���~S�>&�]]Oj���==m�ո�Y��r�9{t��u��ή����O�}\�W������"�ݭ�u�n|�����ĺ�#�_�k��)�b�3ʁs��7%�m	���������ͻ:�����sk����#�K��/�_�{��{���y#�������{>X�7�����;�~~����9��|��'������m\�6?}�5����j�Z�D�}��΍u:<����2�8u�)�+ô�:@:|�KJ��Mearp�O"�(�/ʖ�3��"d!��)U&UtW�N^ɚ��4Ka_�agBխ�M�ܺ��vm A��O��mr�Ȼ��Yz{�O�_�4Fa`�V���z��y��82Ј?N�@�FY��R����h��(r�����<a�9hB����� ����ݪd!E9i�	����5#d���v�Ϧ)�A��x.K.�_~�-����~||�Bszvr������׾����7=z.��/}���W��?���o������Ԧ�9�������s���9��?x��K���������O�O�K�n�_����կ~�G�&=ɭmͫ���M;���ٖ���r��@3%k	�@`�D��B#M!�,S
�����C�9@j��������q�G�71=�n��R�<i9��!	�m��5�u&d��]���ވ��h����C��)ҁ#�,%0����5�l)r��|����>�J���D!o��5:,>��/j*$k��r��ݐi���d�|�i؜*¥�zN
Cj@��1k�/=�B��pc�����t���_���ijnj&އ5�~���zm�~�[��2sJ���<s^9=(���s����-�x�@\����s�TTnocI�om�{-�4Y�-
.=eSQ
�D��j�6փ�aLk��!�Ɵr���*ʒ�gVH
�c����T�v���(�4�0�d�Dt"˰!�h�]�8t�Ԥp,��Qi�5K��Q��*���b��;a4^E�ADMY!}�3�d�-�vd9V��7'$��mY�e�HQڈ��q0��A0�F����P�tD1���p�UE1�HbW[;\]�D�J�����d�+��q��
�G6�v������c��d%D]�k��_U�t�.�.�^�r��J՚�۫z`Mc�qfr��5�:��N�3)pC�|���$�*m�(k����cGM!S�@�y��c�5��"��0�9��!�*�o[���J�YѮZ)�Ch�:�P��� �@����2��9�ӎu�].p���HGz�C�u.�.��^���:q�V�U����ӤjU鲀L���@�ବ9�B�8���G�)��Z;�D#K��?�Y��LR�UL<r)��9%rJ�<VW#�Y���m�ObQ4�J��+4!L2NÕg:I��x�ǜ��BjBi�*���f�L�s�ig�D�?x͗H
mW����;�ʵ��QJ"+3?5u�U��$��7Jis�1�P
�ʑ�zn���d�U�7�a!�)ͧSt�6fN��du^q|at�awEBr���ϡ�����Y��� ��^z��Z����[|`��S65D;::�42��7�&ѐ�� -ĶL�pS��e��L�P d���hC(�'���SvF��X��hʦ|���-�>B6Ы�U7�^��b`�SKd�M��4&;�pY8,�L.ǨJ]�NYs�RJa#4���4��PFV�NVɭh!�C�P._�m���cW��J��Ț&����r���N_��+�a_��Hu�Zl#q�S��"�4%)D-k�M�D�PbX
�:鰁�+��x��J� �,�6�����f*]4�:*ۯyiN�RF�8NHj���K������b8!�\���3e���_H�~�wD�JD�88|!��1T�m��1�4U��l�4�*�єSB�r��8�HA�\'	�M�yzƧPQɲ�h5%U]�i/�@��v�?jBMY!2]U�%����8+m�*�O�#3٦�V����@���K�i�_o��}v�SN)�@�D�H�#B�Xs> ���s��",�6�ũ�Bh��r||��6X���[cqL�+є���#��l�r0e�e�K!�A�9Q��h�5��0�9����@���޴u�����c��C� �l��ٞ�	��bd4�Y0��t>����P��J��2��������P6��?��4;4���au����~rv�&D����'=�����������.��=ٸ�����_���OZ��sj4��!����__Ṏx�{����j^_��,ؽo%ؼ�B�s���ȳ��Ƨ�����{��j}�����O����O���y|�QG�{㇑f�i��P�rڬW�vM>:�M��fE������b�����yv��u7Y��O���ɻ�qzvf{׃�w{7�Wo�Y��L>]U_�yKsy�G�[��������s)�C`+��ɮv_�1_�mC��޷��82��?Ͻ���tUXO^zC�1ub#{�G.�/��/�����������MY|��~��>���l�W�y�������D훧O|?�[��k�n�<��������3MM���GOo��9���q���VRD΀�
�dS�R�%�3v�"��S���;x̦�����/qwZz��.k��	Ę���8�l����/qW6���dd�� �LJ����h8�3�]�?[3|�FU"�<[
����	5e��?b��|R8��ߊ�H4�n"�Q
�DN�:Ɋ|K�$�fT.;������Z�#Y/|j6��	V��m�Nx?e��\�]�ӓ�_;;=��&�uOx�����{��ޯ=9��gw�7/n\_;?;����|򇳳uq��o|㛞�\C�^���~�ۂ�O��}�w���w����������������/���>��Ckq�Ƴ���7�5�[��H�<�׹���
����
�^>���-�52ڨ�����R"pԅ��µ��O���5E��� }��"�����V]1m�4r�Y�eTF4G1�M���b��[@۱~<^;rgGp�r:��C�2�N=�Gh��Ѭ�D8h�aE�������-s�c�B��U�S�8�ZJAJ��٦�p-0MS��M���҅��49�,���ZF.��*��4�v�C�T��{�����1qM!g����֚"�(����.Y���E����/��[u���@:�N	Y8�)h��z�[Q�d|��j�F
��EYQVȨL�F
�\oIa��f��Z�(�x�je!v�e&[:k��XD��WȮ�h@]%����L��F��P̬P�4c��b��R��+�j.W?l�q�R�#�C�b��*������G.Y��N�e�5UWo
q�p�pV��燩��r�8�����ht��+-j�!�P6m�!���"I4b��p�B8�V�g���]�K�_S�j�+�ˊ��~��~��V���k��euY7ń�'����sm���+��O���#�t�X�\���[Qx�|"|�(e�WT�C�$r�K��r�1!u�t�%VZná�8�E��|+�^Gp`�Gۙ�GhEh�[���5�)�/���Xz%R� �'�ɚ����Yb7���:�R�7��Gf �Ւ�Ĺ�{BL��!�'�f@��F�����4�t��Ɓo�k�B�@(�	15��bB"����d`b9H�5F�)[�YW[�6�G0h"�����,_�*
W[۫F�f'eD�hp)@c�{��\gW��l��BK@��h��������2KKִM0���C�r����4~Rh5l:�D#�t�)���q���j[
r���b���%N��a�&N�f�ȵ�z1Z5D3�i,)�66�M!�V.��(1��S]"N��X�9�e��#�Bh�@��.SȀ�E���	��SR��w�MQ)�ȴfR��
��-Y�r�>Q)���6�P 5Y���S?@g�,�I�BuU΁pv�,Hmب|SU�/j����ubj�QH�cHI�4�F�'X98Đ�7�9��(�'aeE�Y>�B��8S�)�VQz��
��Ӱ��<JDN��Ld4#���i
��s�`�
��e�&k����R��E3�,*=?��1��G��7�jC�NFG�&�IqDᤜ�Ӣ"E�z�E��4es�1M9�|~m�YdNj��h��6 �-m�?$��/7N����Ѽ1�0�8�P��Ɨ%d ө�l���N*�����)N�l�rMk��	ʹMK��&UL9$��i9��L?�9�%�Z[Zz~��!�D�(�Q�\Q�� �5�z��.L�\�κ8���T:P����,]�^�^V�"א� 'b��R?OG����tR.DD��>����5p�ko4!����P�Wk!�l:�:׉tj���C�)� ������J�ßi�tQK������8����٨ _��o�v�y��*�K�&H���p[��$���nA������WnkI��%�A�"QJ�SE��,?�7��q��8�hsj���1+ͯ!5��򁺪���Q����ȭ�����\]�?�g�������Co��RH|�F���tV���������;��f,�n�I)n<ngξ[��X�^¾eR�ۭ��<������/,�d!�sd�{b�Tc��s�1�i�����|��=v�������I�(���7����_^]�x��j��;1�<v���/����ސ٢�K:�4u��N7Q�u��x��#�ہںZy��������%������wpz����M������L��G;^�xy{�.��9��0�X� y��Ǐ���X{/�.9RZ5:��K�������~��В�������}�T.k�q7�{�R��O��o��o���q+�w����Ϟ}�����'?���������?\|������S�%�=]O����������e�������׿��P-��H_-������<8!�iH�%�"e9:��k�=|T0�b�J	�D�p�7忢0��mz���1�rX�b��Sh#>�=B��L�`; K�;~��tr�O�X���*]z��YѺ���	�5
U"MxR���,�,Z~�r�$;�	%RW�J�b�;��X�h8��M�4)V7:p�hl�Ӊ/�9��9�6�N�©�R����F��G�E$҄�G�T���3f��e��/�u�/����׽N��)|��u�����o9޻������B�*    IDAT=��'7���G��u�ť�e����|������3������^{��MR��W�������g��v��O+��3)��xk�?��r�t��4�,���əe�[8P	��1m�9�x��$B�X:�~���!Պ&%A�p�X�G�����Gy��8�^���0�,���+�P�A[� �S��B���uO$��R���EiЁ#�����#(��P�sF���j�� W��R�)fn@�,���-���i��B�`�^���7��*�c*Z	S�����r	ⴜz0�,�5���uX��jaNhen=� �G��h~j��òm�߳b-9Q���� M֏[{�U��Е�����1�{0���3U����j�U�	��$���y%�C��yS!�ܖ�1�J�%�=lɲL�q�!�,)�l ����f�B�S?63�B��䷨�dM+��2�rs�tR���,��C���H�CYH:eQL�T{��fv9m{%
E���i���^D�фpDY�����5��ӕ,��t�W$�һ~�%!j�ďc��⋦<RdEr,���R��֏����,�!���*����%�m��nw{�IHg�L�D!/�*��\��{���?��Zm�Z�3���H�ۺz�9Ыɥ������Bp������PK�Ip�,Q4H�r DRfU� #�J`r�s�ʊ3H8! ~嚊&^"_�����(�������8��R�h�S=WDV� ���u�1�k����L��,
�rE9@�p)|QW�B��)�Q�*f�&�9f8O:����ZV��}�C�Ek �)AN[�)�i�B��%�nVHc�8���r��,gt���Om~�ӳ�����D�@N#Av��@Rt����R�h�����A�#8Y�x
�Q)	�2�G㓭D��B�C��h�E���'�UԒ�B�/��VC�Q��\9"Υ��Y
N+�B��m��(H}�����ֵ:�_]�|���!Ȋ �\4����C�e�EQ ��rLk����kXi�f���B��8^},0����t!���3 -G�>i*Q.�2�a���cԪ)�sL�qXm�ubO&�G�C���f:cD |)�0�6G��O!)�ڨ��2H�#SΩÐD
Ef�Y�����ޮSn�����l���r��ёn8L�-Gη���,�*YSd)�$A��1&�Q��P)������O�t��������#�Z�H�M3�Y�o�0���h�!U���a�� �P���V������5H�(~�8� BW���� �N�%brvk!t�8F�r�)��c��r��U��_Ӫo�u���k��!@��𢻾C��a
o+��'w����b���p�EI��8|#BR3�)QV�|8�*���O�ҵʗ��H�B@�������O���:+F�#%�d�m����i�*ꜟ�LK�C�q(4��D*'�
�N��oS8���u��z��l�T�,�rz�U�BugJG"~��8�~dF���r *֏�r��F�ҞpxՉ�R`%�p���*�	�n�*]Ho�-65�!
@2v�(P�����7ʢ)Zi
��|]�&���������BJG�l�J#�4PQ����#�ȩ�d!R���]��a� �l%��RJ��V��o�Y�!1'�T�6J�1)Z{���~���"C�Ձ�o�:�$+�)�����:���Dc����:��E}�(�`;�@��f���\�.�74��D�_���#Tmi��+���\1��pbx�F�-rOQ����{���e>�WESˮt���g�ݭ��>ч���2zX����ݬ�3}"�������p��W�>�������'������q��Z���1�,��VҾ�;x��X��;��:�}ުU�w{tr����wn|i�����������́����W���ɶ��K�����މ�K-�G��Q�A�(H;�خ�p|ߝ��(�Y�rz�HG��Vu��^n���?��N�Z]"��9��e공_o�������F>��
�����������o>q+�������{o�|zp���^{rzf7������ǧ'Ί��{�����>=<����~��+�}���ۯ+�c�k?mK�g�)�}ők��&H��V����2B4:rE�S!vD����nM��C���X
k wqH�d%"�\4NͰ�p@SL���1H�L���tv*V��c1-P{6�&!N���*�t�)#�&7�'���TY	��)�4GW�3%��D�Fk,k4D n*=$kZ	S='�,���ዲ�#�T���S��*S�f���G.ǀ��8S�o��	��R�b�}��htf��'����/�=��rׯ=9�9}��gOO����:;9~�?�8�o3���/�/Nn>������|�����z�G!W�'������ww_���������'�=�sy��?~����Z�M��<}퍽��5������}�0��P��'���:FT۽qa��b�3�bw�L�lG:�Ӑi����B���z�0ʝc���4��Cd��{���͊0������?	y�w���H�d�Y��^ G���hM9�őNG� ia�ulj4MA]���lm𭓔)2�2Y� ��I<2?���qXQG��p�M�cV��Qcn	 %�l�8h���(Pz̢Y
�[�����,!RB���7L��i��-k��E��eֆ3��[bR�F����q2ɕ��w���������C��4E&8-9�A�p�s��5�
9F,�*��R:
p-���"j�E��vh$��FRґ���� ҁL;t2E�F�cx]��]��z0z9�J��C\bj���m,��*��խ4�T �o���ֲ����"�
>D4e�]M:��qD�@��\��a�X5r�;��&I���	��s!Sj�h3����\\ ��rD	6���i6M<r�|�.��	Y��+��I�:P���Y�v����D0 p�S��i,��[KJ[�����J��+GD�?�>I����MӉ�.k��O�~ÿ$�����\{h�J`J\+�V/75=>;�q׏�B�4[���� "�Z29�R��Yc�kR��ܖ�1� ������G��
܀��d�X"@!ӪC� 2}��� &)`��A�wՐ��DK�,����l�NY�j�a-���|��
B��&� Wl'��ˁ��8,�����XN|4<kF�h�9h8��s��s��;�,ڠ�P
ARRZQ!S~-�8^V�I-}�1������ 3@̿3k��F��D�,��𐘥��0�h�"�HZ�Q�tʢ��mxu��j�TN�luQ�N`:�������y�"T�f��r�1L=���B"8pR����R����8	6e�#�W%��%:h�YS��@"lE�P�JlߴD'$�\G.k���q��D�%�c+g[] 2)�L���ԀĉV]���YbD��4� ��,���`1�`8E��."-q�ٜ8��礌#R]x�rӁ��������"cu�g����8r��p�R%"چT]�$&b�K���t���(�)Z	`��B8�)�`d�o���2m	����O��BI�Ou���P�(q>D��*�-T3#���8풓<�Γ5%ŏVzitt�f %�����t���oC��G
�;�R�Mi*��o(�6��u��'_.�-����Q�� B�#���JdI�c�`��~�㷴Q��+�_J�Q�(j �F�붆v�9uũ���+G�o����⳪��P̦��Q�)� ��)>��+�r� v}��'�5J䔋�RJQ���~M&�d�>�1=ˆ���x|QW�J	��o@8e!��ۢ��F+wB�S��|`�C�d�9�S?Y��JG�[iH+�Ȧ�iv�@RVԨ�t��ᥰ�Ғ�Q����nȒW>�hE7�2���(��֤�L�t�@ړ��� �"2[Z��t�t9�5�ӧ9��Y>��W��2ĺ��B6�?<B������~��P�
�[��m��D bD�!�S�B,|�fZE:�6SF�����L]�NL��y�7���U9Pz�,�� rjRY�Mf��G�C��C\����z�`BV���,�M�6����ԛ߷�H�}��W�]{r�j��H�������G��ݯ/l��OO�r��z��{,������u��� ��Y�V�CV=Fy����>i�EO�9S�7N:�>�u�XZ�+����������\��g'��ܻX�}�.�_u{����7���=��5q77�_�$�:��Ws�>�ՏO��ُ3��}߅��yG���+���g�����y��p�z�t������8۟-n�7�\�4z�+8ק�r��S��&��Qk�՞�̪�s}w�)��p�>;�lk;.|!�ڟ��o�y�;K|o9��6�x��h:4�qzO�w���g?�կ~�7�7��)J��IȞO���?����|�믟<��������Ӌu1;�\����ɓ�}�������O_\=qy�������f���>���_�;��r�v�u�!��r��C�O�Lj�]��:�_�RD��J��<4S+�o�!8��
������$B�M?9��6�-�T�n٦M[>�Y8_�f� �fU*�cfE9%��Ù�G�&���NJY��*���a��r-0�j�)�9r�Ю_4��(AL��5�#<��!Z
�	�z�eY~%" W���&�V�%"]JY��M������Rѕ�E�����~��P����|M����o|y����񍧾��铧ǧ7��b�|���ݥ�>�yv�G����.^z7�{�n��<mU4�:w~x|{q|���7��wuK�_��/?���'oy�����qޝ߹���hR���q�q��xS�K����`[4Ê�jm]L�[���gE���/���m�)�Va���n6�U��pa����5VH�
�������~7|?u�������N	��G�4�t Y��A݅�G�E3D-�#�S+��	�����de�p����A�l" �϶k��f�9#Z͈�B��i��SM���Y��de�a�eL`48��TD�;�p�]��#�1�[4�o�|���������@��,a�V����wA���y��sy���2�e[��-4���~�{���?�S���'?��B���w"���:aH�!R�@!-IWq����Wh�rKt�����e-A��Z��N`!C"C('>��Mw�M�TǑ�r��B��Y>\um#�u�R���C�ʵ:|�?��4O?_�r�dY~��k��i�D�jҺX�Cp�Tka���CJ��7xm�`N��L�8|�C��V�����
�K��Q���8�rMUA ��߉�z�Z�ZÔ#�N֏,���Ն,���V-���L���?��NP� ��κ��UN1�BB�S��|ϿC�vd�� �שZ�=�[Mnv��w����u}�`Z�"'�~���6-'}QN-��5E`��M!e�ɟä���m(���0��B����8�'�D};�4p]��7�2��d�Ί�3�:%��P� w'D��UX�rҫ+Kz�B�9�#��VݺL�JDs�V�85O�'>ܰp�T��4��OQ霆�NS�Y�3M��e��,����Rp$���6.K�&1	1m[�!��ISt+�
�)B��	���jR�Ch�I-��fS�J��!N�uU]�Tlӈԛ�p�w��ԕh���o{��t�]��qF�_�p�)\
>�i�^�&���#>��i�E�v@n�h3�y����B����ө��j��)dTWn��j�zf���_N�(k C���$'[��Y�d�$�n::0��ߕ�C
�;j����VV̚�`���i�Y{�����!�,��a��򷼕��?�&Y;���F~H�Bl�v�O�΍���;��W��t�@
�>��R�Z��{;4�̔��(�p��Df��z�!"Eh����G����SL ���,��r[ږ�pW���	d���� 3�'�ز>��?����B��ccM�#H������m7�V
��6�̖�B49p��R�im�$0��B�]Bۓ�5�T�Z#E9B�_9�#n>�t�Gy���BM�ҥ$2RUaQ�0m�)��ִm�X��y�O����N"�3�ii*�,G���h�������:NL4�OsK]2|���0&Zʦ����V���-��D��V�4�h��N6�B�ͧY	��H�$[���NQY����Rల^QN��J�O�%W�(�H��qj[!#N��
!�F�t ��N��Q�O�,-�)ӕP=���k���4�%S0%���Y��b�R�Z��қ��a�%�?�*@���V���1J*1��%w)$"wn��� Soʎ8��!��"G��0�h��
�E�Ϛ�H/E�@��qp"�4Z۴h)@GypS��+dD��T�@�ߚ�K�5��sYt*r��&#`
ufBpZ,Pi��5��jFV
49�Xk�V�E&�aGp�hU���T�f�k��~b�M�:�W"��_�.ڐ��#���o|����:?=}�(5������!�&�g�^��g!�ٝsiaۯ}��}{s�^�v��Vx�r=F�F�9�H�h��y��ۺ��zH���mR�m�׸n~��8X_���۝w'��W'>��^�]����T!�IO���\�z���M��Z:���+��w5��]N��<�/��}��q���{rt�]l��+����󓳫�볓�u����ʭ���u�n=��ً��7�����3��'n�^��S�����{3p���@ߑ2�wf��9pu��������燵cg��+ӏ?���q�����?��t_�� ��GG��3��������w޸;>���3�(i`���H��~~�ǗG�?9~r������>��Љ/�Ӭ�է�v��ol�ۉ7�ki8�~D"-��e��a�o��y�b86-'�][!�Tἂ��d#yK�ϖ��%Z���f�ʍ�/����k8�l�RۥهtD!Lgen��1�.S�J��$�t�Dv˕�D�&��үI!p��U�䳢�����Ʈh-lC��r�zk�p� >۔?�'�(ǔϡ�B~�%��c�@Z/�)�#�5�'�q!�V�K�뽃R�}/a7&���<����g��I���ON>�_:���d����-.��t��_�/�ܼ8������ͩ{S�y�͓��_X�]X�o������O���]�/>y~���ǿ��ˋ��������w|���o�RBo|Ħk�������+�?�+�x?��ږ��>�B��P�����>�GPԦ���cs�bR�x7ut�4uߗC
貉3�I�[��.�?���q�(=���o�*r�\�<�;M����%�VE���K�)�Ĩc����qX8eL>�-�l!�oa-�,nl�.#��J�
�$ER-N͘�s��A97��Hp3�+"�4��YS#�B�deqjG���'�^�%ˎ3��K�kfeU���P��ح�$��L�p���L��r �(k��$�F�p�;�*+�܏~k��8������?����;v���a%�c!���t_�h`�*� g|�JdMT����j,�)�����n��w hҩ���#��K��K�	[�7ٝ6���_��O�S{��x�ߑi�Ъ�Q�&�%�!�U�J����Oc�8�|:��a�fZ���m8c��IG�A�š)�CF������ �Z,_Vj��YE) �FS
�6�&N��8��(TnUچ�iU(�r�5��A0�z����48���1�� �,ʧ��(g�b�:����_opQn� ��5e�=���:�Jd!�@�8��Z���B��H�-g���5@�ݲ*��(>P��FSJ���-_�:!�c@,�|S
R�"���ܐ�f*ˡ)Z�-IZ��7��S��hH�.�7��Q��ȴDPz�p�����D�z-��ϙ"H75�峅*W�)-Z{�j�c�˭Dd����M]�X�,8�Nn��m� 5gK�C��8-P�~K@%�P9H�Pej�*��&�l����'g�h�k�N�U.�~XX�hi���)����z�8+\�Ein��W�z�khIuL�����MNB�����L*�F�Ϫ[)��&�����T"��W�����\��<[����9��ڎ3��<U���p���~�z��8�    IDAT�P~��h8�|N�*��T�@!#p��f��:)є�)�������7m	�JS+��bE�Ї+A3Y�Bt8B_(�#���#_H�-��g߯����FEY�J���d�%�myk��>�h���s:7�9�-g��h
�&�n� ��ֈ����Q�#%��B�N���%�[/��r�ր�٦Y�J,�5 �d��JkIÉ�&d*��([t_�_'�*��� �ȩa�΀|�&�C����-phқNS:�����:>N4Ru��>G�Tz�*�J����c,��cb�v�E�}͍���OqR�F��+�QW��!�H�(!�QH�|���7�n!Bȅʚ����sj��q�q�m��<��g]�X�:�ÁS�~�e�$�Ш%�)�%�uNo)S��}�B�sR6�@m��K��6ɷ��֎L�``��D�I���PӪ�J)1�Tb�i��r�	���1%�i9u5k��2BQRD9�չP �e҇ pJ�︘:C*���x-��RMK�:�O\n�Z�g4�Z2� ᳘��M9�#��"�D`m�4�Ȭ��(�"�BH��7E�4����~�8D6�:������\���d�4SE��Y
DbJ!�	1*�(+W�t#NY�ȕ�n�ip��$H���ހRL�819D�td��t��1u��Y|QHn ��i�_��78��LHQ
!��ٺJ�,)|~�چ�c��VW�:��gj��c�IVbZ�� ��Z�>s ���˅���d�T(��0��lN�R��)ë`�k�Y�DZ��G6GEQv�[q:B�� ��S�D����ZB�,~�pY5Yu�,�Jt)[{z�#�O��`
I4���l�G�mh!C�XM>���=�u��������x{�᫛�WW�o|���ƛb���k�l��7~�>n�^�Z�����e}��x�i���O|��]���=t_��p���G�:c�Q�B��|&�����@�ܣ?`郡���y�>�����M�����������e��������^����R�88Ҏ/���:�vn����=Ib:A�m�P}��ί{��`!B��6�ڷȮ�[�\wto�����������:����{�n���^�ޭ/�]���v钽�zsD���2�r"����k���1�M�f��X���'�����;�N/�}�Je�?{����>�5�����Z��>d�.�����_�����å��z�g�}��ųǻ㯿����~����՛+�^__�������/�~�����r�ֵ%�&���О�sM�L�~!���>�cjė��:3��/�ܬ��ȑ�`��I��n+!D���ɪV��':�h4��M�
��(�9y�DQ!�~�i��D��i��'�tf��#�$?ʡ5�x���e!ɚ�[��������( K��RuS])$e����<Qx��F��c
Eˏ)j��U̒�6[�]rO�"J��8��!�é4\o�h�<���'�!����{���s_:����ȃ��tw{��ɋ���w�/����J�[�}�ܿ�x8���g�ۗ7�7~�x=s�+�Ƽi��]��(�|�_�×_�����/^�D�=�N������߽�������g+��=�ǽ]��=�X�|�j��9�3m�,_�@~�����.�4)h�9�)�U�����bA��:��=J�)�q�K�+��ϸ��JeI�~����eD�ĿQ �E�)-���iG������4U�ŨWC�Y�4��ь`��xY@�2�����AL'������8�V��-��tͧ̇���b��@іO�2�%�)���)T-!�l�i�c�aR ��g�Ѷ�o/:�Z�'} �~{��Sh9,S���h>��IZ��q����[g�^��C
����/�'`��}�L���b��(Љ.���!�V�P��Q^�q4&J��H�LS�b��������+*�@��@ ���4�L1m&D�؊"�EY"�"*ȶR�)F�Nf4(��t~uM��$_4�>)L����P:_Q|��N�o:�S���-]K�Yu�$+ΚV�cP6UK?tL��Y�-
^p=k ���M�.�I�K��)��9�R���A._�"���T�JW!��8Uj�m�.��GV���z,
�bJY!=@��J1��N�R܏��P�RςN{E��e�����U�B��"x��Yj�W��k�E~6���<2��1���B�~.�)[�����%� �>+�rѭ�kJ��4J��@�:t��v��=q���0�&�[���	���∆����Xk�v�3���Ua�,�h�AH�p>�h���(��尐tRؗmEN�+d83�Ȭ�znX��\Sq��R���I8tp( ��Dò�-
i2f��h8K^�4[����������~t�)����9B��*��_Em�V�C��� �A���Y�é�i���1OA.��)��[Y!#���))4���gG��2{R?�;4%�s�קi�����u�uΖ�Z�jE
��?R���Ιl]B8mEj|�LY:���3����(~[��1
A�W�_J��[�T��[:���S4+�R���RVgO"�0Be!��EJ"d�X��|0mu���S�¡�>����NR��ʹ(Q��2m�|KLd�r���p#��zƙΩI���>Gz{B�id�? �[�j������o�AB�#�Q����X�@�	�ӔKA�a�s��)�1��M��'��=q����'�� ��c��?Z��R�p�Y��9
Ɋ ���n	Uo��eXW,��,��:ԀPL��I�%69٦��t�Brs��mHM�XQN��ި�ZJ��y�J���,�V��{@�Y�85 q-b�s��h�Z"����(�c�(*���>�K����~�RD-��!>GJ
,�N��� ��&f�8j���������r�%N��+J�0͏l�����Z)�� "j`6B��!r8B��ʙ��
hȂ(-��E�D�����k�ae��!��������[�Ryj���a��-��V"�TW�
|]�R�ٔi���ҁ�J�`Ia����Z�Rzb�ӷ	��jn!����'��O�a�88�ފXC�����*8)K�3:+��<����8��+�Yfz��p�"(���n�_.;)�t�>�8�%�#�Ϊ[�Z���KB�����^�b�m�+�T�6�Vd͔fU��;�E��c�٪Y�V�O�a5�$�OȯC6�-���t8��V�b4R�e9��pӓ�z���ŋ7����������_]��9>}|s}�p�jw'�'(�4w�xtwz�[?�yԯRz/�G3}��g�߻��]����ㇻ���Ǐ�n �?����L��}��o�<<=YO��7�Zދ�]>x��w����/u����n��>>\������ݙ#u�D>�y�m�������'W����o|k���n}VR�cj}Rt\_W������۲k|�ԟ�>�����・[C���no�<���B�}��뛫��s�.�߿򅼧�~��>����F=��~}�����k�k}q������::@��p�����ő���ut�.뀮�Oo�;�]����=
�0���� ��_��?}��o�S�����?��}���^~��˳��W_�.޿�e�g��y�w���8�����3o�޾>������ƭ��/?�_~�;�����:}b��>]�4ft.i���N<= �wk��Z&d��1� ��v�����T�(<���i�#���?Y���|6gKz��}P�"N!�R4��7N�4�-��K<ͱp~Q�� �9��m�Ѐ�.��j�辝B��鼔��4�J �b+*d�M�:�/7$r�����dU��EcAs����`���C���R�Ȫ�WOYJ8N ��D�N��v
6>;�ZW
C�3��>���ٛ�������q����7Ǉ�����;�.������؛�~��|���=ڝ�s����m��ݞ\߬훼}dݿq�]�������99�|wzvt���~��n�}����_�����{���z/���_��?����l����[<�vvr��.zzn4���)��E�~��R�V����$(djL����4@�Ao��{/H��3Y��{���VWX��-P�w��C�A%�CK�z��P*|S5pj=&дv���|!�H45�CdU���a�"���8J�E4o����d�*NY�d�7"�4SL!w�]䓬V�������'�NG
�BƤ��Ӏ��=���A؀��m�S��acr
�W�?�~��v��Shi5A�ɯ�Ԛ�"��v��;c�r�<��OK���t�W����qFcNDg�� ��B��VͩR�VBT��늂���Sn��"ˇ��x:3���&�8����Q��G[*ۙ����V!
ZB���� C"4�|�\�B����a!�̦6_��P}
��Q��W(N���� �XQ8ٴ��F�N���^T#��F˯�ZiCL�`�8��̀��@Y��ޡwF�v,�[��,Zõ�ﴬ%�N��g�=����4C�=!�nLIUS
�����Ml-③U�Zm\.�6,M>)��q8@w4�#�d�"GA�\���jj�ib�?�����e=B���,%�F��E�s�`�& c�r�8MYS�i��@mN�R��ǌS)�!�fV�gqE����r�l��60<a�@)@
�84�7��;D���+"@~�6;\{��[2���,
�b-f�!j���
q m�h
@uYڹO!fK�A��檽�r��ZB�
���Sv�Pv�v���*a�9vG��Vj
4zI�cHO_"�fH��i�����3d�<]�D锞ZHYB��8|h���`Zϭ���f�!� 8��đ��')c|
��B����m�,¦��/����P�#ۺ�<�W]���->ǀLNk�58YȨ�z0U+Z�C0��!Z*O�R����:D���9u�:�[)B�%H9u#�����T������v��N����厂��R!!���lp
�C�A0�)xx� 4Ŝ��D�&�i4�ƴM��`j��"T���O:5�$Ή��gK�����\�S��I���re��4�]�08xkh�oLi�$�Z��~��<�H�|!�)Z-���D�C�8���r*���-�]e������4�9U�U��k��Rl�*Yj5��i��78��r�j�������kT(�o��~�V�M"�J��*%|4�������O�e�rU'E6q>d�C��,�S�Lj�FH�"~Y,����ࣵ	�4��A�)=�� ~�@N%Bp���Ee!��s��P;	7�>m#�[T��4�"�2}>N8+�)|����	�b@�'[t����S��2)YhG�d�OSC
��#s��	�dVc�mg|O�$~ʦ����J���|���.S��:��I�!�u[(q���D
�W�5F�X.+W"K���l"l�PՑ��d�(\t��J�z[��(�Dj�+�F+jJb:m�R�:a�ʢB����>Y�DGy࠱t8��Z��CM�)?2;���Ș56x���|�ƈ�Li
�QZ!k�G(K(hE��0e���V�O�E�_]Q�E�pf�B���>�&h�ί�X�
I7�6�eRhZz�����|�r1�p�)���ۇ����� �5RplQ�)đ4Jw��V���z6m��
�H��Ug��@#�������Z0$rjpmY\����R��^�%H���თ�/^<���u��	��Bt��[�|���1���~��?޽��GW~���ᝓݹ�I���_��ݫ��ǳ�;?v�bfzvr��pws�݌���>n�w4�P�Oj�����V䓑G�x�;>=9\�:o�����7/N/����ן��8=�^OnnC��إ���;tC��2=iW��[�G�Uޜ����
�L[aؓN�i��N'��w���G�E�#uxs��x�^"=��&ܫ�7}����Ob�?����=|����ٺg�ͫ�ã3���{�#��z}8�"�i�W<שhɪr�ZN>��1M����Z���&�ᩜ��;����˥����?��K��	����͛�|�����;��'�~&����>zjq�����ѻ�>?<��|�����?��'��v���;�_����IVKN-(����ڙ�)�_�)k�,�(�	�.J�-ʟ(N��G�6Ti�*'q�D�����P#}�(��EY���������Xu ����Z~S���Jd=���}��V�+|��{N���	�u�"����<�i�*� �fgfRBuKJ�8Q9��ϴ�MY�)�5M<�B�\9*��T�cl:RM�؉T	j����i"�Զ�L9�F��*$���H7Ȋ�/�[�p�G|#��vG��^��/n�=ϮϘ���;�..����ş��Z�����Ŀ� xzt}t���׾��ۇ��Ww���]��?R||����w���������냛/_�|����bw�������/�������15����ɧ;O��{���m�>6�)�y�·"#'�����LV�/�,�D8qV����e���{瓬�ڨ|4dY���M^��Џ�T�F����-�V,�Pƭ>��;Ő
������@��$�r���$R��k�XB� �F�ᗒ��2��U��ˇ�i@���qo麵�7�7�W���A�V)��r�Z�gZ�I{�YMY~����@͇W��æ\9ӐJ�)�Ț��)��o�;����N�v�������Ȕ�4pS��L%,��GY��	n����N�-�w��rUT���B�s6�rB�"]"�V�r�M���,[��J���y
�
����N �Chsp���R����=��lQ�I��Ԥ�K7�+WQV3Uǩ�,4:�����,���� �J��#���r�(g�a�q��R��M!�s��t�z�R�B�D��Hw��Yǚ��2�B�.Un��8�D�h��5텍�C"G�u�_�N�YG'�bI��hN9jB�7&�,�����P
@����||�XWاW�pߐ��,��6<R\�}lN�F[Ym��0�/~���ك��&�\�B�Vq0u����v��P'�\H�+]�=���OL:�idNCh
����
R,q
�ag�q�Ɓg��� ��G��`�r�gd�TH_W
ڃ��BFdn��֎����������P����'�r��!�D�wXE��%�Ck�4|LCu�)�l�lt��U��"+m�镕,���ťp��ԛ��&�gSx���ѳ�S#�dC�L��ƴ�a80r���[�21��ii�Y�2��Y8�[�OW]�+1�?YGJ��-jR8�p�`@ʶ��ob:Y5"EFY�ՊS���������6d�l -�&��ƚ�bV��1d��MMTn}BHMn�hlmp��T��J���1�xO״:aq�=� ��8�A�l�d5��[�����s��D4d��	��J�8N�9��#���d�
%>{4z.�֠�a뜠�-�~���q����G��!�*D�����tS�`єY�1�0�V{p��6"�u�W�5FY��1�D�X�%��d�8D�1��uЁ�@0B�TJ�Y��8����JRi�~!v�W���K��G���1�/j���U�5_�rM9[񵽩�JGT��@z�M!飜f:p�0)$�"T�)�����O6���V��Z�(X���'�фT����?�(���y��OS�&���!�G!>G��Z�4��d��A0
��!N8�tXc֙fJ?Ax��!e��d���P:~��s�r�0����T��h�}����#�b��g�('�r�OttҜ�ԕU`��QH9!H�>B��B�BP����>r�r�#��Z�MG���Q�D���F)|�,#N ��4Gi��u5�Ꮒ�T�sSj�?�R�Vt,Bkt��aDp�;Qqd�F�/��r���!_���F)B��+1-+�LQ3�� �i����O75�+����!�i!�B��p��g1��̖�~�ZJ�Y�{��O�`[WK|!VMk��Bʬ�ZSN��T��)d���h��Ln���_���Q���	'嵶�7��%��˗yŢ���    IDAT��q$�5��E
Ĵ��TQ�;���B|C�i��R�	U%~�0�e�eᳳ�xYh�Kt�� �I����ZN/�v���T���3��zx��×�w0ܨT�}Ɲ�~���z�7�u������z�{�C��z{�C�6�>�]�Z{|r��N�������z�s��jף���|�¦������M�۟�y��=�7
>�ܝ{����>�X��7/��o���n�?���֏Xz9�n+y�;r���������˚'�'�#S��l��`3�N�:8�^�MV�I�^�0�;5K����V���L���\}��x룗|�ߌ�@�����~��ۗW��~Q�������Fo4�jד��Q�H�����uȠ�qg�3
n��������s�Ä�I��rm��MTjo�}}�����/�?�g��6w����~r�g��������������g�����������)]����_|����۫��ɢ��������^ߢ�֠����6d�۵jo9��SM�;	[B���4#|���8!jEK'ej�{�7�[L��8E1S��)0�-�R��B���������l�|�S�,���䓒%���E�9�8�@6��,���x6}�\$��L	�Q
��4�~Ӷ=�>����!𤄀'0PzQ�(�VVm�Ŋʒ>4:�jC�5�l�rٜIWT�[����Hv Y���B�BE��q�w�@Q��15~ �*�����#������؛���g|�X�68=>:q��.�G�'�~^�`w���?
�N.N�\\����z���>���~��%���~�������>���|����J?�Uկ�>���?{����~i���̿YqsT3w7��������3�Y�V��Y��v�Ŋ�*$Ők��c��r9Bl'-�4�X��$z�R�h��Np|	���Ղx#�E���v�e��v�2z����m+�F�S%D����|x)�|G��l�j�S
�eG���p� ����L�d�_�H��8�"G�7 Bƴa���_�f6�Zf�c�*rR�҅�e�<p�mNs�ԕ��oS(�,`�ܩ�4��B|����Kg���ћ��
8Q�V�aqǎ�3�������6�5�0�_��q�RS�I��t"z��^�p>B�*$R�klhHT-�F;��NG����"D��s"�^�B���|��a�Ǉ�QW�Q(�e)p쉵H����m�'5��i ��Q�B�
�����4�
�k;Y8�7H��$��+7�,=�&.��6ZQ:8����Bp>˧���-�B�LT�.P�(~'ǔ/��[����ąA"�u�;��R� M�Y2�ג%p4�ϙ�$"K����/����	�h����$R� � �W&~�Y�][m��vӓ��>��-^4���4VES85�ւé%�*z3mTT"����HW�|[�T�;�L
-�D4;>f"��i�����+Ѯ��Z�'?ߤj�|YB�X��y��vpI5 U7�N��U��'=�@��nIU]Hz��f�9��T�A�a��:��w���%�J6\��4�NB���+!�(AL��kM� ��i�)d��(��\MQ�3-����ZEj�Bე�eM�N<�pQ���iY?l[$A����9��i�=�����������h���m#�k��"���-��ߔֆ�#$�C��ٓ���<&X-4�%(�6Q�(q��t���\]S��(K��"�Q
�4�$���x��O8f"��,��(���!��ȭ���+R"�|�i*�P�� �i��huK�k)GJm��`"��C"(��Wk��u��|�:ٔV�S"~=C�F�8iN.)�@QL>�0�Fg4�Z��F+��Cf*!/D��1>D���6��Z}Nc�3���Q��Ǭ�P-%n{1G
ؐ��Gs�*4=T"�5ů4Kaz�K�0M1gc�BJ�[��IxmH�G��2HJ��2M���%&��IV�8��!?�ي@�F��j����L�~�,1Q��=ͰE��F���9U����S:B�=��S�~B�t��B�5%$����r F!
E��Á�"�@S�Qu��U\�[";Y��C�E��M�e��Su�K���)W������?*Dh!%F���>�ސ1�D�d�46�b��]I7�ഐ��L���<��D)�,�,>'Y �� �΅pZu~���Js֋��!WwD p�E.ߨb����8��N�X�ڋ���tLV�54S?9c�K�I���L%0ٲ�DVSZ��S���WQh�y*$D|h%6嫒?몄�z0E@��ɇ�fg��JO:h`��	�1���39����h��\�����=��"b���u��E�����e�qTii��6�a��J��l>ٜh�!����{���%�J��,��t� r���cP��68�D�|!#Gn�C����B��)�)���J���7!"���ȶjBk��� �Ѽ ��+�rw	[���>��%S���������f<��E�<�y|x��[�Q�G��Û��������ޝZ��͝o3�z��Ŭ�1~������k��#F�c�ނ�pu������7����~�����xvvyvr���G�7o��}�8?�ەޮs��������)ٍ�u���j���k[ց�N��O�����ޯǂ���j����}X?%z�,]�]�NYo�_�p굛��Dʇ�A��ۇ���훫�~}�굼�kK�rr
�w�׎?����{�|@���Ά:�z��6To;誃գ�����r�\�k�:eYt�N�ޅ������%M人�y��W_���o��o���/sx��?_��!G~����������������Q�1��>>�;?�����������Z�.���b���=��p��C���sd{�f���QO� N�)��Sd=�dџ�MY��9B�
E�(��c�%�5�|���7~�����V��q��R�|��*�'-�A��
�&����74�rj;��4M�G����:'�rL�q�3U�'��tJ���󤚲m�͔�H"3�J����E��Y|!`�f�,<?�QCkWsa5��DcSx!R'���V"��D"4���9���>�~������w����P����ݞ�N]L�nn����vtv���Eŝ���k��N�w�vG���;����7�~P�o#��<�}W��~�����|����Gǟ\^�����u���ٳ�/��|��}��ʁ<�K�%��_�.G�bXu+��P;� *@տ�:��d����B�!R�ā�b����t�:���h��"�]������Ʀ/�#KJt�5�u5���wK�B�������"Z���#���ɏ�A�<.�Os_y@4)���(�9�my�j,A��2��G`�C�nX��2D�򨿖�B�#
��*))tɯ~s���*7�Ŕآ88JL{[��c�-�,)�44ݯR4=�D��m�'EA��ο��֌*���&�6�w��L¤�/���"���M!��<I[�u|j�ݷ�U�ƈ#T����M� Bɲ�U����u8�D'��PW.|
qZf�Z��[��W�q�h�)��S-|L�	Si��V�5EHYT�0���7M��%�~6����,�n;�R4cu�|�i�9Y�Z�)�����4���8��M��t�Ȣ�E9���"'X�/�(���rL�ju��L��$:��^4)@�D�օ)�դg��z���KT��T��,N���%�N�Zտ6�� R(W�O��P�.�i�G�J�����X)��i�D)=$=*�+%
�
qȺ����?[�)�NX��'�B��m�|�#�` i������C���'δWh�"G�B���%�Ҷ��}/_K���=ށ��H9����4�ڨ7�[��}S�Hա)���i� ��A�8�(�/d81�-��n�o�ir$Utn�-y��wFՕ,����ҷi��9)�th4%�� �2����
Ro@�k,�P�G$����i��C2'k���
-W�B�k���,B����#��prN�|"pE�@��ߔm��d0���H6�d��E�d��!��*��ڥA8S��j	3�N���B��i�>�ԪbL`���lRgc��	B��ќ�M5!��L��"���-�i<��\�h� )��I�8� �#h (�r����E�CڷȅB0k���IQ>M>���#M�P�NM"@p#9�$
�V'��얽�,���D[f�%R����!T�tS�S�|
�C�V�*�	�Jg�qD5C3�NK���gK���O���-
g25bcj��_J S�����iY.kt����JL��!�[�'/ ���:�4P���*d�FDZJ������U�RVɧVMC�<lY�����խ���z�G������=`-�$�kE�Y/~Kȉ̗�,�HY|�����/�,��7���W��:E��,�&�>�F��#T���DC�(��&���� �b"�-��)��=!`u��߄�4�j��u�/n����R8E�R8���6j�T4�|:��tZ�Jд��Cˬ"\�����Aj�B|�� )��I�9@��ꐖY�PӤXL��A{b�>Y�攫zRC��%�s�&S�Í��m�t�D��Oߠ1E6e)L4�h:||8'5>�(�B��ъ�2
��ö���1�ĄHD���8%��Mbѭ��c	��#*T�@�`����0̩��,�M��D�RH�m�Z"d)hL��9��U��PS����O��p�]�Z�h���)7����v����M~�h�`*7_-��{B���h#_�t��Y�19���r|=��̝�ҍ)G$>�1����%�Wk���8�j�m+���p�@�ȵ-W"q`��������)�SJd4�Jd��[�(h,���T\Tܺ���m�w��2{p��<���������
=^?>xS����>�xt��C�v>ߝ����{�ǻ��{���n�^��g�zo�=I_7볏�'>�4}ϭ/u}p��T]���{������x�����߷��Jou����յ6�f�%�!L��^_y�;Z�9�}J]�[�jz;,�^m�s�BV�s�MH�]wM_��o�zs�ȝ���n��;]�짏i������[7loo�O�l�y���������nw�����F���֞ެ*k�r^鄲���*����;Z�3� �h��E�w|R�������G�Vu�����͕��|��~�&/��������{��=����Ώ��Cw�6�O��|��t�m��K�����i9oύ��f�:�r�j����L��1����'Z>B"�Bl~:|k!kD���Ζ�g�.�1����<[?�`r�rC�cQ[�49G��l:�!�?�����Gg��b��̔��IU.)��,4�ࢅZ�R����Y���*�e!#�ꬩA��Ds���*]9SL%┕���:/���R���--3�D����2��mсW���b���o-��Eu���������z:=�=���	�7�o�OΟ��_}�������g���o�>�����>��W�o�Ȧ����n_}�w}s��+�C�_<#�֊��]7X�=;�������;��7�>�޿��_�����o��~���/��^�#������vB���]G~�î��v��Z]�ձfEq����R�L"p�~�$��ku��w��6�k��LM�3�˿�K��{㻿���wKZ������׊cC��C���>�M]ykb�Ŗ�Z�N�8Nߠ`
D�NQk�T�p�������N
�4S%��� �v�>|�����RK@̶�Hn�w���k�rY�,��+]]�YN"qX82���*TWq �l�8�i�t�3B��s��yS?>a�q�X������˿��V}J̞tS�z��?(m�Etz���a�O��:�>���p��2��C�C���@����eJ�@Ç������.A���BD#�4���]BR"�m5ڀm;�V���(��㫎�)����1�%�Z·��toF�=��#�B3�/��:�R�B�l	qd�9r>#2�ů�))HS��cJ)ZJdG�1��dS4�hF"�b�zts�]�ʟ}�J���kg,����J�4���ӏ�6X���,���h�r��TN�)�fp���NV��J
A��!���b�ɺd{���d�\u{|�?��0�ȦIQn��.��t��i=>5Y����	�.Ӛ�y!#'pld���8ì
\Jd�����/%e|��9��O���:�3N���?��ϝ*��0�	=dJ7��R�Ug���̚�0&\���X�n��(d�4��,n �)�i�h�|�Z�|����Ai M�� ٺ�h98-f��"
�4��R�'�-u�"�UjF���0���6�p�뼽ČS'8�B�5\"|�P��f��PTz[���x�B8��J�$%Ě�!��7��	%2R���L!�Z�D^����~��&����gY��D>p�<=�!KJ��Y����1b�;��6�r����H�)Q-ʫ�mi]l���h�H��	�7�����1��'Ro�B�ԛt��V���1�9D��Q�h=�s8Ւb-� �M�Lۢ�LsRЕ3�Bj@䲢�1�d�3I�DL�@b���lo�WRU��ۙ���T�VL�jE�U%�d!8D&EY�J��7�M�B��l�Ɂ1�H3~�U�O�2��	I�U!~C{eېYd{�i��N�}�V:=ԕ��8;GVn�=[AJI?����� �^{d�Y��=�5i��\�p��j����لѤ d@��g�ل8�+��i�_��[?(t�)X)S3M8�2� �8��+~�*d-h*Ř=�Sk-e���O�$.�MQ~Y��h�5fj �Iɢ���`հ��OĨ+��X��\V�L�@gQ|)�,:�ƾ��3ZM�V��t�Ǐ�3�@)�R�9E�^��I��B�D����@�~8�!1n���Bee�)K�Ӄ�Ot��rSCh�55ڜ�B�mQS#�pS�Z�vj�Xj����Zg�������9MS=X)�I6�lY��\{���r9����*��p���6+���Bb��EI�����U"����l"���rLe�S�@X��%*Mbʉ�9S�Q!`�,��(�I��N�d�R߾8���I͊Lq�v΍R
�i8F{ȩU�4�r�du
囶
N�t�D�MӉY3����M�P[!"k�!!4!#}�(Oy~����ެ�)�\p���R��J��T���t��*
%��^�9Jt�h��7�a�V�B���F�(NH?P9+�x�J���t�Mt�������榠�{d<��aI�|�5��;i}���b�]1�}��?jys�7'W���H��n]�;�>�y�Υ���mXN��\7}T�Oa^�������{8�ӝ7ol������3�/_�v��3�!}*�_rޏ�w#s}5���������;�υ�7+�Щ�w�d�ֵƧ��9���E+w䷮wo0�{��IT���;�Ϟ�>{v�>�����+�dgs��tw���=�-���ۭ��:�,����ҷ������ѕO�>�n}]��-�u֡�_/������xQ���ޗp�y�\�w������Н)���F�����<x�?�����O��/�<y����_��%��/�O/|e�-�㠫�G�Zywq~p|�L������?��L'���5磝�l��Э�+��|���tf��[��u!{�S@�&DM>�J�$R���v��!�\?�@��&|r�S�����:��KW�'Zȿ��/�#>w�FsRԭ\<3��p@Rp�ɂ(g��s8L��-=�4eY�S��M���4���Q���ï4NN��!���6LNj!�@K?>�tc�8��j�H�~lW|4R�l|���UL'�iH�+�r�'"�e�z��������F�}<�hy�;�zs����3߰z�����������})������N\�.�_~v{���������ן�w��~y{��b�����o2ܼ�ދ���\߿����ū/�z���ٿ;>�ձ/�~����󋯾y�����_�+��Ȧw��i�c��b�8���J[r;c�ldm��_�@�aR�	8��K��h�JT�[�q�    IDAT��ߗ���)�,�
�L����=	y�s9��m}��?��?B�G@dN+u�RtmŰ��`�ӓ(QC�����*!H8�r�|�8�ZO�NX���C��\6�*�!5��
��4��/a�9i*j�.��9�jyg���> 8�tX��`��F]��qZ~+��z��ΒM^��B|�
�6�P"d-a�:/�d+b���$���o�[K�!�  I9����n8�<bm5�><�������BJ�F�����
�V[Q;�Q�,�[Z+j9���6Rô@��1[E�w|kL!鬔�"�e	��m�áf$3_uCV�(�Ȣ��o
4����9[{UK��&��	�+�ɶ
Ȑ9~6�Os��n��cJ�q���0k�����҄p�f4�ue]ש�tSʢ
U���'�]2�`8�0�.p���O�Bp$"C8��ɇ�*[J�~��(�A ���|��.��*�>kU"u��B�-�'?�ɏ�c�!
�rjƗ�|��H^�$[K�ci���|�K��}*'qNx����!>�@0T�nj��̏fZVVQ��5P��,J��pB��s�FNRE���eYKjC��jk���1�9h.ku�_�rZ&A~j5f��H�i��c�Ҵ��49F�%��2��NB�Nx�a����W"A���v����S���n��&p��v���ɷ�|:��c�o�������y�a�R3M�(��M+�P�i�i4����!(�����W�=�4�ȅ�"���NB�eE7ֺ ��(��B6p�!�)Z�)f���)��6��f`j���e���X�ۣ&a%o餤��cқ��@��B�&ďIȯ
�,~�:I�k�e���hpC�)��䚆����|�f�өIR��CZ�!�@~Ky�,�Tz4!-!7�.k]���/f�E8>��lB�L[5Y��9�|��YK��BЈ��/K��
��t��*=AYd�S�!h��R���MS�ߡLPT���i�d�1|QM4�lY@��Ձ��O'�dq��� J\���r��?��2L�*rTI*;!��=�A/Q��@0��J	�)>��@���0AI�lM�)) ?�Uf�jvRrؘ�Zm�����A_z���y8����6/}
�I`4~�I1�!��`�B�ju�R��Z؜�mE��"��*��_4�$^��hJP�����D�I�}&_��7<�x\s���r���z�w&Db���|�dY2��J�|����t���2��8�tS�KI!���6��%泆�t͋	�9͏��C~%o#��Ɏ�HO�u���ϑՎ��s�i�(�:��MV���/��<���t�#W��"@�D8�TQ`�BJ�OB"����N�u�P"kt L�;��BST(?� �J����+mJA�m!����C*�\"��"�1����fY�k��ǀ��g�R@7%>��C�R�1��5S��B��)e����L�_��m&Ш.��:��!��J�'�r8���re�GE>���ɭ\d�P�H)]z�&Y��6��l�rk	��Y�1�hk\_����{�Kң��i輢�B$[p-��ܴ!�PW`�V��5���$Q��Z��"@֔�CNjl���I��:q�z�U4/֒�
���!7���D���K6_���pU�;�~ӝ�ſ���M_I�xv|�[}���l�����n�U�~���Z�[�G땯�QΩ�+jow�'W�W~O��&�#mw@�[Z��ܽE?c3�O.^]ݸ�y��ZS�'=���C�����G5��O�/�:X�'G�����O}Q��Ai�m�#Ȯ}���{���Ͻ�_д��������S_�b�����#������܍�{�얡�l��[����ė��J�����������o��=|�~���<���~�s=<;d:� u�\{�zx~����J��O>��|g���]����������Ey��2������|���?��G?z���g��w�_���=~x~p|��{$xg��p]�םׇ�lՎ��H'��V��MY-���q4��
G
XԔ�F �)!�u�7Bv�ކr�Pj�p#2�D�U�(oi��&��*�R�(�����D��bZ	v���h�����C �m�[Ǩ��!^c�E�5���B~S�hZ���Q-4��PQ�S�HR8FmL����GKD-L>0$�D�@���i��	���IL-��8j�0�tN[1|ө��м,|��$�Gzv)>bd�Ui�
�6UF��aj�g]���Cm��������Y���&~\������'�]~}�^����^�~	�����wn�^��lwy�|wr��O>�S��=���G]������{|��~�����ݫ��w����w����ͯ?���|~{wyz�����/�����W��].;��'.8�Q��v�c�B-���֘���d�O�p�4ᶥ�߶��%[D��
-��B�rIDnj'U�$��nQyo���{�����G?� s$_i�4D�a��TE��PG�0��|���@ �)�a�tzi���sp���qYh} ���zE!5��?���5�VK�C��G�ė���X0c��xU��F:|��"��i"��?'�b&��sY�)N�i�d��&�1m����@�Ii�Y�q��c��p�yMg)/��R��C`��R�H �m75��mj`�r���J�V�<�#+1[ͷj�8�iMۓ6g�D3�#�R��V�i
lGX4��(�A��� _J��.h9V�$4�4���a-��~�q��JA{Jz�����ȏL�(�vO:R��DD1�`�|%�r(@�8,���	a�p:+d��Ŏx4L�5:%:��h��*�:�z`�L�U� �U��(j����V�r��gk�&�qRB�PmH�Ǆ�"7�M�v�04&%)Q�dYUjRJ�h��{o�����3����w.�����ܐ�e�7�{H
����"w4?��Cj�	�J��v]i�#m:�oure��
��V�ա�ʕ�l��ԶmKY�m�E�L{BӴrSـ��[JY|�)
4�ɮ`�l�5z���Oj�~��_���'�6Mr���O���%h b@D�� BR�D B��l˴�*j&Z�����~ ��L>B)���P8D��Ȯ)�Օ\|�>~Ru�Ig�3\c5I��6���km�&�/�L��_�p�p���f����j?��DL�:5���9�7�9 WQN��_�T�U�:�B��S�,�i�h%�m,\�c�R��ɂ4�Ɂ�h��mQ%X���q�g� ��sYj�RuEьz���l��M�\8Ā�t6GWJs䶄e	%(j�e�4���S�T4��*�`}�Zʉ�ֈ��M%���7ͱ{UZ�=;�G3�(��J#8��m�\��#
A`"�ʚ��A���2�_i�ɣ�z��[r�BjUtN����A�պ6��/DSK����1��Z�'�5�(��a��u¦_�ӡ�ْ�N颪�4 '�m[ 8�C�RKh!�L9Fm�r�j*�N�#@�h8�-hj�7-A����v@3p~�8S�U��,��z8��=8}�Y!�QV"�{k����b��u�,B +����.��&�J�Ĉ��|-�_�,g�b�!K��,N8'r46Z͛��mΌ�%"%[eA,62�GzH4�A���A4E�rBr��ׇ�K �\#q>Pz+���$Dz��98���8uI�Ov�tV��&D"� Ӊ	l��8G(�,ô��a�6�>qBd�V�6�p�N�ӧ�[&q'�L��
! ���jI��XͰ���rq��5(I��麷ɮ���uͪ��I]��ecÆ��7U�y��a��C�X�Hk$Q�ȾT�}~����ij&@l�^�bE�}N����'3�jE�pꧢ�eQ0
� e�!�(ʁH�Qzߟ�t�����,V����Vm|H֊�9���00��1�!��OS-.��!�k"�c����b�����T�����@��6e�DJL��i4#��Ј�j��)R�?S�R*-JMV;�(��$r�%���|x�d'�Z��uR�|),�?�麄4Rn��,|%��A����"x1z] Q� ��@U�"��H�sb������?N�_i�(+3A���z�*� aҍ���/��G����rݒE��t[��*�2~��`Z�(�����S�l���p�	��B���MF�H?;��j��7��M3�����t���{�w'G'�����;"{������_D�5�F�λ[�S�3h��5k����g��x��ލ3A�﯏�ҽ?uԢ����[��>����_����ά��LN�����������8=�p{��?��u���C��nͮ�^G�M���s�}�u�цxy��g�ڄ�ɺ_{��Ao�O������'��n��w�\)���G��NvW��W×o_=�\y�����<��n�sd{��^K�u�QN3F�t�4�4��w���`o��,��sd�P��{�h˷�?���A���sz�k�����ջK?R�����җ�gO��u��wj�ԝ _ ������[m^knЮGA�����������am�SH���%8�'C���y�F��Y:�0�$b�-ӑ�G4f�Qw{!đ%�����-��G`���q*�N;PsR���˟_�z�mƯ��!���'ȟC(��߯��V9�F�P'A'[�L��Vb_�/=~�BH�����_.�)�d�a�e��RR]8��i���JG3f�	��?=�P�D�6����ǩDc���w+W�Z�������EW�ۻ�7�._�z�f=9�e�z����_�^�<�8=_�u������������������o~���o�z{�5�����;߼�;q�ӧd;�nDx�ܕ�O���g��ώ��OO�(���}������ݯ?��/����G_�γ��玏f���'H�h��e�i-�v�4N��L)B~T!��
q�vI�(Ǐ�-����FxdL[$�~LM
�V�����k��݂2'����=M˓�����5Mט.��L9���"�8t&]9>ė;)��>�8��΀ڶ0��Cd�/�,���������w�&�HY|L�Rh�|Ȓx�FD��EY)8_i`��Ә��l,e�&�VQ��|^H�m������P]~j�
��-u�}��ǵqC�n��'^	�/����.mM7�1�ӟ:�%����(�7ٕk�����F�r�%�a8|j��SJmǔ�٩����Lb:8q�6�c�Տ�T�ئ!p��G_J�p>�ȥ#�Z�t�%�<�1���u5H��A��C��BF=@�+�7e��98���-�6V��m�Z����L�!�ѡP]�	�w��K3l�x|�Դ�-��DRC��;W����jO�bu���/�DW�tj���)K�u�O�_]���C�^m�"z�/�ψȕ��4~���t�͞X�4B)^�R|�35��ܑ��g;�!��{x8�D�X#Yˁ�h��s@��qZ;����V��!j�ӑkji
aS�O9�-�B�	�iđ��xa4MDT3��A�c��p�������n���R'%J4Z�Q!"m�*�(
����/Z�@4c8)SN
�Z�Ze����ݰ���T45�v�ȯt)��툨(dt�r,�vu�␒��r��B��"�C8��Z�MǧТp(�^�M�mӲ���=�˲"|S#���!��3!�ea2zuX��� GW�j�r�4�o-
1���;
á �/MbQY%�=H�u����S!�Q�&B�@���y�,����p
	r��0 B �ϩ!)��h8~m���\~YI�I?��h��T�#�X���l4m2M�!�+�#ZiS�/�T.�Ӊ��Č��ٙ�D�,�~f!@�'�H�%�����B�*y�2&A�VHY�g:琝)&�I�DSY�7f�a"�c�V(qQN
��	�DF<����#N�U4҉�,?��� ���*�$�^YD� �2&G(�y�#�S{��s�&�F$��E��@��yeT%�Qi#~�Q�@DSNj���s��,��_M�eq�� f��;d�T4͏`TZ�����D �N��B�
�{EL�J�Ψb���N�~JQԨ�f88�C�S#ۏ6��W�5�˟�CЀr�lJ�vH������G���8-��)Y#���`:;��f�_B�_��T�5��<���BSnȐMY8���o�
5bJ�3]��^��@~���\"e���	b��;�:�0)�iO:d��,�Ƈ[_EcK�	$ȡ`䇯�6M|H)7)Ӛq�F�h��2-$�8�gB����^���h)P��ҥp�틻&8��.xm̨1"�6B�&4; ]��zP�%K�^�E�*�O�@��&����!Mө
�3�NL��I+-}�ejck&�(}�F02�d�+���=�d�NX�b�#X{q꧔�2�o�[1d�(A6�T�W���0���0��`B�����p��*��SE�l2���2�n�U�8���ve)�PN��Ȫ��9A��,�fXP�i�F��s�h_�H��`����n����I%Z�Fx�Z����ͅ3J"{�Q�w�ƞg1}���1�!��n��<����NI���ѭی떧g%W��H��zMޭ��o��O�՞/o���Uw���k�6������'9��~>���TO�y;ݍ��+�y{}{��u����c��'��y|�qʇg���}��o=�{�?{r�������ҿ�Z �_Gm[ѵ��K�;�޺w���O��{���[�N��SZ^�|ps����\_~qxu|�p�p�M �[_^��'gO.��>xzr��w~Cxwr}xpzr|�-_�����݁gI���n�׉���T/G����y��� ���v4�YǴwlD!�s��%vr��	q����x����K�����^��<;۽}�������G>����=�S����$�i�nt�^��޼�m��'Oz�p=�ppz�ت�۟��:�,�iC��N<��1-�;�脨�ѿ��\�I�'�䖞#�a|��P��̇7b�zu�Y!Φ�D��h�t�1ggZT�q����L�բ��a	6��~"���?��c{mZ|#�ʍ����~�0[HH����D����a�)�ØcmT�6�U�1֘��j�1Y`�Ƭ�8�C��@*-kz���%�B��KD0J�e���o�gH>rR�@)9p��r|�,�5����8��~��A�+�_��{�������孏�]\��5�����/��=�����W�>|�gԭ�����Ӌn>�>;�}����Ӌ'��'ͮo:���E˖qzt�|}�[����~
�y��Ogs�}���j}�u�"��l߻����A�@	1���mo�P�EV[��4�Ӿ�I?�]�>�PE�hF�njz?����@L�G)<���>����������?����Cj�]]TPF+��>�z�4S�-{�-�4B[�Dfڪ�e3�F�BdVbL���o𝂦J%���� �����Q�_o|V�@�au8Y�#d�Dj�(3�6�$b�F#2�U�4�[E|`�r�p갺R$��z&.�X��5��d�e()��|��o'�����Э��N	S�t�9L�v�u�Ӌ��3O
'��ձ���B�9��T���l�U��&�t�:.|�Iĩ��
!Ǝ�D~b4�!4M�(CN������YV���)Y�:�o;��HcKr�[�0����!�Q���f+22R24�Y�?/Ѫ�?r:!��!�D�СS�TLf'�)ǔ�M�&KY�Z�[/5|8D.��1��"=\c[�5@j�I��!Ms(t�������+a��������嵣��~��BA��删�R��m:F�	vP���N�"�V�N�QV�O�C�M9���~����C_�1<dM&�S㠕/T"���!bsL5��t�ũ
�O~�g��ڄFu����Y�Ω�i�>ʵQ:q4jp�4NVcFS8����4f�8�g8�B�76�k�%���9����c�m��
|�R8�:�**+)��t��h0��5�Ԁ�Ԉ� ɪ��ހr���I�S��Rr��c�BRX4N�i�n��<��Z#<B�3�1+�I���N>���)���	<����l��VaRHٱ|S6>M�Ζz0���q��5ԧ����KH���|:FQ�)�    IDAT��ȋ�ᓅ�hY�Ȝ�A���?R���8�B�.��Fw�Y �
�pz�d�r�p#��ǩ`��z�Ȉk;��F|�'B��br�nRU�3�19�65�*���i&�V(��ƯJөgU\}��g
d������O"ZS#5%����/$�8g6^n� @ҡ���,�IE�\3�	4�:�j�kR�4X���F��\]��O� '�x�F�&���Z��(��@��G�(��4B'R����4Y��������FY�@MWm�h=�(�Y���3�6�i��{������5B�4� �I<&'�I�)����˗��m�+�0�~����SV��K�i� `��%��D��Dc��E�1`�F�u^���5�d k	J�2N|N%h�	J,"��I�(Đ�F��iR4�B� �)�ȯV4S4%V��xSmO��2+7�A!N��̔q����䐥OM�N�F|�@�=Y�I�A6�G��h^��e5%.
Ꮓ��\�NLcu��z�dh1��)��S?�Ym��FM.�u��O�r���\Q&_�z(ŔS?p>��Ǉ�D&� mVjZo�Jp�A9}YU�[��LR�p����M��,Wh���0+Zo�v���Y�i�	��J�lL�)�rF�4�*�N�4+���՘��Q4���K���1!���j��NR�8�19�a�Dt��3LN��1��N��p2���_�F�攖�}'���?gdQ� 4)�dEÍ�5����D0��7�J��(qGh�+Y3��N�U����y�8ᦌ��QTc�̔B����A���6�O���ğ|~��A��'���k7}\��\-�/\��G��1u��Kz$ӫf��?���w,w��	վ-�;?�٬�_�i��u��������$c-���j_�$�֝����iM_���m�u�li�栏�������y,���G�܁t��?�V��z�>���o�5�v�<�r+��Wdn���*�~*٢�i���9ݔ=9����έ��I����v{8��ӣ7��ʉ�SqO�^�����ٱo��O�z�g::��ww��O.��H�ؾ�	�!k\K{��r� ޑ���d��]��
ny��}��au<y�M�'�R����?����G�x~�}��k޺�q~��w��G�JZ/v���C�Ʃ��O����i�QΝ8�]m���PzcA�~�N�f��Va�oʄ�·�<_I�F��'�\�~d>'B��%��( � |����i��G�3�&8~�E�ea�օ	��Yj|Q������Vb?}��B�3~�J@8��-���Vm�$M8�P(�q{ɯįHM�QL�--?} �a�7�L~�$���M�h�����Kĉf��q�74�r���8]]���l
R8�B�����	�\�rMW��B𣁹'��>޵��]{����v�zw��������e��l�h��_�~sz�������������y}�������_<���\�W��O?��Gͮ\���_��'�޽�|�������7��|�������_����e�^e�q���+��X�%0�+�E�*j����[>����6
��b�I����naB�h#Ad>P94W�DL}�;MB�G� �H_Ot���dMBҜ:2��|��
:`!h��*)�鼁� '1�\�@�a��:���Es&�F!�� �2)8�tU�R�۵���V�v_A"�~8��u%�Ȧ�h���7�c�h���R�6�FUrZ��9�#+���8x�8m����!�m�F[A�b7�'��tƻ���x����B�SK���o�VE��_��?��?��C��տfd5%H�����!�#C�)�bB%R�T9�JP��=';�|���rLE[o�
���l�M��p�&[�Fʢ��4��i|�����c��#%B�C|R�G�4D�@~P���U��*��hR0!�M��V��R��2S㦷R����">c�Mr]7�&�p��?B|���	�S!����;���N�5S�F8��C�@N>�8R h���t*
o�v�>���V�_34YνN?x
BYU��pRV*$˫ɷ/xqi��>%��u+������p�g>�c��Q`�}��P�K	��3���9��D
�3L�CT�8�QH-�1�/$%�����!�K�-?>qBZ2�I�G�_��nÍ.GpN[!E��Z�\���l��U|�
�E�����pDC�L9���M�E�ј1�90� L���dUE�@YM9�֛�T!euΜ��E��dY��1��Ʃ����`���L65��B���g�f�,��HaD��)��r,���j��VaN�j�M�P�CZ�6���4uI�d��\>Y`�Wt8�\�)�)M�_�2&Au��t��CY)�y]T���O�2�1eUR�D6�WB���c[~�ۢ5?�D�ǏP.8r��Ac��8Uo,Ec��qL�pҁ�E'>�Q������4>pB��]1�z��L�q���H� _��%(Ą��B6�ǣ�Í�@�!��c"a^��E+4:�K�1~m�,'Dʈ��k�y�ְ�$)W�,��b�0g#��aR���4j��a�D!e)�U[��:B�s�B��R�	�^�غ8�N�U���Q4�i�Ӟ(5�v�*��RK<������ZZ�ʚ1M���OG?A]�k!R�-P:�E�o��|�6��)~G�6�ɲd��z×�1�i�Qz��pHm�,'�pjm�E�0�᷇�ۓ)Q��,��snLzRM��Ԙ�Om��o[pjl?e�GZ�Lj�����P�Jm�9E)�KT��"��Ԣ�L�dY�QJ�h�9����(#nJ����-?H����95)��p&]�Q�T��k�4���45��s�_ȕ_��E�9�>�U��#ȡl��m�[����T+Z)F:�S���oZ����Z�wjd�GNH|%��h��!Bu�д�|"�*f|!"B��NH� ����?-qF��9GP���>K��i�ɯJ��6!q���aD �m�_*C�۶q�K4v��S���B�m�+����P?g����� ���.�_4 �T�0u���j�vUQ��������X�B�l����z84��i�T���[SRY��z0ʪ�B5	gV'Ki����ӆ�+���c����o�zF��G��t��6����z�r}a��R{����=>ߔ�������|��0�',�a�9��;Z7,Uױ�������lۿZr�҇�>x!K�u��|88YDρZ�;��{9�.=.yr{x��$�O�]7Wo�}t�W��z� G@����������w��p=��z�;2Ow\��0�o�B]�~�ϧԮ?����%�~ͻ[�]}����ݯ�q��c�$[�ۺ_�[��p����߅�}>O��^�a{�l�^�m��˃#���?JvW�����/;���O<�4V��Z�~1�vh�+�^9vp��D�wS9N`���h�rdG�GWz�A�跾�ͳ���~�˛׷?x��ס��x��71����ެ;�?���3���?��N�<��w2�]]�-�S��w��;�4�����,j]���sZWv"���(��7RnGF�45�ahƲ�@�6�JJS��z�H��I���O�Q���9����nT����'5Y#%���(�?����9�c��!;��8r#p���h&���d1�!�?S���JO*\�T�"�@QH8?B%�"������m�B�1�	��3��I
�F����VdʐG���BpNJ4��M���nޅ�̉�Oܐ{������0W뒷������~w7��]�(���7��Z�ٳ��L��٧����ٻ�sWb�X���z����u����3j{����?����O���G�����7���\��>�Q�O�ޟ]�k�7K�vqSS�*�9��O�F��j���������,�/�M��P"@%D�:@�6���4沩%ߡ��Mw0=��B�'�'�Ո�M'�$��v��uZ�)�"�z�')JbJA�@�\�i*���	�_!�Ęq$���������2>Dz��7����A*
�SH6��O����ܶ�cʩJ���&��p>�hY|N��oT�/g��3F3�mK
v>��ar���&[�1�!V��L1�8���Ҝ1~��s�hJ�0�՛Uk�i��^N;�Rz��5�O�r�D8�J���S�1�hq��>��Z2�[۔W��q�1��dIgBp%X�^A4���C���*m΢n=�$kd�O\:��E���� Q�B`�
aB�iOp���r��p>K9��QB���3���5̥��Џ�CG.GQ`���p�[pS�r(w:�J��d�.{N_n��&��F�p�ܓ"G�Q�,Qj�N$�3��^+BM�1S��Ls+�x�� �u��m���N�"�5��^d���!�5�ߜ~���w�̟���np"c���=��7`�m(HDP��3U�]�90U��%L�՞Q.C� ����R��(�dxf9�|�c�j>�JA���tS�6&��*ͯ
f�t�.Jr�1��9N�m��N�%��0eN:��H-NQL���J�o�Ip�nd@�ߨ=�d�' �D���Z
B�� >���ƱX�@��\"�w��-��" )�Nt���f��mN��1N�G&�)�嘶��$�Z�ւ���\gEӇ�t%�_�d��! ��چ���r���R�8S�Ƅ_�#To��3dv�Ҕ���3"h�Ɋ�45�A�8p��(MF�4�/K���H�%��*�v����Wb�4�(Z
�N-�u�7���S�RuS � D�|���R3���k� �6��P�gR0�2M�4�r#_4�(}~v��D.s�qF�X?�5Uo����v�V��픥�NJ]�DQ|Y��0mמ�F��v� �1���rjq2�:�3)����{�c*���F&���h�oDc|Qc���߆���J�N*G���è�m��Vm�+�8�>�4$��:4M|�:��y�,�V%���V8SL�,)��#�l�F`�)d�h�Go�+kN3x����RsIy!Y{�r��W�5��IA��[�jҺ��ܦS4M�D �ڦ�Hy��x��U��r&��dV�t��U4���I���fj5���:ߔ2dp���3���Ji*��f��B�3�UϘ8��f8�X������VcJD&ՈS�,���y_�q�MiJ�?��єU%~M���8!_
�����U�D�������Bm�%p��7V-�j5V��\n��pTd��?�,��h"��k�I���ؾ�vN�|�DL��BM[#?N]��W雲�o��Ve�B�ڐ;gv���#-B��m��p�CJi�e�ukL\4B�9S%���bJ�)����\e�v��� g7�{�E��hč����V:N48��Z�i[�I�KϏI�q��d�՘�F
�ig����
���0�U���Ҧ�MG��9�	\9?�e1~M�&�ԛ�,x���ȶ?�4DD׳#{o:��L�NNH�8�/Z�Ap4fT����3��i=�{*=�����]��߽W9AK�u��Ӎ>��|����]������'�� �[��ޞ��D�=8��]�����]_�i��^�wS�=������wnt:S�ܗ�qW�^����co�Լz�~�98�;��̗�>�w��к�y�6����n���P[a�����]�*�~�==_�Q��~rws��䕲� �c�l��|w� �<�sX}�-=O���Y�����	���Ovuj���b������yGYHi��Y�m{n�������n��:��x�k"�Gp�;��a=�?~���o?�pw��������ל�{�����c�>�qw�ч/֣���}e��z�v}�Zk����d�2�v���h�j�o]ڶ���n�"�^�)2�tV�{�Ф���B������MeiRK(��'�0j�UA��6��O7)4�Vi��~u��t2m��3Ng�Z���Q�T�*3���V�f��}e �I!�1eQ�ڣ	l,+��W�&�L�)���9h� 3k	����s0��N
ÜM�)��4�����;��-�/*A��iG�3F�TS�
q�g��SN�܎��L�����o����W�,\=��^�����O��'��}G�o%������O~��ӟ\������2펟>;�<�O���=X����vT{�a���c��~�i����0�������~���חoO��������G�g�Y�u�?���h���l-�oԞ]���vY��j�����+�Z>��HA
���F\�K�����%r$q\	ME���jԀ��p�^�-���X߷m�t �V\%��d2qj��t�`�
�2L�Wљ�p������"D��}��,�j�#JM���k�lǗ^c��4�r���!{�j�,d�a"�SCNh�w��𫛟�Q�hl�J@�D�FG�A�I���-��'����?q�
MϜ��.��IR�=|���K����^��t��
t3�;t�����Nd�G��~��ÿ�o�g�R�nO8��hj�M!u%KKRǱ(S��dqz��1�(p�A�XE��LgJT�Ȥ�9s vO.��$�ht86�稕�~����+�H�Z`
|Y�M�X�Dд��q@5���'U:2Ӽ�jՆ)<Y�D))K���Ǐç�i���!�AT�cƶT"�G�(��	A��%�_���?~EP���0/�ړ�i�Z#_�.�+�q"	1���?�u՛�EE0�(��5�H�@PT�~�yY�ۙ^_=�������)��>5u�O��R��?�c�(S4SR-J
G:�>E!,5c)#B;�瘶m��8]AD����2x��4�T�B1��a�9B8�@��!�����W�W�-M���]��O��9AD�B�(ӪD��t��n�|�ϡ!��0�X�M��Ԓ.���'�l��9Y�V#K�O鲐�c�eg�\�,��ӫ�C�M3ҥh���p�bx��e!G�7�jj4�CD�iT�Z@6>GѦȲ(� ç���D�9���C�_Q��H�1Q��Y4&�cd�z㘖ŉI�+N)�z@f8,�:Kj�����b#۔`�TV`)���3"�}d"�t8�\NL�)�L
&�V�8��c��8I!���yK�����JW�OD��D~���1g��G�T4���)���2�iYE�h �,��>�D4V�)���ztі�CRl?�,d�	M�|!)49���ug�ɧ_��S�P.�ɩ:��p��*�&e��H���B�ZӘ�?P��*K�Zp�8���4CR�l!�ന�Fʪ����Ȋ���5��֔_�J���/=���s(�(�L�����h��Ư�8�Jр\̦�$e*%x��[�
�B����R �DN��M?��t�D��H}�r�-a?��
��������*�(4���O
���Q�m��L(N=@LY��o�k�J��1�f |Y�~����įf�)ǔa���VZ���!��=�p8�&���d���hm�1�
U1���ȁ7M�T�h��U"�����\��ьSem��"H���W�ub*ʟ)q7�b�2�3]qD��s)ӀPY�K�cJ�!~:h8���h�شDS��D��R3��8rd�1�)�t���fXёMG:3�*���V���7��H���z����F���D��(�A1�۪�L����z��戦S��e�gj
�	O$f-�
���h�9�-��dE��S GݜY�J�CAd��͙�/��)8F�p��~9 �2�n��N����S�q�_��V��m�4�cm{�TS���.�֒Ecr4�I#N���ug9R"�28AY!�����5�Yim%2:��H��Ĥc���iK&("��є���@|��'"OO�|��w��I��3�M��@P?kl�í�bԙ�������b�l?w�э����	�3�(z��SEG~�w�r���^`nAz ��܏��#u�}�G7ן�n���4u�I�z��h�~��/����,�oK}v�	%�uu{u�>��(��2ϊn���Z������~��0o�����w|v~q�Yեs���Z9뭹��_C�H�N=j����̝�=��N���PY{�n=�j�j�9��ng�mN0s    IDAT�8����u�բl��w�C��{�w
�V��S[p]U�QnU�u�j��0���1"l����׿������{�N�������c[�Ϟ?{�r�#�g�xs������=�=�W���� ��Y����v�=\��SU�e���\�G\њot^��p���3�
��!��2��N
��W-ܔx&�.�T!SN!4ۢXŜ�G���Z�c]��_!�6L���dSTzd��f
�z�VQ-�����>�QS�X���}�()����(�r�L��jL�+ʟ1L4F��[Kx�D7�##P���g@F*��Z�OW�˙B�|#A䎋���!J�H�D:e� �Ah�JR�~�B�BM��糥�g���
����=���]1�j�Ǉ�=�Klg���n�ZK=|�ū׿���orz����ݹo)�OP��x{twu����������Ӗ�o�W
�ޞ��=d]���p���w�w����'����?=�]\|����}����g7?�����.Nw�^�eX�Y[a�v�2K�[E[a��6�ɏ0&ɏ@Y:?��hm�����Ւ�|��a
?�я�r;���}̡���N��.WR��.�bpi�4��HPl���SV�J�4"�� ,�S��Q��������F�gQu�0s��������p����ۆ
YK��c5�hRX?{�hR7�I���T_Wp� ����Ŵ�r���hI���5���sP"#P+2`~Y�8��,�8:���(�� �,ө����1"xW��5����=`dY��?��?�p����O>�D-��p��n���v�A)�k�`�I9�Y#�r�h?�q 0�D��lW�B�-�(ʊr�_	�Lu}48��D#(W���0VNna�p:�B@jS�%kN����
�t�W���b:UpX��h8J�˵�|4}2L��p8R�脈��#���B�5f��N`R�����,#s>8�栔ҿ�0*�g���VQceVH�M#��(]�z�!���I=�p��)��q�tt��bZ)ߨ�&�?P�e���R������[��n�j��RD����1~}�9)E9E�B� �/R.����0RB|�B���̆M�A�T�N�U}���
�`��6pխ���&+����cs:���Ԓ6hJ�iK����Bd~���zk���0٤s&d��9���R������F8�t��h�:d�k;�lj�$ő��r.�[KvS�>!~�^���B�������!Ӑ�h�kZKF��1�!p���gQ�pE9Ekl�	'"��Z�)�ij���k(W"N>�BuXH.Gn��%˩%�h�9dU�c	��D�S�1�
\��BFH�8J�Գi����94���&�c�q&70'pμ4ҙ�ì+���Kt��~����,BH!���_��"�;-�,�Ѵu�T"�_zR�c�
�6]���1V�XzS�ML�u�2#Ь�D>B�����,�(@L[,�f� �Ə�A6f�J2���FS�)��+�\(�h�pƗn,͔����q�;����eD�01JO�&�HG0�rG�mx����,�ԎIgu�#K��6-Ĉ�0�5-�/���)B�|N��}�\4c_-
�
i�"�����F[T�v�O
d
Sє�2�|#�Q�[2�t8
A$V�_!N=�;�1Q�(T�C��Fu�§mH� ���b���~�*@V�Ѵ�MuU{��q$B(�6���1���VK�C��Y��#D�D��)�&���:�>j�9!d�D�E�l���HɊ*Q�i�9��-V���K1��g/���L	 �4�w���[�D���Á��U�ӕ�|���
�b�ԝ�q�p��^D�K�N��̴�Dk�[H�(�I�#j!�	����=��?�l���G�x=�M�4�����UB�f~��?YZ"6����A��9Lb)V]id8��F�q��B����l:��B�RK�<|`��ą8�4�>���1$�)���׌	�ol:j��@��qWi�">�y��B������g�ZBh������Rh��B���p{>�fN���!�}6�?��?�P��IN�Ԉo�^;��8?��j�4'2��tR.�ަ�Ŀ�*����ҍ�$���R_���5L�sYp�?���g)
�V-A���zT������n���馞��z���܉��n����C�z��Ν0-��(������|�샇5��@�ۇN��MJ�{���<�����.��pO����m�[�hz�p������㣋����wneJu���YG�ėf��[_VqycJ��nO�[�v��$��d=�n)�[���s=bypu{�;�)��+��o}��׋�ﶓ�I��]�����m�n��ڹ��$��c�������=��.��[;�{:={w�҇���bG���ʼCet��P��2�::���8'X'���ρ~{3S-�q���]nߣyp���Kk�I��ۍի����7w'>Dw��F}���|{}�;8?�Y���<����>����n+r)x��f���*i�C\{��1�[����gC���rG�8���M���8B��~�H�ՆiH�淥_�F���d_�|��dF#���� �+��Z�N)�J'��81'$������0�l��~n���U9�~Q��Ve��l�� �������q��[��������d�3zE�8@j�d���Uh@�چ����+���)8���&p|Y)O�C�(T?������nT�����j�E�'����!bc�5�7�|���s����O����E�_�f͇ݻ�w�_�\<�۹�yx���Ĕ�������@mp/�uY���я~�F|���o8���������͛߬g�o��c��'��{�hҥ�}ki!h6�h]l�e;��M[fk���9����)eol� j ؁V��SsɕS����o����#HY���Mo�L~/!�)l�Cb�X�Q)L%�
�/S!��7Fhِ��l��6Q�x#���	M��_��_zP	�1S�O!�� ��`�'Zz�LuS,�T(*�D!�|��H܏���t|Y�N䦪Hd8���Q{���0+M�CSz
��0����F��GYn��GS�T97������%�sי��?��?�!N���ӱ���'���q����ǧ�:X�V���qLQ�z`����=�O82��NM�2�3U�qL7�/_ZY��
)4`�!�E�����ҷ(�)�,��r���ĄP��Jx�HH>�K��r�h >��&�?���{	��[ic������X.�f�� ��!>�����@dc|�LT!Y��r�1�e�|S>sj ȩm���8!���L�٨5+���R��I�D��Ί��7!FGu��Ԓ(Z=�ٖ��p����*)�'M�\���bE^MB����{����?���6>�&E���M��^\�䪈���N��'��& #H�PP�~%L�BD1�An,�Q���h�4e�F`6��lc=~�g��`����-d�f����?�Z�6 �B�|�*B@�Y,�dd�Q>ZǱ��P0�4�[��,�Q�dÍ�LL K�)�b�9�@S�k�Z��Y�OAQ"u�TQ�	,��Q�(Y�Z�rMm]�N!e���$�����(2ex!#~#<2��	ӬV�8%52��&�M�Ӵ	��"o«C�S?^5�/75䲊�[o4�*�V����^��StsbZ�i'f)��ʯ��
Eη|4|���3�8S4>����I6�bZb>&��G0�4ǖ�F���6n�u ����hۥ�>L~C�M1�!���(g_
�P~�~R��V�l)p��K���ّ-=�U'�R���.k���)��0mCкJ���z�s(��׉�C4��8����L3t���r��4��L������v
�1s�ULS��4��?B)�G�Tgh�8� }�)��� �AJ�oJk5n�E�ՆP:�cD�2���ڐ�G�B� 7r0E���b�:�	�8�Ȣ�	I����+��Y*1rH-m�������YHki��Tr�mr�r�%�VyJ�l	@���5�()�>ǔc�V9#�F�f��,����v�B�:5�VVRh�k�Xo@S|H�#©+RBD�56��G�o$9�I��_-�D����G����V>Й�� �e囶�8|:�*'e*b�4��<SH:�ԗ�1�� s�[a�s^ѭ��p�eU�2�&��1Pn�E��R��'��s��1��~/�SK�C�%>��B9��䦓������z@��Α�Ix�L9��UcR9�htꊯ(�4�h��>�n� ������%�3��X��t!�D�y��p�VtY��TT��u�����h��n],���d�ٕO���o��T�Q�)'�ĀԈc�2�.�����IB$���`��A()�|���ㄛ�`�3M|h�i�a:e��r�𙵧��hj]�F���2���9�T�SM)��K���M#�V�S0-+at�K���i�9Y)�x!)e���zh����(4x#�Pg ����I�	���a�]^���"?|��۷�._��pC_f���"{ӛ�]9>����������z!*�����q���:-�ͻ�yr�=�xxr�\o��ns$�ۂ�g>x��^�秇���^7�T�=\)�H����^]���õ����z��j����J���n�|�� �H��mr�Ch}զ�aۖ|�q"��f���ګ�8l+��s>X����@7f�/��xꦮ���>ҭ\KVg}v�E���ݰſ��n�n�k�*���ͺo�N	S��MǨC����:��ԥgڎ)�{S��B.�/_��	ڿy��s�>�����ݵ�z���/^����^�ޞ��[���Ry��ا�vO?�u�|I�Ϫ�����ۋ���.�οx�~����~���SI�~�{'�P󵪇ηV��12!�*�!�Fx�ϊ�q����9N阙�rD���k���<�G+1����@�҄�a�?c6b�'��ДN
�+�}}���ҧn��?,Z�(:Vbc/��c1C��2�M��LM��g�#�N���BF�t:4�Rp�n!�����(���-*}Q��ć3�������z�Ӷ&E�"S�*��c��J�����cYhn�1����G��>L������z�[ߒ��}=T��p�4�]�y��������Չ�(�?4y����돾�����:��3w9�^:G�7y�pu�#���8:?_�֏MS���?���^����_��'?�7O���뻛�����x������O��`�����r�;:V'
oE
YT4����":��Ee����Goi���!�@��d�������V���[�@�놑��ķ��-�N��.~K�-�d�/^=d��-�1r�1���B�8�v\T	k2Y��p�E%^��r��]?�{KGKj�JR[��rEC 
���>Fp��^۾�RCfe!�k�P�UZQ�)f�v�D:#��r��J�lԤ1�2Y��
9�3�\��Z�c�V��L�8)!�8��Y�U��+b!@YN2g�,?��6 �q�h����vF9Т���z R�*���:L�4;��pLV#�N�r��-P.�Ӏ�V:-1�w���D�E�5	ѕ,"@/"Y@H'���FMrبɲ4)��uGJik��>�IgS�7b
�1�0��ь9!F�ycQ�&�$_�\�p4F��*]
�UT"D�\�#� ���!�h� �����Pf��OE�]����{��r�e� ����r��W�!��aե��.�R��D9�$Qx!Y�֩b��P�V!��_��_���
�ìn=t���!��b��?�ʙґB�O�&[`��_"_����=�1�S��p�DL��p5�􍅪�A(]��cE��D#C$Vt��rU�XB���,cQ��i�"�Ё;�Ul�(Ŕ	I1�{��D����#��Ę�����q2Y�
��q�kպ��1r��'�� J��*���ȧ��̯s�^QR��Ї�%���t*�\35 D��eq8�K���h��1���A�k�3e鏲h���B!Ȝ|�Ʌ��yH��ա}PMc)#S�=��g���K��o��jk��UW��s�9�ҩ�)�I\�JKD`�:�L9~Y�R�J$5��4��nd��`R�����5��t�1�� �S�"�e�^�M�!��&���E�D ���D��ޢDe�!��I��*��Z�) �IJ�������d�����jq�"Y�b�J4F�lfZ��;f���7�8
1��hF���zuubj��y���Bd�&�`��ɩh��QN_V"��^JE!�㣙�ř��FH��4�Z���z�F�L��~�A?И��D"OV:�m��~p"M��l��f�'˯S=t��?��4�T��3�r��N�/����S02��bj��b$Ev�m=�m��6���R��,�>���2�d���9��00|8���rV���,Au�8�M�.��Z��r��ֆ��!�/Z'I'�3�ڠ�B(��*�Z[��B���mVaVZ�B��(�t!)��M�L�ldt�~��[E�oi�@�A��6~Rp��O_���̏���$8��h����,�_��H鲀�M;�!��������j>~�|LY95)E�HmLQ�f���1�B5P�1P�;FHg5B�:j�"������)�%"�*2�P�d|�!I���Tc��є���l�C�T��2#���|,W4�RZB�����$�aV�4<Z
F��S��q�KV���bI���FY%���`�3�7-e��|�2e�)2$>��s��!�vu>���RF�NM��νMo�J	���D��Ԅ�����|�߻�*N<�un,k
��,�b19@�6l�p~�p������4�2��
���I����W|d�\
��d%^�SN9NB�#���|�'>t���������>����x�w�;�KI���c�dw��G��wm������B������<��Se��9<>��ֽHdo���ڃ�g>0q��&_G��������_��1�g>���CE��E��x�����\_�2������_���5}������9�|7=0�Sm���o�tk����n{ �_��Ktz��t�[���~WXO���6�k��عi��z2���c�.q��> �������7�"=T���n�y�ջ�d==��>�q��|�W����t� �����;��;C�oy� ���Nj�������o�عW�^�מ�]��y�qV��g9���={~�nX�#qt�p��}��7^���z���W�>��������d�t�J�CMQ�t.q�R���@f��� ������,J�Ww�I�6Ł4-�4��3e"�B��r�L�	�oJK<'���r|�ZE���R�Ь�Z8�I�/4��+
	4J�<�� 1MYQ ��?>)r�|!&�h���HUe��Ii sc�SW��J�C��#T�τ�C��s"�ַCoZWB�j ����6�:a��&Kp [���N�R�{�M-��eͪ9!�|d�Pn�� D�_������W�7��=w�r�s�p���ź�����Ë���>^���7�߼���\��鳏�~|���?=x�٫�Q�G��,�C��G�s���G/�<����k�k�7 ����m��}wuy����~�ko8���Ӈ����9���Ԟ>�-���5�rԞ�F֢h�Z�Z�f|�lsh�ۣD�88޷�)d���dG_��N���D�t/"�Y������L[�]+���ߏiɡ�KLK�pM� p�M[*�9p#��j�>V���1��4�EK�L�;�����]��+��ԌÆF�����+�=�S������mqC�H�_�3���ԘQ:eC�O���P��.&�B~�@H�ru�9!�ϼN28ZL��2>f8) ����T��)_��EVTn
Q�G�42�i`'�Ѷ{I��ǂUHot�����mOpziy��f��kF9N?�ڨ=8�h���C�M�:�t�N{���L�U�/�����(�j	e>�_9d�ِ!��"@TtjA�r��tL�F!:d�&+?�B�p�@"�)G]�iƇ�R�8�� �0��1R��TBGu�hN� �G��U���ڊv[��Cp�ԜH�#Cp��������y�8�|̢�L'Eu=�Z��iE��\�i��    IDAT��:]�R��|d�Ff�.GH-˜rr�����%FӾ�V�N�p�׈s�������N]=T�,�[P�O��O��R@"hFS�k��*�1�|��9�Ha������"�nd�)�@pB���A�'+Q	S|N~`jô�]=�U�&�� D��6�?�Z�9
6��/%D��Nʴ�R�S��*E�9�8d�N�Aꡩ�]]Kq��5|�X	at U�)Xf�T�C�&B�8|`=;� ��K׽=�vu�{��HG��/1��l	{b< ���?�� C�m�-��&�\��=���}���R�\���/s�����v諸��Eٰu�:ɪb�uLn�[�PQ!�JO��D
��i��󥈆��E�����ۆ� ٍZ����,MK�sZ8YL>�4�6B*����� )���rL���!Rv��c��0!��d!FU&�fE럾1��Zŏ����B��:�>\�~�tXC"���&�t�JCJ�� �%%L�����*���>M'��I(K:K0�é�z�h�I1�&R�9R�b�vnpJ���%�M�hB�$��V��!,
7��R���n��
QB�S�2N8K��)�eUdjJ	�,
l�CDij��P=�@HOP�@4��j)'��p�ґbZ�tvqB� ¤$�DXYI�"�5geM�h������>;�aZ?����ǵ#�6�c���6�4&d|�ouEk��ytG��I�w�,ZK��
�Ʈ8_E�)a��&]bZ9l���5�©sR����wZ��� �t�J��!��d�Z���
��n�����S3'��� �l*����N`1ml�롊l4%�����'��~t%eV!Q!:���,9���KP��e��*Z]
���g�	)HA�B�����h��c�,�H?����1���B?ƈ��(D.�2�����E��A'N��|����8���h�sJ�^��&����eH�EH�o`���.X�;9-�|S�Z��qh$�ʅ�ӂ4;�sp�PbM&¯�:�:$NS��8�!BH��@�r+���(��&բ�l���O����鷳�\|���=����3g�@�h8�U@��B�P��h���� ��)nZ{���v(Յ�)*�} �uiO�,4�hvr7�~��Bʥc
a�������7��$'�?��? ���(�r�K�9^p��j������ą +dj�В���e��Q45~��[�4����B~��Hʘ=|D[�(�@ �K�"��L@�A���Z���{xz�������������G�G�njt���ױ�z�� �תՠ��a�'�wO��͵��|���ၯr��zK����=���ʸ����m��z�qw�����x��G������}�چ�Ϫ=<=pw�����k��kC/>��л�2���u�4����E:>�����>��3��#ԛ�L*�d�D��8=8�w����е��{���w��o�����޹�Ci]~�p��������g���ܮ�6}/(֑�>*�͙.��0�}���� \ºY��N$�{��ֽ�� }��玾���i8X�f�N9>f�7QݟC�)qx|pz�Ȕ���ίo�˲O���]�vp����o=9x��ѩ����g���׽�'�w���c��}5�'�Z��G�{���_[��WW'Z�g9��nķ�:�������PJ�I-���A��A�����3� �ʹ��SC:k���6Q%$�VWb�@#}8�h>~N�"�s��$���'�ր�Ox�����%��B
щ�Y�޶�G�`Zb�i��Bp���+G0�\)�@�Q.��s#p�0%X��ִ�Յ�B(�JM	fs�k8��K%V7A�ѹ�96A��PQ4~⢜�S�N⤃3��5�k�tȗ%�Iӟ_��)��ۄ9�ᕇ�WH�p�n�����kϽ�����/�����}���w�n]�_��_��9��������=��{sq���囋���^���ۃjQv��Fy����I���m�W����-�n�*A�n���^F{w���?�-�v
�k��-�c���#��9v>&ܻ�.�
y�S`S�!Y���]{��T����Ob?��O�X�w�%x��d9��L2D��Z�Y�!��q�IU� 7B���u�R�hB|��y�LL{)`YR���.em�A����v��J�犯�lt
R��/��PRȦF= ��%���8��=�gU�1�a��d�Bfk�5��z9�"#�+ڃ|��	q�����\����~�¤��Pv���ҟH�0�9QB.K���O�-�,�!].�w�Y�/��N���S(kJ����^�������zv�
a;�41q���p8Bq��Ʃ1>NE���hY�eՕҦ4K����hB� ���K�N��� e@( �t�,��^�B��Ej�_�NR�	��T.�N'~�8p�8���8|C�E�(�wd�E[o�LcJx���,�.q���*�9��P�6�*�CY�����s�DL1%rp�l4-�IG	>>~���w�ztxj����׫�s��x�xd���!#.�PZ��q�C��S��4��H1L����<89fQ62��lM"+���]��Qk�gt8��"�p���!BeE.�)k��!��F��`�v[G�G�cd�pD�4��B����j2B���!�s�4?+B ����oJ��5\�\Ks>����i�r9r�Q�� �p��L�)�^q�
�:[�Ro��R��i8&��B�Mnե�!��,G!|C�� ��d��9,Nn�1Y)M�%��5�S�|6GbK���-=A~8���5�= ��֞r=���Kq��M�R�=�6�B[��5F�t`�p�RL�����t,�z���(f�u���"Yz�B�20��!8���F�ͩsS�"S(ש�Uhc��W��*PE����غ��RX8�P�r��VE��a��Y&$
���N!z�L��d��޲�j��L�lY@�dq�:�ܦ�h(^[
[���*��Њr�֏i�wD�g��1���G��/י?���:�X��,�P�Xd��$��#�/Z��Pm�ASK(+%eMZ�)f ���r9� G�Uu�]YѤv�D�9%
��đ� Z3|kLKt�IM
��ƯV�hJ�FH�x��)�![���az�H��zhlJ����m	%
%5Y��r9�Ԇ�4q���*3|�H���X�����2'qHj��Av�J��wrj&}`�2B�e��N��[)�N+M6�:D+��1Ҭփⶮ��q���)1[���S-)p�t��gk�NL� ��h�xn�::q('.mv/�n�N� F@����l���2}
����`���C09��ka���g-D�dq�m�f�6�ڮ�uy��E�YS8���J�gm/��?U����Ӄ�6�U ��2���J�ZiΊZ�4��Ĳ�-QV�D�2��������)̔B��4m]R��8�5-hЯD��_�\�݈C� �`r:��&�4$&���l���(3M9Nd��NJd�\���	�Ưz%X���ag�K����*��i5��@��cp�_���/��/�����/zB��������o:���_��#U�~n�e�Un��]2����L!�1)@C9��V	GB�c*я����N:˔.�	�?R�����՝t���ե���Ջ��� Tw4nq]�s��� VƵI�}=� �q�n}z����������r��w�y:��7G{�.����u���JKa�׺[�aR��=�����������t����Y����ʃ��^�=�=���W�8�[Wݿy��P��]�O�=�AT^e</��*�?��K�j_�"O�z��{��K��:9G��F�J��N�U�{.]�[_8��98=Z��vN�����h]̾�<}|�Z��u�g������M�d�|����2H[�ou����f=e9M���M�v�T�,u�S�B�xG�{���k���6}N]���߸����L}=�U�x��������'g��=�p�y]����S'պ��u���F�����חo|;����w��=�K���˫�K۴>��7�m�zեtj���v;��Bu����>N[K)|x����!ֺ�r8���Ԁ�R�S�6"W��Z~���l-��4��"����d��0����,���^y��1��+�����>�B|ʦ�'2��m����Ɩ�Z_���2�C���~x|̐�'kj�L8)H▉�H!і��0���NX ~��8��׏i��R����6J�X���8N:� ����B���d�=^o�r��o.}!�ݕ/��o���^�kϜn�<�M��ó������Y������W�'O�^����/..N�n�;~�P�]��:z��\�	�W����s��װ�2j������\�Ԁ7=S��\�� ��Ѷ�n� ��u�{��6DVN��C�#K�:���+�x�խG2_"�r!ϓ�=<O��f�_�E�wK�m�	W���*u� �EI�p�J"������m
�`!|N���}ZN�l�I��AZ����Wq��5�5���+T�z�7��c+��&ɭO��7�=�C8�T����L݆����N�=diF 
�!��V�vO�8|���1�'��g���"����pl����������.9��'4�r�����kí�ɇ�O <�i:=�:�l)
F����NeM��u8-J3F�� ��Ү	�v�N����������'�c*�r�\"P��6d�������.6��NuYB��ԛ�u1s��
�Yfj� wL!�X�\!Ô���P'FYRZTS�����]1+Z��NHKf�`:"O
0�UJ!"�uV �51F*��'i�W԰4`G��i�V�(�h�,�6�L'��p:�����G��C�P(%�u�ue8��J����Z�lb�3N'�^?" {4}��'h�T�)��Oٵ���G;�('e+��+��<��4�uMS���C���%_9�Lǟ�,R�4Z���D��8��{�,)V.�h>kHwu.j�FN�)X���@��б8�؞���F���u�l,�t{���UW:Ǡ�bjckm=*�n�3�h �t�L��G�)��e�e�D�X�SH� Ǐ ��7�z�� �������a�6ǩ��\���i-)�hr�J���Q�~<��l�s�z��@Q�NR|"l��ʝ(�0N|��ZZoO��MLӗn�2>��&�r8�<���l��S��g)hr�R�Afu+TK�@��pcSzx!�Yu>ZN>�����#�P9�����k��1�S"%rLd�đ�!ҳ7��:x�Z� k�N��0F�)�4|�E��l�:"d�����*�����J��̪� �9|�rl�)>:R��`��r(O-`�!�&Q!c^fZAd�Z��XbEG�f�"��&�O��>˂�F�u�B��,>|��\8Gt��@DH9N-mH�B_��B!�Tk���h����'R3�����SWo�4 � /�c@���]�8SWN6U mi"���G�V�)Š`48�,\
~U��rG6�D~ônM�[Z��C8UL����!�H�gH`����]��i���g[��QK�����؍�NE+���rd��' ��D��#Lz}F(�M�a6�Sn��F{X�~�/+���"�@�A�
,e��D���
�Y!�7�Bww^���j (�E94�@��������@`��s��THT�t?��FUB��S�]_'!lgx�,���y(�L���J@��@f�F'g�:˴�B%�F�,�Cg�DC� ���R�k��1�e%2�!T^�9%L�ZQd
�h�i�h��I�W�M�Ze��p�pֶ���3���%�dic!�l���r9� |͋���,2�D�Ā �M�4�@̊��
5�!�W��E�T+�KAU�5*��c����9�9�5�*9i�
N
C����i'ZM�F ˧Ʃ�0C�X����j ����ɯ���!�ń�_d��a;��h�ϴt:U(C������ʉrj?&�\��	br��	�_�<C��ȐFR×�Tj�C�$�'�Y�*T�{��j�\�Y��ht��ɺθ}ءq.J�ޯ��e]9\���S��?Of:�ř�m*[9�+�\��a����d��������ό���Ǯ��w��i�FF͊�<�A�.=*]q;q�������9<�ݏ��o�^z+���t�v���ͩ���Sb��~{p�R���t�ha���{6�]a\G�Tc�{1������ ������2�>�&u����S7LY�����^�l	����ɓ�Ós�C]�]G�/���!i�b�蘮[@�>���u\��9���v8^ޫ�=}��jw{�v��t���-Sʌ�������އ��//^>?�;y��ᣓ���ޓ'�~��ޟ���H^/��s�������|���'p�3�W�
������l\����Z������3��V�Kl�˖�&�
I1����f��?~�i
U�4��C(
����`Qc�<�y\�bℴ�h|!⻂���T�HaS��B3�X���[Qx�FN4�wi���tL��f!4#��`!�)�||NU�#�����Q�V�)�2��B%�yB�7e:E�)�GS���&2��[q��iA��B�:�(�Ϧ&Z�Vg
_����&AC��K�ߛ�=�$}Ƶ?�x���'���{�����[OA���>���������%��g'�'����o�.���K\��7ޑ�~2��[/�����/~�z��Wmz�?������~��G�p��������z����CA�X������;F�����'���1�@��K��oL)�Z�-T��BcӱF�ňh^X��{Kӛ��9��Fy�ݮ��{gܫ��
[mZҒf뛴&<M�պ2_�!�v���Ea�:ޕK��Z�vY�*�+����1)�W�K�w�Z��U�1����aEY%�K�Ԯ�N������PYM�}*�j�وé�lRM��1�ۍh����.���88���Ӵ��D�R`:�t��_�?��>��s��?���I�w��P����.C"���l�9(nV�D�����]r���%k��,S>'�P��r9���"�H�T�m��r!�"[���̀��Q���4!Y��I�����yd!�����������DdAr�|֐e9��6Y�&��iKv�ק����y@�����8��(��/h*���i$�(Ô5UE	��,����A��)�,��+��t�(4u9�h��2��i&���5 ����k58^tE�eRv>�{�D���4�䙄U�K��^����!ȪP���G��yQ�%�U�aқuA�kZ��^~�I�BS�,>$bh�h�6e)D.��)Q.jm[.GHz)DZ���-9���SE|NG�SW��Q4q�pS�V
�+�B���¾��毓J�����kO�M�?��*�׏����s�id`]��2e��1B"�%ć���I�駟��GB��L�3Ggp���~d��*�:�$֧)_���@��rB��c�SW�����FXi4�%sf�Vw�a��Z�	�<e�6�CsȜJ��O�i�Z>�l�DD#�����Bck[Ȏ�H�O���k��'1$q�A��/�,��sChZ�DKVS
��P9V�8���<��gZ:B�C�����h�=�E+�?�7$�t8�1�9�n4����%K7�l��-��6ʝ~����i��Q��e J�ŎZN�~��"�60#�����D�(Ԟ�8[�im�6d�s��S%MN"��R����ɣCT�U�2q�h\��8
l�IL��Nvs�YLx��؉��"�[]~�|"́��e�U�|�GJ��'�~����PM�Qi���J�F4�DU:"��鍂�GJU�pR�3S�AJk�ä��2q��4����=a;�B�l�Uæ5P-!H#BQ�jk[����稢,A
k����юM]&B���|ӆ5�¶?鈖h*d��1'dj �����)>�(p�ч`4#JM��D[æ3FB$�C_Eþ5%ȩm������,.�����)�`�qF�?�y��	yj���Z��;�c�����UNu����U|�� �@�    IDATdՒȊJ|E������"bZ��TK4�u�v��BX�SV�9<!�,N�	j�S���'^�(������m8����b��Y�)�rF�&�J��b��7>�@Y�@ʚ���FC�7M��05D���15�Xd4�(=�dRc�(2�#�&��Z�P'�r�DE��Nzu��*N�@YU!���rB=d��~rJ"RV�B8Fx��@Y,�hb�䖓?�Q˙�C�Χ�!%XR��$�"5�D��%��n�?��?�E�oyެ�{��)�ƈ���tS�l��@�>��
�
�yAE)C�$ہ�I'�8��������"xJjg8�H����OM=�����s��L�Z*z<��w�ܿwx|t��l��i�����}�z�R��߲i�|�wv���g�Z�>���č��__�]�sX���ٽ��t�Es��k�|�酫g�n}��#�Q��K:�z�����cW�OϞ��ؕ�Wބ��}��/�t���KW3���͸S��N�b|/���㨭�aZw�.��~�8�,�)���η�9��}��Z�R�eWV������v����]�i�����K]�<�F��A-z��?�[�X]tYs�1�=Q�]+��v=��5�oo���}�q�u[�Y�v��LqL����3I~�w�C֙Cᗿ����ջ��/���Ã�7�_~��}:x��C-��|�n��i��m�[v=\|j՝o�?p-��W/�y|jS�]�W�K݊N{�R'!<�SkA��:��y��D�Sg�c!�i+XӘ�KX
����p�ү`�F�]��Yʆ��\5�(��pv	�Kɖ�(q�P�*Zr�8�Ȋ
�D�k�P�`V�tħU"Ȧ��h��$Ve�2�(������q�B0�M�$Ҭt���7���p���)�_���;4�$��,��EZQ^�h�,_��Dc��2kC���4��l�f�����_^�<=�z��N}s���l�}�	�Ż�����=�꿾��꿞x�=9]7�ߺ��Υ8:��?x����7�^{^�;�v{��"���һ��W������e�f{ٔo]��a���3������� `BT�ޖ�R
7��)��Z��'�-�QTHV�'Ջ;G�	�Ӭ7�5���J����M>ꃼA�"�f�+
�ξ���o�Nϰ2IjׁzF��X�ۃ�U��#�19��.���wۇ���J\�޾M���E�D#���GV.����B��u{$n7�w65�*5�8��QH�v`��I��Rʹ�Y��ek����0ei��*JIS�}�����B�D�R	!
	rhj��qJ��:�O�p�>��s��s�cƩº��(ؽN!强{<�����S�#G]G��D��HӞ�m�\���iǨ�k����U�#�s ?��W��C	ġ�������FNL����!��R�(�ͧ�O|�tRJ�q�Oh �19�7�瘪�&�5E#Ȋ�[xU8�8F�l��9��@�4�zÑ����k;��|�?�t�(� e�#Bְ�*:�L*��G�z��:���~mp
��t�#(]z��b��*����1��P(+�g{K���ex�34�m�4P��9���a]i���>��?�3�6�A 2N>�f��_����1�"k�R<!���w��K:!hR���A�%�`9:�s
�p|Ȍ��q�b©bY�RE]���U��(Li��R�`��M��)Wb��`��(�?�Г�_,��hl�y�**���" [ZE��V=)��|��	��@H�BY	n�+�)2K�kh]�4���VR-
R&�C��Ƨcu^����P�� ��xL5�Ρ)Q����(JS�dU�"�&�);N��B�0m��d@�Ϗ��)�`�|!j|��o�*�Z��TH����r��P�R�hl��s�L�5�
��)�G��A��b���Q��5�R���)ȗE'BE!v�~^�~�!eS�&�E�i8�R�����i��׌(A~)��&:����U~;p�u[Q�����MY�~(�c[�5�,�>��\:�*�S"��D�u~R@���NS!��qxcw*��
9���||�4Y8��dO��{D��B�XL1�K�4'ML4��Z�(�_���Ƭ�j��ɡ�H�E��e!��c)�e�+A���H!�'���	��p�B�8�q��\3p`���H��'hi阦���M���9Y����Y)���,SNU*�"�i��8�@�D�"Kj�!�OL~�t�~\O-�օY��gBɚ&X"���䛖kʡ6�����@�L�#Q�R�PH��0��|��)$�2-���
m��<l*��|�I����Ȧ���)c6vu
I�اI��)�ǩ"P��8��O�$|�9 K
�@k��#�V�2�(�#���+]�\�:��^J= GHM�����(P�P����S��rk�H��<>��$��1�$�7�D0����Z�5�D0!lǴ�B�&E�Uә�N�K4�hX>�D�b9,Y����t�ʕ(ZhJ#�25�
�ɑ�IbP6���X�4G����H8��#��9ja�\cd�8�*�=�!�
�"��>�P���.��l; ԕD�B��ܴ���JE!`�'��5�?�%Rn]	���C\4��;)qXm�e9�NL�0���3Q���I��L���B�b���贍��|��I�E��9��tҶ�41!)��׼Ƣ�Jx7�/���k�_B�Y?���M���4U���,BH>��Y�9$X?�hX�[�N��|9�[�p=z��� ��ɮd�c:����}�����=}��azs�7D����;*]�t2:P>v}*�:1�y�B ���'����n���l�g�7W޷�������{���7��}���=t7�.���?%����ώ������ѱ����r��z~Q�y���uʭ�o��A�`���BJ����Q=��ݜ���r�'kt�wm���r�^�{��(u<9���y�w��x��=}tryu�ww�
�[�Q��:�ΰ��C�(;ܡ	tP\��r�'%Μ9�k�ޞ��o��o_�|��SYO��C+�.�������w��nN�޹~�ʗ�^\�=����b��9}ts���}9����n�W_��푯/}���:��큩�Q���~Q��s�9B�:��($B!��i�Ҍ�ڮ9�Qh�f�� ��]�v2�2;���\����G�DL֐kpr"T��#�VLh��KTˈPbVH.�NH!�S����pH�JT:>MrY�e�+���05HC���n�a|�]��(+<��I��F�7���D�h%�r" �l�s*�j�%�!����&w+�I����E0�N�Ʌ$�H�P�C�/c~��q�N%�p}�������{�[��C���O�>�����������z�}��37����M�u:�<�m�����;O�<�xԥ���#�����~k�M5.az��!����4�a/R��z Z�g���<'�0i_�*��! � kQl��9�a�dS�qYV��>���ƙ�|L"ޠ�-k�����XE���he�ײ%�uB�Y�j��#>-Q��h�"M��F��H	�	q�2(K	4E�á`p�X��Dɮ�o���p��)�+QxH餄 Q��Zp]�2�)����Ъ��g)�z�F$���7�-���5��6-_�Q�����*�:osD#H�V�Q�75b����� <}6�3����Ij�k!|;&�#
�_�r4Q碨3ʱKa,PKQ:����C��N���!�s�A�!"
$ժ��ڀ�zbE+��"��EJK��wd�F�lS���P�O��#1��&W�5� �7"G+�Y >�Dd�K�(�D"�,����nhB�g�{�
�g�`���:4J���ZZP3nj��@�Z:��\r�p��RH�ΚEC�N]�mW�.�Z������<�:�5)�>��˃�10��A-ێ�����ǂ[-%��� ����qJ{4Y�?G���7�@���:T���c��Du�jo��!,_�G���l��9��q�6��g�Ї��@��%�m�ÿq�[���s��ӊ��&��������_QL�:��q�A�gɒbUd��SȚ�(��8��nK��V�VV�i�T��Q"�a:!S���0�S"�/:颁�k ;�:�_Q���t�,���P�6�G�Bt���
���5U�¬�>g*H-ߔ!��7��1ѐ�˪[��ө�I�l:��V�V+-�#1��Vm*��RH�6ƙN8BF�,���tB4���ag�$ގ!wZRn���V����
�Ⱕ�ߢ��ր���?�)'�zi
�e�� ����4���LG�8��2?d
4�f4���Ԥ�ц�Z�[�Z�6a�JLpVA*N��������@�� )7_�&��1r���KB����G&Ĩs�)2��֌�:�WQ40�DSѦu�i�r#d�~��Y�\���2�G�b������kfӬ+!���p�9�M���,A]�iCj����(&��juҍS�b�;���7-w�7�Gh|�B�lQ�Dx�8Дm	]�.:d~��K�D�m��m�)�4K�b�"���N�C�P��l1�g�I�)d�"�N�Q9�V�����零�r���#��CmwE6�D��)M��B�N	��5�F�Vx��v�TQ4
!��ي��[�l�|C,�~hV�&�i�!�q
-�M�6j�v�����vj��qA�6�#"_J����PQ>��=?o�@6�X�V@H:��-�7��r+Ě�3!u^!�������R�3��'d9NK b�76�%�.��VSgd�\��SN�#§Ca�XRVt�$+�f�&>pΖZeS��di�	�~�IqjX�����B�@H�>��}�*Ǉ�q ��hJS�Mp~8����1#����k5)[ѩ%��ϩ�h� J��7�X �2�rMEC�J����Pcd� �S#�2��M�/46A�^"f�|�f�ٴ�	�)Ĕ��:��Bp��BL�A!�엠R�B��_���� ���~����BpNuQ:��D�'�)E��=����'54~����*�_9���o]8��rX8��i�������|8�߹�u�]�[>��<}���^lKл{�H����iprz��Z��@R�85���_�y{�c}����?r�e����]��~b�1���n]1=��v�ׇ�Z��{7�����Z=�:��g��ެ����G��n�ۻ>>tYէ���Ϸ�={콚��W���r�;*����8���/�<��.Oz.�pir�J��M�ƿ��\͸���v�u���޾��.�o��t�򍋔{vTY��f������w�3���o��v^���6v��Z�[�NONo�o/֎=d��өy��&��v(Iu;X���zt`�J��_��	����[�;�����ơ=�r4���ï/�<~�������Z�}��~�����ٓ���˛Wo��W�ݬ���N���ߜ��?|��ü>�w{NPwM���~ؙng��c3\��uFmd�ej����S�� Y��$�t�6?�)'q6��%�_{�ɚN2`6"X�$)ΔK�N
��ZYI���R�9l�r"�XE`������r�g�5o�)�o��$e:�_hjpR�u�����L��U���̧���kOЌDT�-
gkF.'t�eG!~��*�u7�o�~Y1�`�ILd�\-�h�	I�.�=�{��O޿8�/��no|
��_�x��^L{{|�ս��lzB�/�=vO����מ��vu��K�/޼�\�wt��}�v���,^��U�WIo��LV85�%��?�z�R��yKP{ނ�sb�[���j�e�[<�C�WO��V�
'��'%Ԁ!� q��S%����>�KN���!P������3��_��_�e/�Ps��x��95�[�7����� �V�^�]ݔ�[��5��k�-�)�o �Z�ܖ�
Ek� p�OʒY6W�_T'Fǆ��:�"=�U�Ǉ��^��6T9dg��Cb�h@�8ӧ~�L�ZB�(!Sc8IApX�6��1�_ӔOa�iY�GӒ6�e���7ռ�M��9�+���aOl���䡦1'�S�����G߾9��`:/9�% >��`��fjQ8M5��)�� *�m�v��sIo��R�������R��M�@�$�����B���e	՘���K�I!j�7�ҁ��פ��e	I��c��@����*�Aol`� ��<�v&�B,P���84E�8YV�+�P�r�ҝ�|��c���^����S��Ε?g �@�L)�A�(�E ku8E�@ݲ�iG�c�ր�C3��ֳ��+�ps�����F/����R��,��.g��������l�?��ϼ���!`]�̹z��������Q����B�j�@�G��_Ơ��S�S�L��-��M��DvR"���"dW9)x���W������" s�j�Vi�m��ju[�
K�nx	75l �(�N���|s�XY���4L�ʹ�� ���^��퀥���s�����#�Rϣ�1���v�9��h"di�.��,��d"�E�u�X?�T��T���ӵ�x�����*R �!��#Ԩ���L	~4��������r�tj�PY�4~
9Y��N� ���\ C�:�V� aE!FY�!�7eM��|9��1�@j�aGdp��U��t)��)'%Dt�;��!F
������3��7&2)�E��*,���*�����_Vk���+w�o��Ւ2NdS���·W����89шS��Șr;O&��X2�L����� d9���T4Rm��oׅI���|���-J'p|?�[B6M���t"5e	"��u[���8Z̔Օn �3� |��FG'���#��K��v�)�R��im����<��XW�pSNU8ɦ�VSQC�,Dh��@ȚV���O�3�|#B6eLbppjIbx
�p��)-ec%o��dU�M-����rB�" ��b
�J�SԔ�Rt�=�Q�zm��Xc�AJ9j��,�LDM?q�4�C��AF��N �.n��T�	l�5�-g�Ka��\�*N��e�5�Ϗ�8|�? �c�V��
�v(eu�RS�DS���r��������׹i=�?B8�N09B�@Ѧ)��T7m���A 'Ά�Ω�)CF��VQ�|
F��*�.��
e�m*��C��ٯ�X?����|��WwW-� �C��*�9dk3ex�cQ�\d����3��Z�nL>�8E�@��V��w��Y;���lE��8���s8�W1f]!L{9�5Y�g�G0 �i!��DW�@ˉY.�t�Q���q�/�@��������8I�_����E��PG�ߎEZo&�[��/��.�sD"~����E~L�����n�8�:`�t���1���$�u�Wu��ӛߞ��FY��-���5���(f�8�KY�x�c@p��jL���-��o����NwT:o���t���p&�t5[%��k݋�����|��~u�ڝ[%ݑ)�s�ˣބ޶�+ʍt�,�������z_���]Z\�ӓ�o��l�z���������S��=8R�វ������c����a��5�݂��m��_���s��Zu���O�:w�s}�������O��k�mtK�O�����������7�{�O�&y��[C��E�;6��v��l���W�ޭ��\��u��ܛ�^���e�_\^�ZIn_���x�����n��N���Q�p�L��lR)���;���8[֯�.&�����vr|�ĵ$�}r�����co�r��`\�u������ŋ�_]}����쳟������������>����Y�G��ꬖ�)k�y��[��!��(��(���%��ҳ�@�1�j�����*v{Ck W�(p��ko���ݬ�!IEf�2A�hjS:��#́���G�L9f:S7��8��)}tJ�Ihc��n����00Kd����PCi�)T(5��s�X�c<�=� 	�H)W�9'ڒc��h�*J�=u+�Z�\~�r�B!�i>�m��7"�uY��	�2���m��    IDAT����~��_���or|���ɻ����'����<������#�=���|����kM�����x�&5~r����g�'W�@w��-gϿ�	��T������'�|�zj/(���g�}������Z���]b���Ak�c��l��m+�h�ҥؐ�g�8��I�*�~��6��gazSQ�p��%U|7��[�w��Nbӣ�>�HZ��[����I]��>Z@��W}}{��೎�WYOĖ!��ѭ])9�l�%IA���h�*���l�M�O�_o8Rz9��0ю�BJAz[&j�S����.�ӑ۶v�q��K��8�!�u��0Z�eEq�MJ�t~SU8����W����J���Z&��B�Hs�[����ސÁB���	}���M?��֙���4�����R���uQ�ODudYh.��Z5!�ݐ��i�9!��<����P�=�Yj�y�×�F��*s8z�A��������#p��2g[�d�iY�,2��6��@k�_.���G+��҄����x�
A�C�t�Bh�.�MS��F�V-�cB�:d-'8}��FkoSN��S:��\|����?:���@�X�G�Ҟ� �v�����K�	�\{"��(�PVbk7Օ)�!p���Ih �3�B��B��Vd
TΊ�����&��_yD��9���1�a�� pR(jړ�VX�G�]�p�h�fjOJ��0�FK��A��9YK�	䬄��Ԡ䰍��J)
���sF�� bZ�����N�5jg!�$�/�K�2���駟�=հt��cǨ�r��j5�陬\"8�8�XQV4Ĵ�U �,NL�d��D�D
��Z�>!�AhH��5*�)Ǐ���n�}����4髉�/t�IQ�#=�l;��E9��=�;'S�,�N�pR6+�h��J�fQ�Q��T��8�tL1��D����EMe��,�V�m@�Zr���0��\�m9����1#��Pֈh��V�ݖQH�ȤCf����
i�58�� L�,�����	�A:�S�#�N���/���g��j�@>G.�5ݭ�U�|Ö�C�Ȝt��e���l��Y�4�%+�l� 4(�EM9�p�i iA��.�B�zH�?���0k@t��_
~�if���:�A0�%>�¡`p"���[d�B�m������(@���'��g,�PN����rY�)���RV�V{V�4��lUZ�(��X#�A2�Ӟ���,��G3)[�ߴ�8ēO
+�̏)�MT�Y��,���	o*�Br�!r��с��iEh��O�Q�Z
�p�Q��
Ab�P
�~Ѷ��)�#��,�3�u���t$*��'+MS�n�����uX��i�A�zH���-+�%�Ζ��t��M�@K��!�|ddgP�;��u�V�N�5���h�$$6��s�%djFY��&���y:��D �Y����+�&K�� MGs��v@ℬ��UhE�����%�s�B05J��.!C�ŤSە�t�mT�DL�:a����k�|��)�����72Z�c�h�j��h��Y $0!"*�r���i��G���>|�Ҭ=
R(H	����h�(;+���"��6���ǟ2�&Q�ߢ��Ĳ��o*�=���a�k`�Y�9ÄPc!�fvAd����-5V
��!h�O��S.pw������,�~4"V[�&��@�A#����6P��Y)ȬtC��#�M��d�E�$ɲ��e5m[�re��fe�w6D�!�4�O�M�c��L��'^05̞��Z�/�tu��ۇ����R��ֹ��w<��~x���)�-��6-�{@W
}�����w��i��*��X����+����xwp{�^��眮3�݌�����������w/ߜ���Ή��Q���ҦO���p{u}{ys�%Ý�ޤw���Ǔ�u?.�㺷]ա��Upt�g㺭���>��P} ���'���ƇI��S�A�?{�����[�7���g-�H]^�����X�X{��Ow@�߆�t��`��v�rMֹd�m|��u& 6BLG�?cm��w�������t�ݧɪqs{u~��*m��ׯo��{�wur���u�ҍ"W��gϾ>�r�ԥ�K��޼���|�"��S��?����������7�]�#��a��.k�Gu���ęS�hY��������Mo)�1YS�T�(��'�7J�i��波,����A����o��
lm��	�~ͰF�8)����'�Ԍ*��&����'��~�C�����mxU��R�}�[_kӄƗ����� �,��mO?�_h�1ӪL� N�%R]`���89��Z�Kو�Tt,5��l��|�
Ɋ�N��0�&+����N���'�Ml�q�w����l�㐫�햛���[��o�$�������y=���?�'{�����w����)�G��}v�����ӫ��/֕;���W�#ʽ?�ڜ���OvĽ�O���X��q�I�]S��m�V�g��^nX�6��J�N��'ֵ�_��؇��g
�l�v�Bi��k��p��t*M_碮ӹ�ŕZ���}�w�m�L��Qr��μ� �@���?���)@�B�Q�Rr�G.�6Zsk�L��OД�Ε��	B>���f������?�������󯿼�'D^ �N�M�@=;����bיww��clS�t u��!���5S
;x����?���r'�zu[E r�0%��>GJY,Z�8��4�E��7րǑ�`� A�G��~�7�{4ُ?��k�KR���o:�ѥt>�L9ۮ�3�q�/�4�Y^o��p �՞�[����`�-�u��g���כ�Օ%�B����=�}а�@6��[WB�:@Y@4�	V��i����r��5-��҉� d+ �p�=颲�c8�*&A[$d�HA �e�V(dh�V�o�K���iH����h({F2:�d9C�P�ȭ�!]
�܎f�,N��4�)���:���6��#�U��8�8������t��������������Go�[|R�#X�f<��,g]�� �C�}��r�?���(JM��r�i{ȷ'L�(�_���D��Hi]1���� ����#�1ʅ��uUX3�� $|T	��Ϣ����\�~:7<�{!��7-q�m4[���T�JS�aj�a�9�%Q
��1�q�Lz|�hB�"@s�
!�)G����T)1>�O�z�S�(�=���I��:�́�vߡ�L�u�M�bBj��:)�FGiN"��r���F$)dHk�IM4�)�&�@0*'��,�*���zN�ϑ�Du�w�ћ堵�R�h1� 8@ǿ��i�JHpz�,�֒2��t�Wh��b۩�o�R('1�gq���NӪ���$�Ӵ3�r�)�jU:��Q]k�7�mc
�p�@֙�4$B��8H��<��X��,�i���p��~�pN31!�p�('�t��Y����S��LY!�A-�T�&
�T���
�J�٘U��uC���#�*�B�p���z۵��X�_�|�O�ٴej`@!�u�"4�P{eA��4�:,E4�v � Z�Z��NT?|�3�4&0I���44 ��PR����]N�t���U|�A�M�3u!:�k�H3�tV��,1��q�4PźŔk �*rJI�J�IP"���"Oz�!�M4�NQ#��N���fp���R���(�!jP��fT����p0� ��A�ߒ~���9M�Q��r��ILvt��ζV��W��h��̗n��Z�dE��٘쮎�&�5���'��@}�1>��G��Ʃs�|�pV��к8�,�S��B�Ix"�,��iS��5�S�/�΁qM����Rb�U1DV"L���B��϶솦z����yH��-f���f"�C��(�J�ϧ68��C�ff	�!rSf;�!u��QV9�
IA����W����%�E�SRB#(ʷcB��[��9բ��Jv7�Q�&�N�|8ﱀ_�o����4>p[|ӱh��p�8�����6Y�QW@N�%��Iv�[Eӑ��1�����5 +��{~VB�)��FY�e�#S� pZB���h�:��KgM�UG��@�X:XSR~_f�#�J��5U���!b��)�o���d
�l:l�]��RS�@����q4)�^od�J ��I��z� ��7�BpQ���\�KWzy}quy�4�#ŷ����;$��e],�^��f0'{~ X�$X�냾�m}����$o����ͧ{���d]#�Ֆ���n}��7ڝ7��pS��._����[3��m��������r�=:����ىSu]������q��ޯ�0��>ztHٕ ��n�f�X^6|䭇����Ua]z]]��Z��=ٓu]t������g�|Ǘ}~��w�/���+�{"X���p9�|�oҼ�{u�����}	�nU���v�Tс[@����xu :L��#���,�f������1��wҹJ����������ٓ�G�Sŋ�u�������_��}��ɳ��{�Ǿ�Բ�/��_\]_x(��}�gwW����?:v�[Q]͉�s�f4 �Yg��@�Ѱ�M�L9!��lp"��A��T+�҇i����hlګ[�82U�)���Q}�q��';:hB�A��C�V
�eC�Gnǈ �F���g���x��_+M����ɦ�z(s�JO8��t����� �w��i�pVnY��C�-P"}���b���-��h�Ԫ� �P�R��z���f:BʉbVq�{�$�[���1-���q8N0��/Z��#̺���~uw�}�˽�˻k�}�����/��<���ƺ�}��{�����_\�y^����N��_�_�ｺ8�8������o_�߽y���|�"v_��3��l�Y�e�U�����EDFf���dw�h
�P�P� $>߫n� qA����+����@�26d�ۙ�������3�JjȞ9�3��1�Z{�s֊��vnx����L����՟�ٟ�ǿ��8ƛKO{��]ƶ{.��О�aK�\�)����6�k������ȡ)�m[�3�0w/�M�X�7��'Ϸ�*���[n�JG^nyX���.�GKX>S[g���9e�)�����=�DY
�|��B�ز��l� �t3Z�Q��:ZRBʕ�I��N�p����������|x�����8�z�k
*����4Y
q�m�}�h��um7��S�rZj�^ix�
�"�+�G���V�_�4"�F�!��G��e�����l��E�m�R��Dkt2x0@_�*�W�nL��F�,��]l95�Zl��AJ��4��|#e;��h�PSE�K�q�yS>���cM�D��r�R4_]!��RSΒ����(�,>�Zh�i�*��T�#����|M=�]S��I�[����Q-fj���:�h�|!���p`�wPz�X3��RDs�K'N����B@)�.�,�td�*|4����f�����X�8|�QV���Cɩ=���
I�T��(K$U�� �C�1>���Į$i�Z��:OYH��3�3��"�s.n����4�הqz"�:ǨG��L���{D�E�>�di A4���M#�C0å�28q���GC��Ë�Y���:������EI�.;�~=3|�jTa4[BR��+�}sI1z<����gS��4��"o�޼�e�5�i-���Im8Y����=䎗ޘ(�8kE!�FR�D��-�&��Ä�1g��L
^���ȬW��ŷ'd����ns����IX	Hk,9�󼔲��O3f�у�!p�M�9�fl�����rN�]�϶����nI�k8��g� 9U�o�	�g�9h)OW��q�J�Z��R�C��Μ@��u�r&��fm�:�CC����L�x�8��8!��Y�B�,�F4�+$�K"ԀLE�2N����>�n��8|�F|κ�� ٔ�p���><�,#�,�@��fxx!jh��7-�̼p(p:94	�F
�t��H�.��7��$2)8�F�0�)����k���DZ�*pVr�1Y�Jȍρ4�ĺE��ES�j-Zk�.D�۷ҍL����W%�(\�@>����ֳe�p�;Iդ,�h�u�O�@MW����c�G�ίCd��i�m���ZQ���lSv�¯#�>G\]8��Hm���D!,>&�Q4��"�iQ����3�M�h�v�Xo ?G	�^&�j��u�g�h�BE�Rzq,�*�h�8e͔�r8�P?�;�8BJ71��8��&4uC��T�͔ N���[�D���(=K�AD�pfԏ�ܶ(��7V�#J0�BF�!W��XB���%�a�@�	��s ��Bb��jۘ���L7u Bcʐ�n���� Guc�C)Y�	�����P�)P4�Nj	��jiMq��@��})�T-:V��������AD�RB����Fx�ʙ���~rR@���F|~���^e���B~�&K��!��~jY�(�2�c���&��ҵ�?�*���Ɯ�ƥ����q8��^MZ�����GK���P�(D�w=8�mjT��p���
�� �n�1ۢa��
�vYhBʲZ�)N�rL�ଔ�t�b�����h���� �p8��
��r��1�|��)ӊ ,�8u(����_��_����=%Y�V��VB���L������K�LgW�J7�a��`2>�D���J��<������"�� �7��-�a���띹�}�C=W˧-�O���v⭶�|A�������&<�\>It�o��+�vs�+��.��/�>�y�onZ�>-y����IJ������w,��e�<�OE}M��r�jY��\r|���׸:L{���{�Э���7���sL�zZ���r�x���� �חn��6�(�G�No�
8L�'�����2RZ6vk��z�k�^|��<���'��%N���}���"|�-���w���ɱ���WmG��م����į_�L�ф;jFG_��8
�	����.�c�2:�	��.�W�>��Y=zu��}X6�£����ONnN�O?�ݔ��q��u�}���ݯ~�����K�~}��ޛo�����j�g�:i���pNK?�%(��|��@L;]��z�����у�!�s2�S�o'�K��0�W��π�����gV��~x��h�b݊J��h1�����*�(G��F�BV��C ��ƒ��yp��~=Ӂ��Ϯ������"e�Rn��Y��Q�dC	�a�ɺڳ����U�e�Cu1�� w�!�8�8嚶���T��Qb�hȶ��hk�J!�ɪ.��a�!1[`�L���'�]sn�.��e}�������O>{�#��-�/�^��3����GO��>yt�t���������w_}���??��[���#��"v���������W��ʫ���.�V���ә?��?�����
���ԽAk��@_��U�6z>D��z����gB;���p_�-b!m5>f:SY)���C���$w�Կw:�v\�Y�UA�>)A^=�-�b��H�z?@Խ��.�D��t���V"��F*�_���2���!��+u��"��lLr�y�_.���ܫ������G��NN��zo����Ǒ8��sՙ,}z�Ѥ����c=�V�И�| _�L���� ���edh����R�-Y�� �M�����	7�^��J�g
��೦8��l9R�-����~����B�����M�l�G8^v�����°�v>�^"�)�\
p�D�J)$�`�4�=�,�պ�N8�k�-�\�~�:!��M0�2=�BЀ��S����1�@�@RF�P"zHDH��J7�kZ��|�בD)�>D�,�kDJ%"D�I>e~��"d��z�Bt�p��C��J,�����`Z��N��q�(G-��J�ꄘP�����1��*6V�Ȭ���0q��BBL�l$�P���$��\��Z�q�9�t.�����Vk�����>��R���ט�e��M	��o�J�
�{�xA��ҧR�(G�Z�z�������g�*Q>2MƱpN`�P4<_�T�#i�&G:P�v���d�V4r�R&Ԏ�FQ�/
�����L�    IDATW�%�T�@0g��6Ӂ����"�F�F��_Q�(Wtih�"�GS�&��0!|G���;�mi&
LAb ͤ����r��.L�Z}���D��4�6e�(5XN/��͸���/�~�'��.k��	G�S0�D��W��V��C6]�y������6AS:mT���"�2��9BE���b���&���Q��V���B�dK�(��%��t��%�Y⢙hx��ȐpS8_�D�3~��i�Ќq�M?e�id�f��,S�Q	�G>5�ï�DJ�/�X�8��L[�Ǩ�PݖR) �"��7S �����4�@c4�*q*!kr�U�SuQ�q��W��0�,�@�6��WEQ�H�Rr���VZ��͢u��1f����( �[��=��JLj��S4��gi��#�+�t�&e^kBu"��8�����]̍�.�t�9ĥ��g���6�s�#]b fj�cL���^�S���������*jD�����?��E7ۀ�5Y���4Gp���,D���S�_n��!M'�_'���Ǻ��'���NV34��HG�8�޼悟x���3��	�Т�V���e1gKR�j��i�b���F#B`c�*:#'�tS��꧟Zim3 ���
��Z>��%B-��H���h��i���U,��@d�jmF�L�� 45*gm#�8�-Mt]gQ.=�b[�Dk۴m���usDj�h��1��Fx��@D)՝('�Po��M�82_Q�!N&���I.��98�K�@R�sl>��t��D:����� &�J%"d�N
�P"R����Cä8�;�@�z��b�Om}��|����ZK���c�7�3~U ����uDhs��a
-�r8�lJđ�`,�!0�1qY�$�'BQ#�NH�N�6Ӵ���t(� GT8��1���%|[�TbUL�ڈ���8Sh�<B1�^�F������xUň_h����
Y��O�i)�,&<e�sɩ�	4��T�_���\W����)��H���Ο���U���"<+����D7	��$�f�ȩ��緢pd7���w��{Yh�&+��G�;V>�x����I���g˭�K����?[)����ɭ�Վ�*�]�:��,���W�y�_���C>��=�Z�ϯv}����ot]m��؝���_����U�7����/�����������|<=�8?�����3_S{syg��:}��/_��W�-���׎�����z/�.�ֻ�t�`�π.k��r���h���=]�no����x��w�ON���W�>)e����;�lj��'6�V�?�Чu*lc�������D}�ԇJ�o=�%��tŜ<��lN��c�����D'	G
)�H����՘˳���Oo�?x�����2�NvV�۞ڞ��ɫ���=_��s�����ǧ�[���������j_��W�}�}d��ҟQ�R��;��!�&*����d��L�����P��S�7�I�&2���YNR�T:Ac|��9�h�)�˨��8h|V�)gD��iV1���L0�[�Ԃ`�S35#�QCF����&�~� h�o�+�('T�fJ��#���>�cd�7��!
��C����^cx]I�4
�9�%��ܐB�hZQ�j3M���Ō�I�B#���1++�e������ܜty��;����::�;<<��ڻ�8=~���w���/�~}�h�<�%"��=�������b{��|��=y�g?���?����;�x�w�<�:?=�w������7=�tW����wa����-�ּ;��������曾APo�B��j�޹�v�y�a��V�dY�i{e:;t>>
[�D?9�y;K�TFG�Pe���Z��yDs����^S�2Wn��r�$�^y��[�|�U@�_��Bj��9��jA.?��e>CF�.ѭX_�r��	��cUF�����)�����ǿ�����yz��W�~�9����/<��瞟�0!�i�~���6N�3�%:!� 1F��	��D덓�3�Q���m�i�9p���-q#h��x�*�k�a�9�4����(�5��0������+�����@�C�d!��/��g�XB�ќ3�r��&ʀ*�
uI!#Լ�@~#��,|g<Z����4%�u�e�����E�p L�t)��a�R��*JD�;"S%���P����N����h�W�,��2:JW�C��)D�E���@S�/�2� ���(?��-S�6���%�VΡ�~��,��er(���ey�?�h"�D4W-�+�5�e]���c��![{NT�����$'����!=Գ���P`��q��o.�@S�}�҇/��_��$��U�w +�e�.������TH{-35�i�O���Y��̔���!��D��ʭ��:A��c�nZʄ6k�+!*��i�R0�)�N��~%Є�Dli4�N�t;�@L[��pSu�q4�����׉Q
�d����P��#d��&�r����Z��^I
��hE�����H׳���VA���C�6�[�s�Yg�x|�\����%��4E)��J�㬻^�H��ON�u"$%�u	�>G���X�&(j*��B!�p+�CJ�:��i��Q�o7���Zo9-�n]| $� ��)�N'a�R8,r�U��j��[�R`}:�sp&1����1G��Z�_�Vw�Ǉ �f:8�J��%��M�9�)4R���r�9��Ջ����8)�F 2ߨ4�08�!�4�/1N��h|)�L��ə�4q� j�Kכ)��D$r���<��#��8�^���F�����r�E2�(�z0M����BEK,+^�&T�4+
L��b��8Ԅ�GJ=$k4-7B� �щ)4�1��)$�� �B�m)ЖPTb��z�/�Ƈ�[{ƪ�����^�h��+H��r8�P��,)���4�B�Ԇ�iL#�7��L�`
A�Y����0r#M
8�F��fVj��b�JL�r�[�NL��i�����^�Y� �1�*�1�@�t~���J��/7�Sb��9i�����7-3�ҥؓ� m~ʐ�&�����<�&��߯����$$(T�8����L�����&��P|�=0�7�Eʒk[�����a�KR!�p8i��R��i�o2�1���beMԴ��s_(�8@�����N]�VM�2���EII�D�V��4EC0�N��8C⧃�"Љ&JY�|���)u�?���h�'�c��B@�ҦZz]_.rF�Ҙ%$��2���ol����J42S_$n_�핱��Č�0E%�e�rT7�Jm�e�O����T]�5�~���#7���&9�|c �iF��BjrJ�V]���
M����Z���a���k��bB���;IME�l/B��TV+�P⢘p��h4E�4:�~2m�`m~�&�Z�	1%�o�����+��n�X��k,Mj�L4!|#�)��B�%Ɂ�P�Z*���I'�#�99:� �d՞�.>�a��W,}Vq��+M�r��C��j���˹q���#I���N=v�����/g���#F=���z��j#������/:]n���؋_�z����˝���}��sԭ�F}�쾿z�g^�.O@�}�n�\�o��8([������{��������5�W[r�ɧ;}���/��_{�p��ᔱ w�q�u�,'��Z�����M+�w4�����c�;�����/=z|��R��x���e��A���Vz}�����9<ؿ<[��ig�wsᾖ�=�C哦�RѨ�����AwǍS�%���A쀚�R]
[�T���B"}6����g'�/]~��A�'H�KӶ��ǝ�_y����-�={���Ϟ<<}�u N�g�6�:�����m�K��m�z�hc����%��{�,�6�g��(�	Sk*q9����J�K#�V8��H$e��mN���B9����ި� �">�\܀��[��'�Y�&�`!h2d-�l@�%�@M9�"Ӈ��ljd�d�|N�Ek���5	�'&�I�+#P(�"�t�|!E�ϙ6(�'���D�F`UBꁬ�͖D2<�tS� ΀�	���(W�U4#[*����>��i~����KWl|N�Η>'I���������Ǧ]ď<�^~��gpO}�ꃏ���{/����ݯ�������V��n���{������?x�ͷ>��߽qz~���_==>��?�y�c��g�~��g?��믿�ߛo����o{x��R��t��G?����ɦ�՞��ꆸ̊j�B����J�o]E�l�K�b�"���J�??�&��y.�a�f��ˣ]դ)M�39ҿ��o��Ї~��}[�����'5Li�&!�����Z�t����jH��K��!k4�4���mw��HA�)b$b\~��޽��=�s���ٕ/V8~�m�_x�h�{���R��72��~H��4����dI��2��/�G�|�R��[�h8՝��Fv]��j��7�|Hx��p������qX�+�D� K�%�����{���)s,��Y�,�Z^H/fY�ʒh��u����i�PU��v�#Ѩ�(Ԟ� �7�g-�K�TY| ��ٔ�P"B*+aڹ�Q�u�sp0E��f:�W�8>^��KBt�a��`�F!�6JJ�i	�^�s�H�$�)� ��ǔ�nǈ��[n���i'�F�P>�d!�'W��@"ׅ��FYF&k
�Ee�O�Z�m�($h
�����0��������v�U�R�.�ql~L��ہRdI�JlRR8Ǻn	B���Qfϖ�P�lǩ�k�K/����_r0)L-�;��!r_��;��;�.M�%L#MS�pL�8��h#������� 8���pL��$bd�N���F�ͷWpkD�Z��ǘ��ͤ�G��q��;^N���}V��@>�(�A�>M #LsuB� $k��T�lSY�I6����)AJȨ
B��9t���їh]R�HH�*eqL������P Ҵ
#ӏ\F
�Hm@DM�д޼^Z"�VH!�O��)Z�3r��D���i�r�����r���e*�����
1J7�l4m9��(�X
&��9�9�L863���9YQ4�*�����z3͏P!#��U���1#W�N���j��)'�\�����P-
�	���(j�)�}L�jE[�p{(�v��頙R3�L�n��0�l�ߴ=��j�F�'�O�S��	�l�k�V���)���V(�R�8��t>�(rLx�N3Q��*�ij�AV'�:LMH]cHJ;it�G�hJ��#�
�q�D8�����RQ>)�������%KLTȑ� 9�1��4�:G
�M3�!K����D.�_KIQ(J�~8)!�P�:D�� 	�>�#�$'��AF��L�T4��N�|��G��~DPn1M�f��*��	k����9��)��+G���p�*��i�����3
�
����z��6Ѯ�t�M�i�1����jʥ���[j�^���ş�)̪��rF��4V:؊�v>A�������8���C�
���ҵͯt!4�7��w����Hd|���8�	��j�K�7n�(i�����l���B���Eq�!8S}h��1Z�tf�#Lj�:+8SW(�!@���Y���9��jr8�!9�S0B��ȑ��!S�zf5�)k�!	�b��M%v�0kO.�L.��9X�R�8��^�Vјu�<�IU�%�25C����'�~�B�����tdS���9-��� !%BL~>�ZJ�\��E�cF.�60�2��N:�R���\W>�I�Ϗ�O�����������,-�ɭ��s��Uݢ�e�scә�i
q���X��B�;���@@8J�O,B!�~*d*D��P:!�a�8�*%&^��m�iQ阦pۅ��\���@YU1���U3�;lMʮ+4S�|��MO���>r��h�5��K_/��r8v^�]��,?;I_�}�s�hwu��0.ˇ;}��p�w�vQ:�Y-K��Z�����aGm|4������Y�^��Y��Iܾr�s����'WON϶���=�/W�1u�CP���wޞ\]�.��v��n��������OGo9=�c�+k�b�����R�=�]֛��T��u��>��=�{���'ث{����-�ק>�����W��J�O|���H����˷�J_n%S�)���m��ˋ��	���f�Vw!�UgiG�?p�w��+RY�v�/��x"��YV�������C>���w��ջw���^��|�����;������V_���W^���~����O�8�88=����Ǐ����������)Y�s�ק�j�M[�)ـ��>��F�u�pDВk�,��G����\��8h���7��2��F�C�r�j �Uc�	�L��>���VԴ6�0m�0�'�B�M3�!8�p��*�"��5i^s��@>5����x��Íֹ��7�B�8�����r,Ĉ� _���%�1i�L�B��g�W'��n���!�_�$'�T����cd�?�'RQN>���T���д���������΁����x^q����ǿ��w?��Ͼ�����=�ڿ<?yt��?���_��g._=���m[�˝���K�}t����N�מּ��\�]�n�zoߣ�7�|���q��Jk�Mg��m��W_}�SCh4��1�`4�{��-ƨyxk���)T�u�Ϙ�8�-8�u���t������{�D�wq4��/W�;������▆���n�SX����ۦ�%TRH� �*�WN+� �1ZY)ԙ�\��UQhI�4M��,��S
޳4:e���(�����_V�:��;8?��?����ٯ?��׿� �̟�^�'ݽ6���F�)�j�>��"�u����Ԕ� � �o���|�:��>܈#�3�>�8S���L�o�8�q,�`#��\��Ƴ�jI����(qօ *�H߆��GN#石ӹ��ڹ��ژ,��i�&��(d"��ݐ���z0J'��e%�0��v��OSn4� �1;��!�����L�&�b�9)���s�L_u��L:�NPLW|8�)�
�����Ɨ��A�+
dT��� r)pllY�|:�5��"h�&�L����/%7Z�8���jʨ�3�u�� W%P�Ȝ�%YPS�z��B�'%Z�4�il�3Ө�T�GKV!FH=R�OE��0��pj��I�τ�"K��k���C? ����9��J =�d���(������� ~���+�m�#ԊZ��%�&�|4�B@�&9?B)1�	~�(3�u$;R5�PѦ�b��,�B�����U,Ե!0H��)Ǳ�Y�� #s<�����8FQd{�o!냼<^UKԈ`t���;@���FИ����g!���A�GC椣4\��+L��C����#�O�_�i��Xlp��I���	'˪nD`i�9F���LJ�Y�L�YTH�I�if�"%#�*�6�L!��uUö�5���i��p��J:��|�� �?:|Y���D8�M!-f/��¬N4�BJG��Ø�}��1:�F-G9gs�@��69u�DS�Ө��	��U�fZb~4��D�4��>������֫�Df�6�i�^�uM�L�ҳÐp����c��WZ�^,�}VW@��Aa��8FQ�7��_�ܖ���J2f�r�p����Q?�j���_J��ӘS��d�	秖�g���8�

��Rc��)�v-A�!�零'��'�:��]���AȏɯUL����'b9��	)�A��@L���B�jY��ґ9�*'�a�*"Xb��U���[))S�UQ�!X�vL3���%}
��)��3R�h�qZ���U���(���l���򴁌����*j�n��Nx�ն���&E��S2N>|�-��P��ih�)�RD+�N���\Și�Ѥ�B"�Ưg>G.�'�)�I�#���D�!<$�� vΔ�Y	S�6,_zSBx4����Sc�p�2��#�>�$}'0�(���qt���I��ʊVV�Ǆ����yڔ�a�d���8p��k�g�B-D�!�p�S+Ett&
,JJ.�fL�7�8'D���$�r���*e�    IDAT8�zJ�����E0P4�ֵd�s��g�pJW%�%0�(D�)�1����k��w�8�˭�q�U'UQ�D�덎s�}��6�#���4���c��E�#ki��r�dI['Z���B��O3��G���V�\#�eƉ,q��X]㗎5A淼�����z0N�ͮr����8M����9V�9
@�RL���_��o����ږh�r�@�qZc몙@8�N�mh2�'��S�e�˧	/�=4\V����c^\�v<��z\����'y��u���o._8�����n�W����3IU\>���Y�|��5��-�8N;W;ˇ����0�ӧ���v�Ã����=\�����90�������m=zz��n}k�/���N���c�R�>_���ul�^���������\��b}���������u��v���1�w9�7˧B9[��ڣ��?w���ի��z�I�����g�˃𻫣'W�Ҷa�>�8���[x���R���U�]B�����,Bs|�6�rC���w%Y��Wow�ݐǁ����/�a8��?~���;{/�|���;�7;:7W'�����=�7�����z����O��������?�yv�0O�}�0}ʚ�W]�uT�r����)tk�)p�#H�e-�\����Bc��c2
�^�B�~io�^bՓJV"�"2U(����R��NˤSK�`&ȩ43���5����
	�E�h���*�
2��Y����;�gZb���$���I�9��m�-�X�t%}V��0YjA���+aZ�,N��zYdRƤb��
� e!Íp��J��ϙnsf��/�fRF6R8�BUѡ(D�l�29��A����7;�}W����O���÷�e������[O���O~�/�ɇ��H���_�����K/}����K>���'��}��ܽÝ�w��]��>}p�b�.�B��g|:׀�c���QGV��������������Ehn�j^��(�[��g�抔,N��Rk�Wȇ�Af������Ȝ�F])D\T3q�t=4R��q����w��ַ����|g�J�9�F<��|@BCL��k�^����8B��T7��%��9����C�W&��r}W�����|D?9���G�Ͻxpxq|���w�?~�ѯ>����;�������S�����o�)�*d�<���g6d:oO�8ȢFӎS}��8� �_���t`QSN|4�R� l��l`H�@LK�esgY�Xk,Ck��>:�C�~ KD��r�l�l6c��[4�����'E���2���s�'�pf]�r:����?�����_����s)�l��1��ɩ��3Z|�"����)�mw�p(8�R��2�Zb��e|d�I\]��u>��c6U(��HE��mLOp;
)�R4L��	!j���
�Q�&%0׍?�t���Zi��"Q'Z��)�uUSHWME��X��*�&�1���2�˒n�@�GY1!j�t͘�@K�P��a#��+![��&X
9[�`]][��am~��8Լ��Z*QA���}�$�oډ�ܳ�J���������k�=ԡ�
y9�7����|]�w���p�d��GD3�"�	�5�Ʒ�tp��"q�m��˥,�qm�!R$��0�2� �btD�!�αjE�u�
�!���#W�6�F!��h�+��w�l;�a����!�Uɩ�N��>8�(��R��I��O6AdY�����Hտs���k S�I�!�l�v���U
�J%M5
Ff*��G��J�o����Y��*=�����֕)���JB$�d��G�#�ե0�)_
G�Zh�J���ޖ��Tx"F����,_��̎#r���_:�i���g5�_
P?��X?�8�2��[�d���3�q�pXj��S��v��B��ÓŇ������HM��~bvv!T�H&TJ����M�*Ѵ�S���ϙ��[3��8���|��4�v"h]��q��YM&�/gҁY��EM��FߔH��FF�[Q#��ĩO"�,���΢p��L��4�)&�q�*���K�0!YƑ��1$�)�l++ķ"�F�a�F��o6ˍl�R16�o����E�Q`��}:p�n�,��@R�!�vI��h��c��l,$��6����i�o�#�Ϛv\��^�ru�4���!�`�O�� L�΁+��ԒD�����d%nZ"K��eA��Q��8L�關��P����}�!&+M�*����R��ܶ�T]�v��B��q�$�ÇG�a�/�M� G���Dڴh�cY�/1Gd�	'"��(�4r��V�4�6�%�"ԩ�ե��A�\Ru�X��9ps��R�˙��d��D����d�MSo��	·�F4Y�-s4�^"~f+*�8k7%R�1[�&B����9}��	Ռ)<N�ZH�3�����"���čR"řÑR?��J2j�H)�PmTBʈ��aL
��|����9�,��Ցsj��ᯉ����BUI���|����of��4@$٩E�E�v����隵�;�S��C���C���L΁����D:ƩR���1�J��^�p��y���?�������������ۿ�;]d4�hz��p��'D��_	MeeU�kp�*��㈚J���;�tL���Ás�tS�~5���Ց�~�`�"Y�02�y��t��0���yK.Ӄ:�Y�C��JS�W�Z��ΥOR.��gv{�Zէ|���,�w6}Xh��n۾��g"=��D���埯�����Ƭߍ�}Ic�̝Վ_�.}�춿��l�<R�ݺZ.zJYyjO��|�b���؂woV{�9�>{y�#(�>Q�s�'�Pn��7�����N}��g�|B��̽뵟>�i���:==q���SR�呦��Z�|���Y��ܧ~��[oܿ��̯?�Ⴛf�=�J�y�!��ѝ��z���ڵ6�ùg�ˏ.4V;>�j�ly��hcف�)g��FX�ׯ g����㑃��Ζ~��Q�' ���P�II_��_�{����d��;�>��}�|�Q8������ӛ-:g��w|��ON��~��ݻ�W��I�sO�>Z��9�x�Qq�:���9*m!cB�'�NL��z��g*1��0���B���K�`��T�[r�3䘛#r�0�U4���VK��o~�B����i�	���·UGPB���GD(Y!WS���8Å�t�Fz
�켐�l)p�I��4�>e���"�4=GH���T.5~Yu"wSH�䔒N8��M��K�Lϣ@�*�mT�|��h!���?V����0Y�N�h:ƜSVΧ��n�Y���G��T�~S�� ���?��?�n��ǧ���}��z��l����o_^}v��u��Ó_ry��O<� 9@ƿ�gR�ݿ��W_;����ǧw�?<>;}�����?x���������n�*�ζk���3���K/����ozX�g]����nK��������o��72�"w��h�*l]���.�e� �9MМ'�DXgo�*p|��;��NHAd"	vU���~�gL%Z��bv�7Hɽ�jZ�^;T�S�����J�`�|8�3x���E�dI�
������������n�Z���m���8��<Ǐ/��������k/���7�����Ǟ,�-����ZhV���ѿ�r)�Ĵ9ִ̞�����.Kch�b4�(�L��*��nW��d��(~��̴%ꁩ�l�c�s����9ka�reՆ��5�3Y�c������I�Oي졿��ڡ�*�8�мm�a�NVO�U��H��?��?��?�o
|�{ｗ�ס�U��P��$�*)%t��nmY����Hr�\�ꢤ �W�5�r?>_:)�xS�����(��U�l�t%K!��*&�r!��pY����t>Y�@A]�+�D[���(� �0�!��.j��Vat�����B�>�N��i�RW }-խ)��2M��kSf�w8�Rh�#T!d
�1Y��0#2�,�4f�
YHk���$K�(��a�����	E���3��H�q���)�����h�>�ДB/��o���L=��BȚ�s%�4�|6�>k��zh�ʲvLQ#�V*�o�`*��2�iѲJ��W��~S)u'}S{��5>DV=s��ۈo���!혫q�&��B�2��e�q���Ls��8fK02��"PƄr�곊�E��D|��8G'fH�2f4SedRN>5� ����.�A������Ѵ�a� ��$� �W��cB�%ڄ�v�T�>�)4�Dho��d��1!|7�U�S�89��6EG|4���ht�b���@�Y#ZUB�������L!�i��-��F:mZU1���[8ddkH�B! ����L��2�uq�|`�R +2:�X�EcF�G�Dk��`m&UKK4����Af
��Iөˁ[Q ��:�{QL!��<H/E�U�c'B���*�$U?��M9�m�ֹ�9��@]U���)DV��j��j����D~��D�	�� ?3�c|�Q�Z�)%��b ܔߴ5�W��21�sd�K��&�S�C�;��,�v� D��UIa�(ш�������M��R�� ��7H�U�F���%rj���p�5LysCD7u��u��W�� ␍�(��/D3B/�`R8�d	%�{���8�Z���n���Tbx�0f:����Ʃ���S($K3�7Mj�XW��Pk!�0��FG��6r�	��Y���|V�Hd-���H[!4k�3���Ҵ� kե
��}{@󍵍��7v�)�
/Tthu����9����Μ���:�U�,��1I�B6�^�tp
�'����5 ����)��I��[f�)�u.%�B��h�a:q^	�����Ԅ�U��i-	��2�:R�h��o��_�D0��L
�$���M�a���9$><2�T{�0eUt�Y��S�t!���eZ�T?���DS��'�؏pe����@S�r�66�g���Y�ʏS�!~��=�:� �XN"�pc��L��Ʃ甥p�_N�7�u�UM�W"_H36ʔ��i!�r�>6�� �A�kW�6E�8m�hB�G�PK|�=�����������$1��� ��]�Ht��\�VG����f�)~�������U}��B�$���_���Ӥf�D��OS�hu�Bt8:��:��L0"'�A�kR9
�V��Q��C@�z�e�/.1=����ɝE�|lq�%G����Q�k�t��=v�}W�.����[��^�.>�փϛ�e疃��������������=�������h�Y=Z�v���j�`��w��<�9_�$��o�������n.=}�M��u�[7�z�76}sY����͍�t��t�>:�Eߵ�TԲ�X�D�o�>��)�9��M���[�O>��������׷W���גǸ��ѝ�#߸�á��.ρ�-�;��Z�n�ew�����n�?7�O!nԱ�X�������.���K����8���ԡt��g9���9!����d���������w>��<�}���w���{�3{��c_���������ǎ���������{t����r:��qR�1ֳ��i��EE���g�Ԟ��R�ӇG��'���!?����]1�J))Ob�S rj�K���h���gӕ�7�@kF�5|~א�"��d��wM0�r�*F��I�]BP�Nr@c]@j���GEN�(�ll��W�T#�fJ��M1'�NY��~L��8p�|"��^QL��i8̺OYd�icd�J�Ӊ�O��3`Y�l��hm��b7l���|���O=��7j��l-:�����ӧ�����V�����j�-Xs�/������[�w�=}��?<|�h��������������ӳ��ý�%�:w;T��@>��C��Yz7�Mzv �񁩐g]�8�[s{����1;� Ȣ��`,"g�|>�F�[�#��*�MW0�lz�K�Gur-��\IIXEM@�#G�i�i��t��5��-�_�����cd�r=��g�iU=z��._#��_�1�ɛ���?�n�������~|��ݏ�����:{���ۜ՝Õ/�M	^{���ʿ���tVmy㼹޽{w����@����?���=��[�X7����X=�RL��98-��#�0	�V́�0<ǈl�-��᪘�J����!�wD�Xu��5����KF>qSL�8x#r��׾q��g�,�sSg��L?z��2�����^m����?������޿1����ȵd8S#�̼Ɩ3a���~t�Rk�V,�/ˋ�W>���Rj��:$h�oߐ5c�A
��l{e�JY,��(�s)L���J�H��7�R�K�s@-�q��� ���B�Y-U$&�fJ�I4�5�O�|��,A!��>!M)�2%�Dǁ�.�pc��.a�?����i4�gBF"u"�S3ќ̎H|�d'�>�!�A'��/J��M3J�)W����,�hG�A�(�2&Y��N~���|���}�W��*�r[��������&$Q�*�"��TV���o�uK��hi�:��Z)23U���ǡ����9#Ĕ�QE�)�Ңed��$��>))m���ÉL�����h-!���pm>�U"�U4�p�^�zӒ,R�� Ku�����!��Z7�+L��e�Y�R��Y-��6���_"�>���ej��hR������^an{^��s�9\�_~�e?Q���"��0g�v�)7�UA`1�Y��A�/Z�SeFYpQN��"�e��i�nD(��NN���\�F��ji��*D�(Ytq
�#�o���V3D��Ʀ(�i8�m�A�}�>f�jL9Gn�3֏Q�h�/�ֵ��ҟ�M�p���:!N�3"Պ��*��#Y{A��z���V��Z瀔M�4��H��@ G3
��>�yD�
��CS�>�2(�?�(�a����8�(�-�u#\J{"D����)�2�4C�*�Bc���(O"�	1"ą�)_�4�4MSt�dF(��O�։r BU�x����o��C�:?���$�ӑ�|dS��o�j&�X�eF�O��"B{���pX�DL7��`�k�>k9�-d*�)���&Dд��pS���Ҧ#���(��� �I�ϩ�PӤ�B�1�C�b�ǬH���&_�4���?�')N)h1�k �)`>| ��a��t��҄��\F��FC�`Jb:Hxʲ�hF+
ᗢ��LME�D��� B�F:�t�Ң$V�2�rƢ������t���U��ҁ5 ����d�ɩI>���T����aJ�E�Lk��\S`0�>��PMb��5�hU09�,4���6�"��
Ǵ���4�)�*�7qdE��i�
L��R+�B:��rSL~��jڪK�d�L���)�TH��.����b��p|�ҍ��ժ�|�Z��1�J�IΉ�H�r�&���B�r��a�Y% �����9Q��R�f3ф\ ��M?��簺-jl�*&�«�>�f��Ii8�aʊ�X	��l�6�*d��9��,f�j*X�%R0�LjI[3볐1��p��)��7���J����Ӈ0Sx�F�~Mvߣ;No��V �Z{9mf��������z��#��Y��)�n ���{E8(,>����/���"�#�+?�,���B�>�� p���u��[~�~��	���L�%�GR;��y��܎g�>�x�l��]>��Y���L��CM�;�<���vz�y�Z�����og]>ȸ<����65xu�#�[OND/�������ݚ�9^Dt���K�p�ʯ�K�m�k�H�>�y�cJ�r����c��3������y���[��zk��fo����P[�'/G�q����8?�AQw�?��w�
�`��\^�]n�-oѻG7W���S���J�x�W�CP8�/�="v�ދ�_y��>\�6��s�����f�����X��C��w~`G��,���|j�W&:ܸs��,�Y�R0;8n�_�����,����'����������͗�����1ؓ�˓��?��_�����G���������ؾ�˫n|H���G������-����j    IDAT�~Q�C�/cm/���B6-�?Q�E5PJ`+�7�:'E)�%j��S��ҏ��<I��SL��U�@TI!���Y��f�l"8R�Y阁�q�k�o!�E�MG�cJӫޒq�����)�z���is��H��Vm�����B����j���,�h5P?5F�A��rd�ɇ	FI���-D*5��.��2g�ҩUR���8Ղ�ۻ�iVu;]�[�Ѭ\�r�M�5�/es��i�hL���?�p�,�F�B���ӟ:R>k~qr�&�����?>9>{r��/{Ǉ{G>�~}gu�������ٹK���{e_�M�7o����o��ж?����GO�����O����[��H��<���_��_���/�!��/4[�m�E�7���w��K4�����)ԣKC�ޞ���(uu�L�i���܆�'�Fjp���H��z8/}bB���ҽ���� 5����P�
�P�43%��ySW�hL� �qB�:��|�Uэ���>$G:����$�tI�� ˟������O%�l��7B�;�[{7�����k/�������������>z�{������9?j��KGGGޟo�%k�v�|M�������x���}#��_��?��;�G�|l�q����� �Bۅ�a!֕ӈ&+�r�o��13�[w���V�ڞ�p�gF{X��1
F%��02�6B:�hʅ���@���*��G��N��+�����+��ǔ)��艎����O�����sd4����$T�Q�r:a���	jX{DZ��uJ��9�1��ʈ́4�����d�ۦ�-�5b�(Z�:��\��PE��0R rb��@F?q4`+���q�\.k/�i�)<Z�SN��L�ń���L)[�X:�R�,���,
�T��f�8F&�HS�P����N=�i�t|�5r�N!V'�a��m{�S|��Ȳ
�#�)]T(q�1�uV�gZ���E�;����=Q�Ȳ���D-Y��������*ȭW�|4g,��n�:�� �I�uFMΦM��sf�� ې�8��	����%� �U�es�ئ�*�=���}���:i�)�`$��>5S#B�b�3�w5_��[o����c*žA�oW]L��֭#g8n��W�k�_44 i{��o���p����QRD�I��V��"�8ƺZ+,CE]�:�i�%�Y6n-�nt8�f6~�Fc���%���]�����{�Џ6��X>Yg�n� 6jJ�`�q��6e�UŴ�ï(R|CfM�K�ş���"ʑވ��v)��ߪ9tb�R��vt*aʱ��Cֽ=[v]w?���d�bَcIV�mLBQI�TQTx���W����%�E���$$�$H�Y��|�d��������vufu��7~�7Ɯk��^k_�Z��q:���ք�0�7�^�(�0p�8�6 BG�Ys͚@Z홼��K�Y#Cg!��~�^�0�Ė(2�]���\��`���/��@!h��0�B��bl9墚Q��@���p=YC�Z��t�G��u+jī_Op�7�6�4=L �y�;�@4���_8Z5cri8���psޭ'�&����Q&[HQf���汐,mtDU�b�	6)�J*�^C�r��N�t4��\2���0-_c��]j�\h�'P#���*[vs����D�dL<�DD��%��/�L$�^K�K�a�f��ƥ)IOS��4�x
�Ԓճy[C���;�o��Hq�f�o
)$UDUm6W{�,����g�g�E�^����S������4Qb�4�B4|
-i����a��6�e�ak�(�+�� 0���!+�!�~:M�𫐋�ؼ�r�zj8ɦ@����$���+��x��C���#����,*}�a)�TK�Ϩ~vS(�a3�M!o��8��lFx=Py�jcDXEl���b��i�0�0���@�h�f�s?���q�[
ޢ,C�)�k����0�8��n�'��K�[8�-�
�,�\
�E����&�3��Nm��i��e/�B ~jz����Q�b�C�24�a�1	F�WL)�!Z3E�HxC�f� o�zM<Wj� g[��S6D&�	IP�.K ;�@|+PȈ���/W�4'i�>B��B�R�2�WdTXI��l�R�L�������>N|}�t�4y���&��'�>4F������;�|�����5r���g��bt!eh����b@��4=:�pׅ{u�6��b0�@��
q0�C�.p M��(��/�m)�k�l�����H�^��"hU�H�kk+�ۨϟ��Jq��MJ�P���_�P��PuI��<�.�M�U����݆9qK�딾�ʶ��U���_.�c��g]";���I�vi�'x�����~ẫ{����~���Jzq�i����������몴ۆ�'n�wq~E�U6rr�2WS�)�������V�>�*�öݺ���{m�}�������ý��_~~}y�^��<�~r{�[�o<|�����W^~�����s���V�����׶ӡ�ų��ɺ�5�C=���M��!p��v1G3�^�c�9vh����
]��My;!��ŅK�������?����w�ҧr����'�G��?��o�/~�u����T����Q:Ÿ��#E%�
S�,�ڼ��t*�bk�z
���z�@�\�!�2_6ph��*��\_"�f�hN:������Ur���&�D�	�DQ�<�-ۚl�)�ћr6�XC�����yۇ+0������@G��\s-ёB�+��r^j�IF
s� ;�ư�jp|L�N}|.dHe�!�y�"�M���z�l��.Y�m �E�.N��8�rQ��B�Fb�1�q �!��DA ��K�Nv�O��5Q�ȨO�!�!�w�Ñ2��l�ʠ��*��/�����'n�����>��������i{��u�G�C�;�ϒ��6W����n�%���Ds�Ʈs�CS�2���=��AI�<�j]���'R�޼R@�ͺű�(���7�Y=rA�%V�R���4.���w��6_�g^�f�4׎�BcV��HW���"����4Cήn�!}�)8��A�4&ЃM_�T:��e�}�RI~{o�+�>���y���ó���ٿ�w��_���/��_�������{�������]��78��f��_q���-HG�{.�Z|Kw��+|�gۛG/�z&S���#�b،R�֛�E���P�Ĭ;5D�[
�L�����#A÷b�쎎!��3Dfk��dL����_��\v��y�b�����x��I�.���]���!l�x��y �x~P�#��x��2[�{���/���w3)�����)�EF�NUͅ�;S����$�BC����4�АEA(�i�� �h^��D�WPC�3B���h�Zk���K�/�w�sY(Q��t�L���i�E�Vp�+�SN���վ�G�[�#X%6��(�� !�15�lL-MxE�j�(�����G�#����,��r���������W��t�D���+�B��ew\0y�P��$*��+�|�M
8Y�����C��"���_
��"Ś����� �/�7AtxS��b��l����N� \!	�+C�U#)L��&�+0D�������#R=�J?~�h��\)��N�x-�%է�S;�#¡�ܯ`��1��.CL�5k�1R�֜�!W'��wy{mw��/��pp�Q���x�S�&PT�z5�:��
á���q��x=*���1��lm66ٌ�z�(K�-��D5Ma�!�GVC ��&[_�9
=��->���A6��3$�@dF��ʶ&����Ր���w�� �8M\T�\5'��8@��Xv}����Hq,���.;CC�S�W��fI�w+o��ky�Q,[C�#d�φ�0����C�l���%W���ƌ���siS�p�j��3
�t���ް�ak�+/o�aӁc��iV'#���Ç��d�UR8�V����q$�g� �˰�c�űfh͔!G8CC�J�g�8��-�n�ū�L0N����\�\�S+�>e�f�sd˂��L �����٘��>N�R��UIӷnf*E�7/��K�]m�MNPI����_���쁐*O?УUlR��s&�`d���ؼ�Mm
�@3��g;��d��!!_��a�K��,��)$R`�"J������@6C�0ᆚ!/C��k���N��#�V���\-�(.Q��#OY,���h��(E�B����٩�@��UvL� 1�&�[8��T6A6^��i"�Sxe��xȮx卬zت��6L��DkX@!8�eA�	/��^��S�BrA��5LM%�賓���i�(�tүo��2j���?C�zda�i\3�n�4�
��BE
a���تm�G#������Po C"k8zH"ك��v�R`� Jé��ڱ���E�р��̰
�B�;՗eR7D� �fdÌ�`k!��Aj��b�2:X3��&�MՌ�R��@�[_t��b��͐kV&v
�UH�W�!r����Z��e�t��0^��fJ<�X|xKĨ�1�G�R��
#���k��+ ~6�7��=�蔥�k1EbU�!������Eqi�!!�ևWʒ�[y�S��&��	B�M���@聘��ү ���> [�ׄ#$R
��8pt@;
�
Dfǡ#$M��OzQ�֯e�){����f[^w(U���w�r�=N�p��_�����Kվ�}�keݥ�.b��wx}ẼK�n$����G��;�>�iQ���ܸ�sd������_����9˅�wC��?8{�~�Ӈ6���n�]�=�n�[�Ow�m�6bM[v�w������oY�q�e�h��7_z��W�����w*t^��[z�}�dݢ��UW�}
�����~�8�O��__]�H:�q����zYTba�tkcK�Y^�=��~P�{l�vМfy�㰘�kv|��K$�va�gp�5�bs�kKt�d�.=:񉝓��_��?��'?��G�=���?���)+L�1�U\��>�^#���5�Vu�o	
Vۮ��O�т�Z �Xry�,��d��]/��m7�aUQC+�@6&��@C6����KsR+�
#3�����g���pQ��D5DH
�GII	t�]�d���F��C��WĹ:�9L�t �uЫ�9�<�b��X�
^�[Y�m�QC"���o�
�Q�t��a;�9���0����3�Z��>ʁ�bwC�v�����5�wKr�H�V�x�!���k/1�i�����Z(Y��̈���v��=g%"��̅�����������7"��J����O~��߾���O�<�-~.�����2:�d��ݖ}C����ֲ=��4;DR�ՠ������~��|v�>�uT��Aav��V���W��K����4-N^`�ְ�KͶW�"�� �Jr�t��W�Z|54)e�쑓�i���b�2���&Wa�Pqu�k�Z����Y�*V�Rh��&B�Xd �X:��w�ᡏ�`�+7�X_�~r}vst�����]>z����_|�ރ����?��粵����yݻ�`zz������C?���������ř7���V=xx�bzz89:�]��J�(Uve+�	;�!jV0[C��oK4�#����:�pج�-D��蔋*��7<p�S��&E"ӌV"�h�=�e)����A�%�=`�"���I�t��" fg[�G��E嬊��kkZyYxۻ����|�l�lȚ۶��M`PR�)�����P%��5d�=m$�Z���x�z����A�R���T�auBx�h�b�2,\aD��+��`ȖԚ粆��!��.E�I�����/���T�"�q�Dֳj'A $A��E�����eX�U��o_\��08���@ۉ��;�!��>������գ�$Nn�Ś�()R��$\���N
����H�����u�J�����Gp���C.c�������ft��ѡ*�
ۢ)C=�����h��i!�f��K
�I�jH���r!s��iR!Z�M�tzƬ�YTd)�eIM�,�p͂�;ke��8&/��Ny:
�G�ڎ�ٰ�k\[��eg�\�eQ�7~z��e��Izs�w�f�u���Ԋ�l�DNA2�1�v#BY�(U�b�gQ���Dx� ��j�!����g,�͆ d��)�"�]���obij��bed�!�7���VF�Dp2�Z�bKX

��e��ږ��$bd��Zi��E!�D����
���,�n��P�i�EQw�0��1����SIᆅ�P�z����PLuN�B�Φ��sW��r�f'<d
��Cʎ�����]�zC�JpD	���e�TS_" �!�|{�J�©N�f�10�!84�F���
���Bp��ep�gsR�M�%[o57�-l�)AH-b8RD���154C����%^��ƦYHs7�(Df�L���~4�V#W|��āl|��(����b(D����l-�r��������>�a�g	mG��Zvy����T��!��HA��0B+_��:e^-����t����ÞY��_�tx�"e��DH���#�� k��62D`j���)WdQ�q�ԚoȮ8<P�ƗhR�=�NV޲4/^-<��d4ǆB�a��]CA���
l�l���Xx����\�
@��K#��l��pd���X!@��)�DՀ���E1�ʀ3�p��gWۊ�8�e�a)�������r�g�4�* ��NI5j�Ҝ�c�ALC����Ϙ]>�Uj�PI����D��
��`�+���|ަY���-H|H�*�X�@=�px�d��,v�Rs�5/�l"��+r�D.��9�"h8!��[��Ga!SC,eR�F5�4��X�YLy�>�QK�p.�e�������d�$�X^�/	B�-�(�R���X/�f��;�
x�aV�jք���'�@N�`�C�l(�'�)o��J��Ѧ<^C�^x�2��ҥ��'�N�iVҸfX:x��Pǐ8Cv�0�!�.J�Ud���l�&5IK�HQ=Rp�Z�ʴ%���ro��zg�@�&����v�6)舊φ�+f����B��v5�����^ٱ+�����P\�Ȇ�<�b*���:f]�"�QC�"� �ýu�r���D{���֝�\�<i�|��%P��姼��b����m/_�d��^ޭ�\�lӮ\����zIA�S飼�7Ⱥ�y�q�f��H��X�5���ۜ^؞���������܎���uO����{g�=qm���Ǻ��Ki�+g۵���/߻��ɔut K����YV�8��J�������]?��믽�կ=x��/|����.���{�kw�nO��ǿ��O��	]_l'+߈붡�/�U�soG��!��X5l{��r.G�:�^�/���#��i=��-f��]�r;kme�e@��o�o��yz�؇F�ו��C��1�+֚�ܸ�!�(�UEY�4��f�P- �/V��|{�$����z_��U�R@�\�����X{oK�ք�gJ��N�v���l�.�m�Ǥ�m���m�*��hf4KT��+M�`"A߂w�����EB���q��.c�T��V$�&���@��0#6�!v���l�����#P8�F��t@'YDH��aDk�����J��0���
o��Gh��iR� �[��C+��tԠ��\`}vC���Z$h��pL��@j�l^�@���O��9}.�V�C���>.ׂ[v5�NNo��Q�Qs([�b_<y�~%�o}��&"����v�� ���6��O)x]Xv������fLv�%���� �,rۣ\ҵ8�$��ok���bIA4�@�hl}�u"�2�j�))�2L�#�����=O*�mM�cC�f��rЂC*��T_���������E�4�PEKT�>[ ۂ":e��t�	�t�}��߼v�=���G��j���_�����k������v��?��O�����[�c1������������]{�S�~9��S�����{WG�?�{x�����>��C��7t}�.d+����uo�l屹Z��	o�z6�^�l�؄7�f�c�L�T^}k�."�=�`�2:iR`=n    IDAT�k8Cj�����,�\z�51��NR�2��z��m;sQX���ܛ���6��G��8/M�!7{lEW�,�m����㟲ư\mkY�'Q�Qyi��7�M��d��具�\�qC�=�Q[�S���qkp�S���c6���UI��@=���EPS�!Ӛ �Ѭ^���ri�#v�è�b!�1KW޼즐Yٖ�S&Mex�f @�P�[��$2��t2&�>B!�L����*�T���5�VU!����Av^j͔�4^"�@RN�\�dx��,[��g����x!��������������ȦU�]�>%�m��S?RlX4j��SC�&�-)���A%!�B�jq�ZHކcg��Š6^�;�4�c�!èM�I�B�"�5C"Z��*���b�
�pkk��[(O�V�I�.5��B�a:Y�l��מa8o�"�Q�C�~;@�o��^/¶Wt�5k��	ֻ=׌���<=�6��5"�%*�	��M���dM��,0);��~p������m��!�I� �c5�V��aj\8p�R+���qd�W'��
U�p��+x;�h\��KDA8P{�ĔzSZ�MH`�tb��ǔ�0���2f.��e�J$j�P�#� ��B��$K:�.�"���^���B�A�<5�5�d�M�8��q��F�n���ɫ�d�
��Te�7Ô�A�Vm��Aֆ�&�G���jf:�U8!E�se��&���nؤ�Q!A�V6CC���Mа� �r�B��&��f��{��Z�ķB�j�hD��!c�\p) �N^�:������㧖�>��l=2p��b8\��R��t  ����dd��S�,l.-�ݾ%���Bn��y˨�2æ���H��M::B�MͰ���ĒҐ�T����R� z�yFRd=����O�@x��i�KDS.��:�h�5H`C.�t��w]�:�Z�� �W��zv��05�Xa965�q,�Z.LF6�^-��@+�pв�^C�c$�Ej�z�G_=c3p�,We���N6�~V�rXx.�!�IA��/c+�Clކ%5�f2�eak�h� 0��D�#���	���B�j��Y��-#��E輔f��4!��l�6��ř�16�e��dD�(�j�їפ�1�?�F��YS j�V�!΅��n�5dPfg�����	�7YC�z��e��GP����WI�!$�@K��a [�fC�Yy3k�D�e-2��p D��F_|Y�-5/\����?B�>5F.��S
R�D�	�p(��X)�3D��
Ԓ&�Q�cM�G�\���#������
�[9o��V ��^��q���pF�p�!�њT���!�
�����]HU��G�m����pM��ͫYCK�Xx�U�D4L�zL}��:R���aQ@���B2�-{�;�Zt�ȫN���˺���<��[�`ij˞�����f7���-W׵�Ua�ķp/v����mh���~�e~n����߉�̥ �OR^_�W�8o�����w��g.}8�����z�{}�wX����\�1�5��d�@�h!�"�����������#;�U���뛓#?��e�w?���GW^8<9���;���}?���n&�F=�]�{�CZb&����,�����n��\=9���s�����_������腗>���>�����L��ž+k�����?�urt�� o|��Z�#�ȃ�[��Nk�Wk�0�:4]��D�e�uj\�o|������?.7�Ή�������:"��hWG�C�X�w� ���b)��<9�8��z����=?����/>��/�qgK6jUY%"N�n[0����Z�� W.^F�~쭘�i�-��jb�e�C4��n:)�*�(��	"[�j+iY�!���\E�=��c ��HYI�Z
Ț��<w�f]����A�:F."uI�!�ZN�k��"!��X�K�rV��E.q��)_�QfW d� �e1׻�"�Ͻ)o�ibU^
F�4��"�r%�����/�t����*��
��gH�W��eL�* �p��x����1�Bd�
���Mv!��24�4��D̎��Ԓ��7��6��#C������DS��}�W�ܷ���}GG���6�+����6���K��� Ȁ��)[ml�lg!�������*Q��v��!��ADm��Q��&+�l� >������M.*CRm�pa*��^��� B�`1��ض����7�x�7~�7�\����t�Y�l�Q�^����z����7~�`��S�D�� _�5Od�P���������$�k��}d���s���z������hr�;��?��K�|�s���O��ß���w����5Ҿ�}�-�d�����99����k�<a����[ozyxtr��ٓ���?��ܣ��=�'�K�f˥��P��+>��!8*z�(�I2�H�!Z����K��!�-Z��ҁh�N�3ĩ}F��
l��zE£��%A6&���ks�x@Z1���󗟓�gh;�CQ�R8�R��}-ӷq%����Equぷ�d(��*��4g:R�Z*HpJ%�N\�c�l:�ƤI��Z����YIx�u*���1j�I�@*����Δy��nex	��!�^���n.��a���f��*6����;�jC+���_T�zmD4-�,
Dc��%�Ea��E��p9��bj�Kq[4�(U)��@�ٵ���CoHY����k�,��0�pk^a\�HA/V���o۟�o������?�RUb5R���Z'��i��o
z�an�:�3�J$��q��]�˰"�
�k�2��c-����CIp���[�1v��(0ԩ�0�9�B�ꏩ��y)n��\�O���S ��AV3Abq�����cѪj\z�J"���>�fmcǗm�=�;.��{��/	�˭O>Y?q�EA���.�c_�p��h�.}���WG��+�#o,]�0�ʹ)L�@�=���
���U�(C!s@Mʬ�\+W3""Y���*����_�c�� 7M�CR���@��rYX
�`�R8�VU�*�����~�!0��e�#LW�Y�A�V��쀕Q��&�h��*�!0���f���(4�X6CH��5��Kc��7d!k��Bp��$n�1�q
ѣA�al�@|8���`XF��Ng�e��^2��[�ԐUUaE�V��)gԓ�ߐ� !��\b��Qf^=pd��  �fX�1���I�-�,#�M��YF�aL��VL��y5���.����!08�����	�=+�p	mK���{p����k�
�hB*���@���nM��R�aOxx��-o�
������D��+&�)��V�O��`����,5;�J�#�!ym�MrMA���$�XWI��8�	��9�Vp^C�8��ƛ C@��K/ְ��b�j[µy��D�S�-m�s)�QS������P;��AB2 ��4[�<�!�hɊ��҄�iq�����&<$P�����E.v^F�gC*8ZS��sőΰ2v5K�&�x��i�*�DB�%���J�f/)/~���h8��%B�� y��O��RөC���45��z:��%�6!d�0p&cEr����BLêb ���C��!�Ȑǖ'\�)�,�Ԑr��p�����`�)S��;���z�tM��5j����)y�i�iRe��)�̺@�ȼ���+�!b���\���:���3�dW�.�����248�d��0����U��З1 &��K!Z4�B�U@Q�.#DaG�`�zC��(���QRS`pE��{�G��"�%˨*F)v�@8�|4�+�����ї������r�b���2�8�2����&�a=N�"�+,B^=�\x��S�bػ�V,re�Sos2Z��� Kz�6SW��BT��a�y�^kWD6����H�сּlt��!�W��bq�N��=+S�΢@�@�+Omy�ˮOJ
�q��Bhz���f-�\
qrSX"��|k?zI����ғ�3���!7')��Y�O^����E�w�6��&��onn�������͓3�<�qPHF�r�hݾf�qv�k�n�/��	�����Ɂ�K���nw.U�i��{��؏`.����͕{�W���Z��뚶]A�������������m��j���%?7��㛋�볫ǟ�ہG�ܫ�b���>�t���ʯ�ytpx�w~z���d�.���֪lw��8�"��jo��;�A�6���[\&��
���&^��1B6d�R��ב�6D�^m@v�?�k>�{���}�r}�������/�qm��jۣf]O󰠬U��\B@���,!5D��l� y!���xL`!�g���!$Zj���3��k7n�Y�\�iX�R��pQC�� ��f�f���m��.���kM��naZ�����>��t���X��UtF��>�X�:Y��
��/��H��v�׵��	D�n�+]������2Jg}p�ckIA�)a���_U\2�s���ˊM�+�!�!s���>Bs)�(^!5.F��p��&�d���Ͱ)c&�ڮ��E(�!e�շh�Rӗ���!X^!���ʠ�"��u��+_�����G?��'������/�;4�c�8:p.������*ҵ8�Ⱥ�AҮp��u�pd�=I�Q�LO�.x��E\�358͎���!��5M����9�]��Ě�~=+=���YS�X
M����;d�2/4|��s���Gٟ�ɟ�7�u��d2a�TE)	�os�3�g@,&��r��`
�N��dx�\����V�lOa� �7
PYR��珕u�+�O��}��������7O��z�������_��Ob��c.G�O_<y���}���Z7���x�����y�{���sG�����_�Go|�7o�ƛu�=�#�Ǿ7Wy�Ʃ��U�:M�n:l�ތ����1RP#W`��rq��&��"�aH�,z.C.�ҰJ
1�#hlMF^������g���)���'�l>�y�:�6}{�v�]CQ�ZC�w�}���B�@O�J�'��G�bPp]^a!v��I*L=@)4
8z6О/#�����1�hFe�߼�bqLJl:z-&���!���S�,(�1��#���d���K2�aF�N�q5C�A.y��c3�d�=�Ka��)Сi��q�$A�h�ҥ)p��L$/��F���~�M����8M���%P��0�7��𲨜�`�V�D^!&���]�m
@
�`2�j��F�9�MM��'��g)R`�"�$�3-q�x�4S�4.��l�,���7i�$�*�Y��G��C&2��(\Hkb�)��>�]�A��_,&p�Fj@:zQ�'K
\ڸx��a�Y��:�;�E	������i+��XI|��5���y�l�<���1��g��_�4�g�g����w�^?X?�m��z�-�V��Nϯ�:\����K�=�F�^�@�w�Uvy�[:=5
Nt�p�Z"��[4s) [/D�!�:����	�J:-k��KA/�a��R^�VI�EG�E���a,�tف�8�L/��3D����m�ˇ��5��h8�{ܱ'���\��م3jpF=����B֡s��K5��T��f�O�b+�8�p=>�N��E�8����<4C�!#�PC&B9BI �"�_..�^`Q	�֐+��2��T0��@:SO�Z��ϟz,5[���VR�&���q�X���!k�;lዱz4e�a�Kڱ3TIY���D+�A�ت�g�y5��7�(Dc���"v� lq�p������pM';Y���&j�Sp �<�c�İcM���,G���z`sa�А�`��&���D�|�Q� VF��J"�ܧ��c��p�!H|K~w(�\���g�'�/єͅ#$Y'n����T.$r���B
(03pB�X�l"�Ze��)[����K'I9W:\8��j� hzYJMח���� 
���U�	aϢ�`��j�g��,�t�I��f�k(�0��^�ۓ�*ח:2B���'\��*P�) �YCP� ��-hu��1nqwsiM \��-c�~�eB3�1f��F��0v{&=��;���dQ\!z�V..
�BH� 0���3�$L�)p遛ҝ&Po��0C_�rUU�8���Jf��͝����+� Z�q��!-,�9E'�>�6�p�&y�ɫ��\^3	�D��ʈ�Td��Bx�$��r.�V�2��U����Z��C&�F�0��p`%�ȧg �U*�!�l��e_�O�Ğ�@�Q�Z����\}���>U[y+���J����d��1��(W�����*$5CM=�C�!�'~������eWO�f��0/�D��R#ġ�%^�0E��p���B깐5/�},�p��ٺZE��'�2��p-&�^�����J�,A�>������l��IA:�,ȁV^j4 ����E8}C��\e�v_��O[z��ݟ:��������������؞�>�����9|>��<>�=M[\�<�����%�;{*�}y�օ��ۣ'g�G���Oqz%��E�u�u|���k�T�R����ٹ��~l�ӛ�S�tuw}E���މ��]�^���-ׯ_���'�)�2#w^ݶT�����?6�'?=I n��E���~��w��_=����g��W+Ѿ޻ڿ<:��K�N��ϡ�c�����=�Q��D��u�ԃ��[y�b�ِ� ���AԒ�l��\yp!�E!8����њ ��MA,����t֭S^m{X/6�O<�����;��%��ӏ}��b]�����.�t�}X�j�7��!��2��;�0�����Uȋly\�#���E�5��p4`�p��5��	I
y��c����� M8��ΰ�S@�t�4�E�:F�i���Qv�ŽL͇v<`1���o���g��z9F���t�(�D�������hn��S�;]��Hgw
�W�f<)��\.y��+fꑑr��,uk�ej5�'�@�a�R��C:4�0g���dh���C�5d �~մ�KC��MaԀΈ�,��7��E%�=��5����-,}�����J�a��;:ol�޽nZ~~�d���3G�{���[��~���������=��i�����,��UdN������_��C ��v4m !Z��E�G
fY�K�AS�>�l������ !�y��E��6���2VFI��z�	����m{������}�]K��4��]v'�!FS�R�R�[+!	4Q��$ӸT&W�VP��!;x�5����%Ff�R�E��:�u�ZO������CԞ�|����������������]~���^~��ᗟ�w�ȴݒ�9�:Z�A�D�./�������~�x�w�{<��{��|��ߐ��o.�~p{\U�]aVSo���L���Dfc�ߺIhj���qV!O��
�G�,*M���fk�d��FY%�����e���b��'^�z	ԋҤ�J����k����{����R�ꄫGs�tP<��1�V��J�n[z�����#;?)�N\�r)� �
hm?Y4���bq4x�P@�x.Q�`��U<�].j@�B�m  B���,#C��V@����h��a�� AЧN���@!hf�-#�i�p�lI'��(䕅��`ψ��#�T(�������sA5:�������Y�Ӭ�6�J�d4_"h�,ن�����ë�S�`F��f��"{ǡ,
������������)�����P�
./�--��2B|�{���$k��j��=����MJ)!�4��K>��ׄ��"aϫ�Զ��A�N�������dX�jV�h\�ͷ�S</�	�Q3)\�ȘZS�������������cWj��?���ַ��;��;~�����������������s>�^^^�{Qss���������^�=��ϋ{�'��<>�������	8Xo�=\/��x֔����U��V�::�+OT�	"������YL�1B�c
8�n���dW�m��g�T�9۟�D�鸳5
B0�� pF;�*p���VFy:��"W�a��8�+�5B�����r��o�8BR���    IDAT����fX{h�6H�^�@��N�����I?��\��v��*��R�h�yE���O�2⋝�C�D���
���h��~4������r�#��C�d��
X�[b8
c�GA�!���#���j�ʕ˼T«�4��c��;↢�3��^���p����N�V^�Wk��gR�T9P�VmC��p)cc�'�� ���8e/�KK�c��/ʐ�@D�ް�g���j�&���o������U=p}8�ꁆiVg����Na\->��V%��j@�lF�/��tx٤";�&R=bE	g8aZUQ=�2���G�N*��%�R�⪀�	L������9IŖHJ�
˥�*W�\2��C�אZC��\� ����04!&�2o��ğ)(p�hb��0GV �%jj�nI��$J�b��_��2�ț`=��Q�x^)��3ӡ	��G(���)#ڔ�Pm r����'�7Y�h���� �����?�e4,���(�j��b�-K�8����K3x-/|��2q����%K��*	�d<Mr�!�O�M�L"��1H���B�sq����d p�g�h\V�m�1�tP��i8 N��T��\-��"02Z-Y^C�8��]G�+��8�
�zC�U5���x�ld��0!p6��8SX������p�rAt��M�+)4M�&(�y�Q�a�3T���Br�T8$;M���.�'#�r�2Z�8�໵!�j��h��z�	$��8D2x�V=�z`��H�M"6B��+�=
솻�������P`Rp�p8�tqrALG��:H48�ٜ/\7��Z�k���IM����J��
���B������#�Z}C�d5�z^d��z�`��Է�	���~Hrmw��[��t�>�Z.�[]\�����܏��>�c����&�����<��Z� �7�Y���g�Ǉ�O}���T��ѭ;�~^�G1��.ή�n.O������^\_��塛��.�+l���}vu{����Ş��}�G^���y�5G�>���+�Z���ks��V�p��(�}M�8��_��=&������/~��_����U�>�"�B��8;zྪ���kR�bW�~�j�Y{��k:�^���@v�%b�������:/��g7�\zқ!��p�b�x�"�9�*|�ϒ�wr����h��������	�U)��c�K��W���ov�N��(K-�������l}�J�=����咔���oj#���&�+���`��Nj\�'#�`ↅc�I�
�2�eO�)��؝�Un`���E&eʮ������}��/l�Y�k}�,��������X0�HAĺ�W�#�x�(C�m���-�Z|o�1%�Q��`��-�~4Q=�JT��*��纮_����Jҫǋ���"���Dx�e�I7��*!h1�	��d���s��b30yK1,�,)�8�\�rE���4�p}F↓�1�ї���^�*��0U����*��t�x8�YR�_�yq0�]I~�Y��O?�����Q@��׿��ko�����o��r�7.��W��U��W�ԥS0�~h{�*p�'qQl ��e.�0q
��\q��6*�Ȣʛ�P�"���
i(��X"n�&%Q�j��'4kK�O�QtkS��%]�ƨ��X2*&�WD��ރ�H��5���͜C"��J����>��v�������ӣËǟ���۽����{G��N�%�����Z^\ܞ�{��������O|�K֛�|��տ=Y;և5}
��c�_羞���,�޵��=}��ѯ|�W��+�=������}����}򳏟��]��n���?n��P���[��K�s����l�^�C��!GO�,�������k���@�5�>�~��şh\��E��N�ENY�cGǐ�6�G��f�=`#z+��9�����6�-ΞN��p�2��@�[����������j��r:@f�
g�^5ת
�`�Iِ�6^ڇ�
p|�_
�|��=ڛ�֟���5Cg(�&�Vy��fX���pG���U�F�6P_
��V�d��D�����P$B����f�ӳ
�l���z:*�c�jqMJo�yє!�^TFv"F"�l�z��&��TG�tp
"Z�,)#0�*qN$be�Y�l�B�q��Uj�bKd�.�j��^:�Ο����I����}"�n��\e��#��%�Uv)�����랮���f˥���*[��gX«�	B�����C�RC��+	�a&C�w�p��FN-B���v�h�/�j�ET)�S	���k��FH��/��/�T����ʹ��r�����]���G����ͯ~�+���w?��g����s�_x���}����7�?��S΃{G���'����?��ǟ�=��~G��޾3�7��^�/�9�RЫ!O��x������������7�xI�0'x�ڎ�*,�ځ�V�Ԕ���n�א1ᘆͱ��N8v�@�������=��w�}���,!u����Kjr͚DH��Q��EI=���y��6�O
��V�~��cfcjU��^�g���i���7�;̆���d��([�r��V��$#���)d�%�!�����d�y�Ų����A�P,�25�5x}G?/$5^�-�NK-e�d�"+���)�Z���`Ë��c$��
̨N�TZ`��Z��V�����N�'��⎩^ͳO�v;���t�0�d�j���oѸ��_3��h���^m�����l.-��=�6/4ޔ�����*5N6�6�e���R�T<��].y!��VaY�'kXyc�2c��S,��)KZ}����E!0�y�_�\
p�0D46\��-##[H����mW�E鵒v\�M���p� h�&"*o`��68�
wh �,�3�?E!G(A�"q ��x# �LȚ��2z�l^��ָ4F���i��.�Pv�a=CK�k�J��h�PD +�F_�J���%D..�u�h������hҬ���hH�Y$B3��B�
q����Y���!E����)Tr�Av�ȈS�B�!D�(�-\���55��p��W'5�Ȑ��
�ȼ�ָ��@ e�ޒܝ!�p!E	aT/���`��j��W���\R���]����mS+<B������-
�Be��w�@�:�� 2}�^xL�H!'ǰ��aj�����P��KQ��*�X������W��AH�M��3�zӔ";q�B:�VI�ɞY��o�dI���ui�ͅ�~:p����7��I'���&h��c:�ʨ����N."<o��!�B�9$20�!��H�b#W�.�dW��-�.-������ӟX W�P�k@=pZke�c焐W�i���-�������ד�S�]��M�2��Q}vu��$���p��Y�H��i�2��ia �7�p�ĽAZa[w&a{>�h���rO�����ĭH�R��7�|�z�Kk~��5ֳ�	�w��D����O,���K���ח�ZHN9>�0�?���7g>�銉�O}d�����泋�=�=�{�}��7�o������5���'K}Y�՞_;9�Wٓ+��bNV���և1�����X���~�F��rp�(��K�mɽ�}75�mY[�f�r�ܵ����dGW�g�$�����Y}ѮOE�^<�<�W���{rx�c�>���r��Һ|�)������mQ���ӛ�)Ho��;�ېke�KU.��Ǖk���+�?��\b;��nh�	�z�+T�]�'bc�U$�)0�L��7aʺ~����
��g\b"PF�VC��W��UQ�jk7Y�V�a��P0Dck�=���M!�(dv��я���z��e�aYv��M^��Ƨ`:lm��NYo(E���_/�9�S���2���Gk���՜���[[��|����}�]�J�h�m�3v�����w�I|�Is1��dx� �&�͠N"-Zj��ʲt�G�bٮ:jeQ�������*��?�)Lj2DIb]ute��4����T�LĚ���2fׇ�bMT�\Zy �z����\�@|�Ʃv,���l�}Qh�rQ|c�]f���C&�]IE�q�˨$䩇B:M͒Z^��fs��l?�8
�����w�ه�|�*A�y���閹;Ӛ���o���Ӊh+���:�$�h�eQ@:�>?�N�[J�$�D��4)��ڦɞ�f�f^'��ɪ�|#���0ZCvǮ`45[.+��9�5��đ��֩�۵�]l^��xMRJ�ȥ�& Aņ��i��NDnC���>eHdߛ~|t��8�����~u�����;9�t�ސr�`������� ���M:�'�7G�>*sߡ���'4O�я?;�,���{����S��q�0<3�ݿٻ:9�{�?���_P��~�cT�]]~���G���$wq�w	AL���ؘ�	*��iW���)
G�j��v���4QZ��n�D��O���H��U����:�ᘌȆ�bf�y�)�){�����j�QS�@[ܼ<z!��G�3�m*6e�]"�gq�ő��]FW
�9=����1H�q���P^5��Zl���ZR-��zd�p�f��n�к1:j���Mx=�-T�y�)�����p5HC!����f#�%B
8�*�%K��6��6���u�4'6��65�k\�dS�t�B�%�Pd�Ԣ	�Ooٳ�R�6��Dn��BhC�y�QN�����Je�J#U঺V��������D����ƻ��q�*�3��3�ܤ�G�u�_�j����De[j��Q����*C�\-�^�K�d�d���syqx)�񒋽b��z�� U�5`"#��jmٌ�ovb�LI�В��6d��ؒ����S��@E���֊��������f�_��_����-����a�$�-�s~�]�׿~�w����_y��_����'�N�n���.n���|�����O�����>�̾/��s9)(�+��#� �%ة�!/o���7����7�^���<8>�*�6���E��;n����0����Wv.���� ��dm?v;y�{�ieL��:[7�!@�!��(���K���Ms�·T�����	� ���Lv�z�B�ʒm�p�WX�)����MGJ���.$W�͂]��S��';oY�D�-P���d�`6��R�!p1��φ�����MrA0�ٓW�j�`�-)�������hU¨��R��w���\٥�WX"�CYg$�\��Ϳp�S�p.�\�DVd�Q%\��S(��l��t��,b-�V�X�Z�ht\Ȇy�$�[8N��!q"�y�!h*)q^C��+�(8��Tg
�L��G��&X�Y�U�פ���lg4�_���)�c��K'��8l��髊r
��t�b�-��՟�c�ƫ� ��Kb�����F�iX�!��z`=�@=��z�M�!]!8��6jZ�}��gDS<�0AϛN�I����Уi�����n��1L�ѺÛ{�d�/PcW�����1"\Dd��	�G6w��siE1Zf46�
565�N�#5^�GMx�%U�[8���pU?C��&#��'58�.�bg�F��.K�8txg���2�.#P?|Q��G���3�h҅�W��(K�O_�M����@�3��p�\�g*�T�A���!s5#H:����DiՐZL=��!b�'��W����h��h!UhȻ�_l���)HQ_v.Fa��t�ˈ�BA��Zv�ADU�=0�"�דJY��P�t��L�)8��\1���v�T�pK���H��B���DH�3!S�<C
8B��Cx}���z-�XF�t؉�oʆ�WIh��<S�z�\�ւEJ㚌!�}-��@�[����R��oy�/e}
�
,9䔫�a48��t��6"q],���#K�]�^���zE0��#�E.i���x#p��qM�"�.�kv�@� Qp�����2(��6f�B�m�������U�S���v����r}��5R����������X�l�ۘ��e]�R���~��/��|K�pw{�%���^��"�Y���7Vl��4���O����ګ��n��Һ���,�[��J���\�ٓ]ו���'$ �'��@R��e�$U�:�VD�SE�c�w���z��pDu��VY%Yq�(�"	H����Ml]c1���Z��[k�ܼ��{.߁tUw{׳��3�֕_z��]�ӗ����G����k��Kn$^�_�_n�_%�3�S���qT�r}�(L���2?�9�s���ڥ��S�p=ؓ�ܣu�wS���a3��76]�_μ�k���'B76� �46��;�Y:�͕f����܎�Ok�ni歵�Z�t�;F�}�X�O>����Ho�S\������돱N�Ѯ	DnY�z�K�]�e���hq���&rW�$�qYֱ��;R�1�(���,�I.<�3]��b,JwYҟ	ו! }�!a�2j��ڙ]yy�/DKP�$y'9X��|�!�* �9�$���-�c��T��#,\-���f��E(�E� �'8G��=�;܆?o;���股+3��*qO��E]H���򬩚-�.�=C*��3F{ÖӶ�V_׽I�}C.Q*XF�T��`�����k]�T�;^��a��J^3�xYTE�U�R[�iT*;�v��l���B�blȔV3K0��O��ٳ �Hw�-0��	"�z��[̳l�,��,B}U�h h	ݔ�L���\��X̳���;W�ѵ��3�*0j�����Z �Q�1�`���oX(�����R+���:E��h;�� v�R;c �6� �x (Zv����J!��F:1\ZR #F# T��N�3*L�F5̙��R*�< 0��ǅN�9�7F�4U	����� �A-����4ˍD�@F0Jl�F�y�\K�������y*��YO*p���񢩨��[7v7|�-��������7�n_޾q��Φ��y��O�6�,息����[�:{��o�>�y�
;wn�{�{����3ך�6��񱾽��½��x�ջ/��y���x����ܸ�����������y�����W㖆��!�6��a]���^���e.ႺF�
�Ă�"�6���IS�̛������(�h��
�˲�40�2��C ���BEB{`n���G;���~pkY�t�N��:B�W_�������ރ��������.JoE�5(UUF���ql��/	
��E9��*��b���<��ŌG���@`kQٌ4E�9�B�ʋ���j�HH.`:/{�d��#x��U)�Q�X��(d֖���1h�Z�!�kU�����%Ѩ{�����+��ɡ�/]��� (�������k�!��r�'����.5E,���l`����  )#��آ�ٽ�c��,v�������lW��6������� �Ư�\�N�*������_6����
T<]kߪ-�gIx	�nީLXv�\edT�S�a#�P�.��R���KF�*�9�����ð`��b�D��u��\�k��|�v�(shqg%�FE̹���	 ὂ����w(O|��>w��I�7���\lm��� ����x���޸�<��q�/�����~�����?�￿��G_l~qr~|��~i��O�n�_._�t/��pƷ5���޸�魔׻3+�d�>���U��Y�H�4(cl�yMB�`I@X���u���*Q�fL˥Eh:]7'
�X!-�@]�S�,m;��w@�,
3��R�
�M L���˥˨�Rk6d�C��R���:SJ��f��XL���â+oTu��N{x�D�ЅW��RI�eDR[^!�����u����h9d&Ul�����\EE���i���g�,���`F�]"���dd,$]`F]Rl�U�"!�,���BgD2i��B<��$X��!\�D�#d��.Ke��Լ��Yf��v�n��9�U�WT��P�\�e���k��%
-%|��H Q��%��dd�C&H�<,�dI!�a&��@�Z����H<����`�g����S"��0,��%-���Z^,/��N�Qt�����A�t1�Ÿ�^3/���p�ȵ�+���Y�`$� I�fRW8o�*���B�*XKP��g����M    IDAT�R /a�%ye�0!�0 h&Y
ׂe��D��g�\��I2�.|�":cŨ>p�u�0y�u�	;<c��{�3z����4E<�� e�:<Q5���kg ��6���K��,�J������i��\�ȵ��74]J� ~ :���!C���â5x�p�Ʃ�O$c�H�1#)�,\�kW���0�N�1O@�0fI�&����V�Nx�\ c��W {�	�'H��aJ�e~$����@�Q�_;(�Md��*#�#B���
��E�Xm�V�#�FWx��!�I�Tŷ��J]a�N���Њ���,3	�"W-/�Q�Fq"jhtQ�,H�R�,tHBg���F�e�0R� y��t]�.F`^��@F:*���%���t!#���`ጣ�eW��ϨK�x�L~v��ж�,D�ԓ���Rvv2K*c5�`�`�<-�*�t+*` ���ga�?@�
�.�6r-Yh�?��+$q�E��0PlZ�.A#6]�IK�EX�%~m�u�Vx���7�6�VI�V���+�.p�t�酱��<] ] ���Q�\ظ�\[��/�n�N��)��x���	]]��W��y����}\��y~����K�k�v+s��|���l9��r�)�0}Z׭A>l]���}�'(u�t��Ez�����]��lz����g^C`|q�WE�Ql^�"k ��>��>O��~x�dn�}uyz�W�;iMY|�����0�o}c�UY�\�E:�gR|=ӱj���]8�}�sͷ`vn��g����O�-�~~r���#�٩_�9��̻�rzr|�W�����l�$�?��O��l���7�.׸���[o��G?��o�ڦ[Y�.<޻w�>�Iw�����#\S��{N\.��L�5���evb��<�z.�-R��|�ᇮ����o�A��I
f��ţeW0E�_��v�E �Q�n�Y`&-}")U�s�cӲ�()��Γ���^�ce�7/�e`��&k­T�.� �!���z��������կ�^����E|�w�v�f�#�K��]'DkQ��������]������J͕4+L�*]���;a���0�T��� U~��}�޵.��wG��1;�EH�.��b�5�\v�����'���E71pe(���.�~1_�+:N��	@FằM����v��}��	�2�3����\��sM/̌�j�Nڙ���ײ'����o�;T�< #����b7��������#7Q���1!�R�<v�)�Fn���v��d�	�\V�v�ޖ`����?��m�+��Yv��*o�J������YBy�1�`�KQXӨ�� cF)�b\�6K
��h*ڨ�s�&;���[ݡ5�kU��㪋�0��y�F��J�΢��"�������h�øj*�3-��+{�Y�>ͳ��/�o�y�t�����f��ڿ�?���O�������ȡw�x}}g����������o��x|��������m�������x��מ�p�Q�[�;7����޸��{ӫ�j}�GU	�ura˼�«�����W�_�q�y��7�9�1�EX� �ጃ���ϯ��o�9!L.]�XugT��) �yY�a��hn��(dz)�(V3ڢ؟)X,����*�.����rS���N� �jS�=�΋D�(��
C����(���KqB*��VN�]B��m�7	���W������R	�0:�3v�a�7�X�رQ�r�k;&K��#�
F��	PI��2�F^-ad�����+��dDB�N�I���ҭ��*o�LͲ4��q���5j<�&M�tv5��.U]m)"��g�D��}���eIY�)�.�5ʮ[�C�b�T�.�Vи��j-�p{�vBV�t'S��!IQ�]�7Qd�������*����Aa�r���o��W�y�Ev%	�`Q  ��E�	 1��Ki�Sҵ	�S��_�K���*���m�Au�Ç�,�pň��u3ɼ\�Z¨��"W�r������Y�2l���rMr!-�U��v���j�[V�
��{Q4Յ�b�K������>�y�'T���̆s��������oǛ.�0����5̫[�n���+�_����ov>����m������㣵��6�O�6����oll>:����jpd\�H�C�'g�+��%'K}v� ������W��!O�YҲ�ʖ�+�t��|m閉ѴkG��V����&�!;�4u�&�t��`�%<e��ɂVK�e�J% ϴ ��Ŏ0Ω,A�H�ǯ;�14d��LL�ռ\���..-��-6m]Q�6��36�V` ]�k2Y��L��?N���X.��
�����. ��X
{Ƙ3�o�1��Wu<`��*El���S�00Dx ^2�b�K�J�2(!,$�,��K�k���c�,q��FH���	ɞ��>g C���g�&��Ψ��+�����`#�����vJ<Z�;S��T�:WcaY��k��	�6KTH�.���=�W^�FI��Y	��V9#�NJ���bf�&�ff�9��R1Bt��"ᢔb����
���p��3b�<,b+��#Q!�f���8���J�f����p	�NX���d�v�K\,�,�c/6/���0�R�Q��0�`,vE^'"��(�l��g���<[^��P:�L�2xrF3���%� �
U��6khM�g�)��a���&GK��D��eY
�s�`�S��!�%���4�0QI���(�����3#��
3�8���Z���ޟu��q5#��j�b�!�S%ف��T�s�*1��6R�10F~�6�1j��rE�n3��N���k�0i!�7j����X捁��U{������7�B��zFQy'��@R唘�,��
��>3R��`8'�R'��B��N 3�(e��(�j��b$`����;S�zX�L>0��bW��t`^�\�e�C��b�ņ��¹"cY�G%j�L#��+#]T�L�2Rx��ld�e���DE�GD��"���!cCkU�XKa��,*N�@
�,��+o�b���M�e��B�*X1�ޡ�Ѻ��^����X(�Q�}���0�Bj�Y�ԍ�ޜ��V���\1�+�b�5]-|�#�u��b&�D�B� �
��p����%��9����#K�(~��ݽq�e��#h/=�ugy���v����{�g�g.aܸyp�����#�>�W5}���mx�8�y?<��j[���w,�|Gҗ/��I��W�mʦ^��.��v�����[�.9.�Y���vO���⡱Jr����2ʚ����K����sOC����]��WO�M��sܬ��m-ϛ�L��7}|G��\�M�'�O��ӳ�S�����Ұ�c�|G�˨y��q���CKfQ�Vю������%���YN)F��OK�B���R��?�x�:]�p�B�;a=������k�F� u��m0�ݎ�V�~�X�/���7"��B����Ga&��%6��Ei@`�1΍ >@���rL�ӳ�����:��RX�XK�����ZI�g����<���B%��\����j0Kt^FQ�g̘E1��ͼ�uY���_���V��-� _{�{���f��ߢ�l <H�JK���(	3o��-��tG�n���UZc�4:esU�=,�}�����QH-��s��]1��l9�� �F
v��Hu2���
&2r�aS���ҋQ]�4�.��d�(20�׈�R�k�^T���)�J��t�\�ڌ��(]"�v��8W��f�����jGk�<��N���V%�,��՚:]��di#;n�h;�}:�DZ� �f���Zj�5uv��fP	*b� ��.����?���t#��b�Q,D���@"#Be�QS�ad'y�2�
Ha��$��-����di�k��N�0�;�������g��D{T�:��PJ�"�աK�����e/\ˮ_�Zi�:>��+�({[��h�h>���Zvq��������+�r�fg���������?o����4��7�x�¶�.=#ݓ������M����<?98�u�;����x��p<T���|jɵ��s�}x|��ȍ�.ϟx~�/�|�+����O1����R�hF֧/ �Cl �8�<����);���huYx:�x�G�f����Yf
v:#��\�V!�W)xY�Ғ� Ym������/��f����Ε06��������W�������ٹծ0.skS�6R��,^�6O���a����+��(��JeԕT��;S �AB�:���� �@������1�v�`�X*�v�X^��\E(������)��.�x���%$�Jf��E�^-$#K���ԆP�(fa ���UI!&�Ԧ�2�JQ��g,�,��Rȫ^�5�ZHv���B�S�s9��T�N(�Nᵅ�t�K`?h#0��J1����.�O3��_��M�����,`W�px�B����9��v�?z�g�\>oo���p�(�׷?�rC���`�4�ꑎ��6��N�n�i�e7�	F2-�2��,��E�!���$E,e�c�m���&�C�!=ag�?3U�,mn�]���ZS�Ŕ��k�]�	k�Q-�o��?�����?��K��y��Kw^�΋k�w���щ��m������]�0��!���v֞�}����}��~t�=usryqtuz������?���'��~����]�֑�n���/��p�No|��b�������8���x�򌚑Ni�f��T��B�غtbδ!���fՌ�؍%E�Ң8d��@`����T�ɢ�zRI��Z�(V;@�
��hS⡋҆���rtL�\	�	�X�@�^�*Y��g\-&<	�6�1�J���i�
��+��ЦLT ��!���QY�H�j�3#]��X�(
�� hu�
,��غ\��E���m�1��LI�
���tq��;�(��!u)�֦�*<B�`�t-ay��pT�S�^+oQ�b�H���2��j@U#a��[���*���y�K��r���:ԭ�`8Il,�b����Z:#0�F�+0���e�9�B����k�U���'����Ho��k	X#*�n���8�)���<�2�EUß��͞B�MgOd�59���4FQ��֢�g���B'�0�t�B8�X0ƙN�ɫ�	]/;%�;�W<�J`\b�-������C�(�Hp.Ac�X����	�.X�Z�y�)o.<�%�3�-#N$᫜7$E�'���^.���T��mF'tvx��g�2°��(�=X���nQ`�>L���n �0�m���J�y�2�ې�y��1��T�`sȼ\y��!�6%@z�$o3�������W�a�SaD2i�����Ω�"�(�V�
4��w,��œ���jQF�\Yt�4��:NmS"Qj����W�Ws	/0Z� *�s�V�(`m�t^H��f, ��;pI'y��@�t	ڔ����Nx�d�0���Y
�A+��X�*o"/���$�<E�;	c ���(�`>����$~�D`G(����C��d�Bѥ�	���Q��6�֋�X����W�I��8g��?���{]��&`��bD��N�UIjf�F��\���:�`1�"It1�S�����۠(ƨ$23�s?G�;13��=B�sn]\��R��2u��H!�2��K�% "��iHD2N��M/@��������C�<�U���]x���w.��~�S8FƵ��֧�ꍋ�rCҟ���w1�7�N=��j�����$}pw���H�B?.�^��r�W�^ҩ/���tv���[����n��<q��w>�7������˻e_89;��^��>�C?�L;����>�]s	W��[��W�k;2z*�)�g|���C���I#pӐP���+B���;}rza$t0�1e�}9i�0�����gq��E� v���J�kPތK���QC*ƕO��tGӽ�u[b`�;"uqZtJ'����k1;����i�P&f��p��j��P�tv���CH��K�K!� y�ٕQ8���	&/����Q��׍
I�Y@�U�𓍋%<e�G7�Z�КC����� Y&߽qs�u<To����n�*�"��n�|�ogZh�� ��yz���:��f�wB��!p�M�]��kJ3�i ��ԆÈ��$iv��Wv�m�н{�\lwӈ��3@�S1b���n�����J�ń4�*��5]�ov�����M�:��)b��
ϞNI`�^=ڦ��]/�3"�����n<��0D�
��!���u*�Q�-�� e7�����g�6������d��j��J2<Z����?�cݍ�Rlr�.`f؍.8��VܽU��jޚC`[�Ȃ���ҥ�dd)�Bb�5.�zTB�d)�y��!��B�����>���\���v��c1o[]jo�*�0䐘�h��n�sI�Ґ+E,RSR�f���M�����x�Q����if����l��f/�;c�]����ɦ��W�z���}���-O�Ύ9���o��zB�����/�}�G���ɱ�����g�~;��	���휌g���j?��vy�ʲ����R��m�u�3F��������mQ�S��.��i~P�Zs���n�-dv
��R7��3�����0�Ċ�0�2{�/u�y䤥�����I2.��,��I
@���ӅpU�XݼtR��p�γ�D��q9�H<��؄�r��_��镁��q��:�KD���lͼ颳S�dwx����)�E
:��tf��1/#Bm) ��[%��N ӵB*'=�<���˒a��b޴�P�4:�*�zHIv��bˢ3K��E��3���3FW�@�9^.-#WST"<uqr1Va%U*�j����照��\�n���� Y�� ��/�n<l�������\��u�"�0x0آ�0Z�#Ƌ
�eMg���A[:C0o���2zu�B����#��J$Jk[�*{����k�cȨ�d�i�D%�Y?|F�i�4{��d*uCʸ
�3.���[���@�YO�F�F�^�il�F+�6���EX��c��E�^vBA�b��e�ߞ9::�����o�����?����{��ş���?��;�f{~�K�����~qy����/�>nm�^�G���xkx�����w�vxg��f�v<W��������������ٟ���~�������W�\}���'_?>���-���d> ���
�U��6aK��Kr5�Z^F�dD�6���V��l��;&e9�i;�1pNqD�F�_0�"��.���D��	���H�;ۆ�_L5@���d!���I�H9��K�.b�ɾ0]W���. �XW�@V��)��+�rV2C`��LNx�2'�.���\�������sE5,� �L��ӆd�q� -�v��a)Ex��-�@Ө��i* ��-��ExY�!y;Ƴ�Z���C��ަe�%�X�t�R�e-��՜��E�����% �E��[M:ek�s�TFHmCF%�(z�2VL!t�$�l%���a�C�	SHF�����g {�:9�!�(�X�\�c��ehPUBf�!����I$q
�����!�+I!�H��S�-u�f�\�H.
	m{2�	�AS��8�����a�$QR�j�B�
��92
g����JL'E5��`Z�DT :X��3���{F�U�,vcQ�dԎ"�?�θJ;�!dY�t�=x�X&��Q��	�)�u	N�d�kYj)��ɥ>���
�Xb�5���
���Q$r^B'����I� ZF�
��"���O�"�9"5�(��B(��huF��ڴ�⧻�@0̌�ZPch���D�Kt� #�Ra $�6�nl#�24`F�x�q&����eѥS��oٵ�$�5 &�b��K�����r�qB��a��Y��UWK�o�@v]�8g �����/c�Q�D+�@7��s������`F�G�2�H�6�A6{1�7�xb�A��gg��Xތȁ���uS�W �.-�8i'�*?L Fz��/��e�%�WT���]!�,��@`^-�&�H�rѫ9�*U -Z��r�	��0�z-��N#;���dD.�\�������?x�hg�Va3�,��T���8v�*    IDAT�n
p�!�a��y)�N�y�R��p�U�d�JI �#�<�� �e�7.��b!�����ׇ�bv�"�j�Rw�+x�e����u�ðh�c�p)�]<7�ƻ�M_����랾�Z�]r��$�ָ�y�����+���,؋��ǖ��n}��U�9~l|��Uْ^麷�ҨoU���N��"�������O隥e?�0�=s-�a���Ʈ�ͼ:?����Q���"�S����䱸���¬������T/\j�����x-�8�:�ܕ�ʺ����|c�]Uo�7v|+e�Oc��i��\�x�1p~z�~�
���g=�w̞�1Q6�Hb��M�R��#m��LX�̿%V�0ES�Z�(`�[t^���2����E�)���Bt��3�	Q�$Q1�3ݗr�D �H���2�uy)��$@�\`3W��;-#��d,V���)�H�N��fd�N駱�,
�1KQtB���5'��h)1�Ĭj�Z#��` ����{��O��O���7���ڿ���p��v)ֽ�O?�Ե�n�����Å$QL�߽.̮G���(���q�:0��Q�|eM�� �) �@��J隶@�f�N.-����0o����`�X]7�x�C3(!�s��=����f��Bm5�2c��R��ty������ץ4:v$�]�b���E�p&�$p���,�nY�\�R@.��?�M%�6a73-�Y�:�L&�@,&_�TH: �#ۨE����s9BF��(�����.����BxeHJA�J)�Ր !b�I�p-���8g��ʛ-ccYh�� �(.�����(�bT�t�Z�
�З5�ϥu��A0��q'� �����Fe,ymnv���� D���gT<��0
!t-B����W�Y/���A����o�l���+�=����������^����������[��������?]������l�o�B��x����o|m�]����|�SA>�sӋ����xl��8;�i%�˔q�e5���f������x����s�XO�j�����]�^��k��2^��#�)2���U1-,d �C��N-$��&�d��m������BT �0ژ)s��ꂕQ���KD�����+d���Og��j�"�1�q	��X`*L�azPg/�Z+�+�)ҁ�"�.�;�b`$m<��Z/���V^$�L�Bt�M#�z��ryu��U|�U�=/�@^��!E�u��e��׊5(�P  �!=6mF�\��'!�pB��:Y�PX
.��Om�b��$d����?*��,eL�
�#�3L$�i��4K�4.���s��L!addAE�%]�-<�6���y�.��w�ZW�6c��O��j>�KD�h�Bm^�ʏ% Q�~������V�ڏJR�"�ې����IYfl��d����6FYP�hS��сIF-@�Q[w�Dv�U;].��Z֢.�2��U�슟��h��W� ]�8Nv:LQy���Y,}
KT��@1����q�g���-�V��?����������1��]��\[?㍗���>������^�Ϋ�wn>�摇������ß�x�wX�;��㇏<5�`�������ue�oO>y�3����������?�:�����W_��_����寿��������G^����xC���<�Ӵf��	�9Ʀ3i*��g�i��	��7�4@0��Z�6���^-#�YkC2�n�ͤn)����.#B0�J )��u)����.��I/v�X��0�jTlr�-E�f�i��Zx�̧qi�0�0��T۠��!�抅��������t-�����KX��˞+�Z<eԭ��/Qe�[�����%s �Z<���B'*a��,dc����:<#p^.¢�D�+�^7|:0{�2����D@��*���I�R��~*���愅^�&gbpFRmڲ�r	Ħ똢�����uq�]����	ɫ-\�~�D�����ԅI�Q��sѹt	Wy�sa��0Z�	��vx���[v:��#Ġ&9�m]���<���-KF0����.�,����bx��63Z0$�x)F_8�@F��'� �eF8;�n��|ೀM�³����*Y��W�`��˨���SDI��.0z� ,�g�Yxs����R0sUU䫹 D�6����ri�HT,F���$$EF-�LLg��C��'Ί�!d�3$X]m��E�e��еa��P�59�b)K�8�#�nN�+/ B23�j��NL�x�s�(�)��`t�%hL~�ȫ .�j��c@&�(F]z�q�"sE��ސ�0��ai�pu6`F)) .樦��]��k- R�[t���b>��-��@-&��Ȩ`
W�劙�.@�t�W!<�VW�B�!�'2�a�C�.����`����Sbk)���vz4 ��6iY
ײ#�j�Y)�BGۄ����Rv]ƺ�Q��`�хa�*v�t&�V513��`>~:�=oQ��䬫
��Z���;�b���bq>�lZ���!�Ȝ0V $g!��WV�tlUE'�ؐ�jY��M������Z��MH���,NE"Q���'�\6� �RH��7�|��w��\�+�.%�V�.*-<E�YB
/5c��p:�
�j��=6.�:��֞��s��8Q�H"gG���Q[%�U�eL�M��pbVF]vK12�����q�Ӄ�}�ҧj-�G�m�m���Z�D\n�������g���鋚�e.�V�թw���z=�6�O)����7<	Ͻ�+�ݫ�q	vo�3\O�ON=���r|_ӷ<!�{:�DY�yp޷'OB��D>E������7^< �_tk��8G�OO��Ϙ3���1	[�~/�N?��y{�W~���G�=��H��R<p�����}�M�A���ʻp�v�k���)oݹu����L}�S���b�X��S�Z�^d��;*�F,:�M�і�Q��a������=�8Vp9'�p�F>Z���^`q�B��%SX<0Our�+dRlQU�.�
|ŀ��-c��K��xv'�R�	�ش�Ҧ��,��0d��,�
8Z
p-�d�e�.����/�kw._�B�����_��E$0��� O�5�>,��J�|��|@q�QӎD��:�[�R���ul�fA�J���R%H�}4���^.��b���X\�Ab����,$�W1�t��ݝew�r"u��2]/���V1��*�m���^�uה��N���N���KtBgצ��ar�L�U�� �����O*FIa(\SB�������PHQ,�X�r[�H�B.ׇ��g����(�0��@��B�)5�h;�;�Ă�L�=�6�p�y��P�� ��S0A�2NWOxv̎���W�0����+���,���Ar���\+/�B
;��$z�w ���fV��x���O�����Ć��o��,?��*���*�����9�����(�@��,�(<��,`���I�8%#`T����E�� S���ڌ�@K�u���4;?;�8�~�!�O�������u��ro}c�������#�z|�~9��iFQn]�mz}?���ed��ǣ����#Kk���SJ7�/|m�u��˫S��|{���/}co�ܜ>�kԾM�&��i*���НF0�b���n��-h~D�rQ��
���(���0?,�$	 $WH�t ���4�hՃ3Lc�|����R�����'�(nmڋ��(�������v�tR�� �NΤ>����eA./N]{Ɂ���#= ���,������g�Hk�����;���+��T�.�]6�H����s�x�ޔ
�@(�"��a�Q*�` Q!Y(`Z%����f�F!0Eaӭ~^H-��Ȩ!�´석7#�RM�,ɒpd,< ɂG�(�8)�C�DW^%ѵȅ��*i����p���7f�),:5{��o֑��ț��U����s��'\Nw��p����z�T	f�����m0�mf�v�(̔��z�/+(�T�i�H�e���k��t��N`�������:B5N3dg',Z�fX�,���H
�T�Bt�k��żp\o�X� �lD�ȵFo�(�������R� ��+�zI���'�/�+/���}����?���~��S��k/�>�Bty�IGG���Y���aԭ��q��'���O6׶��uk��;�<w���շ��)���'W7o��^��޽��7v^{�}��q���畷�����_����_�|�us��}uz��ѱ��f�m��A�6��!(X�m�F�mz�i��N7^ô{������<C��t'�^m�a���������Ħ��L��E+�%κZHvm`��,�r-�^���Q�6̬$%��R��.j$�2(0f�zx�1�Y<�)�J!�,fT[T+\s��l�R���Z��P ��)t��L/�R�t��\��U@�THq�S0�\m!Q�@j�D2QXJ$��.v�Y�kz�ǟ2]�$���AHt�K�UƼx����d��B�ҵ����bZ2�mK1C
��t�3�Q卧a΁̐9|0Qf\��v�j���M//%�X ���ڱ\3���h���jY�h��q
��ތ�-/d��t�� �e��^�=)$�l�I�V��^,ZR�`�P��!'�(R�DR.� �2j	f��	Em�TW���x� 1���R$-@̺I��0uZT�k�2c�F�P1e��:R�ȳ�@��e�����W�u	����$���N��Ж�Fwb�3"4!�Y�3��)��؛�-L-@�Q[��Q��2
��X�%Ҳ ��[YvQ`\����U�E`0����*u��dg�R"l�Q��'O�iUұYU���<��Y��l]K=�YxN0-�4%Eff�Iځ�$�5hj��Wl �X)b�7
]F]
Q�,tF�Bo���mD����t�x(3�!���۞NT��r�U�R-Z� ٧�B*���6���q
ӥ��.D��I)` HHv<���QèK`�� �mJ���:�g�S�zI阵��N!������^vQ�,��C��P,׌]��������6]�>�%eW3����,Q����g0��R=�`�jnCFO�іH^�N���,�t�2;��1��EK�m��Ĺ��+f` )��Ӊ��k�g�#�qV\�%n|>���e)���~ ��Mw�\m1����ȵdr�,Zz��"�y���n:����tx������n����e� w���%fmF,����t�����T�k��zyv���}z66�{�n����{�'���������^��^]��;n3�����k�㍰o]ڣ�9���'s�:T�k����\-��ڸ<ܾZ߾|y��%YO���+���־}r�9;nE*��ָ��N7!77��5x�.q#Ҙ�u�=�k|C��,��|�q�4��{�VE���3���0%O����:s7����������g��5���|�p��!�=�֣��ӔLԆ�V^��NN�dV���^ώE�!CI�bi�7-XQZ2���
áku]&C^�]�p���jY� pba���� Iz���YvWH�s�K�?�:���TRz Q$ =���7L�� �aXp2�e����kug%y�4�9u��!#;�.Q���E ;=�R�צ�����^�y��O����w]�{{�{���'����=�P�5�nV�S�c)�\��Y_Y��*�+����(54Esea\�A(�t�[�D8ZBYj���ͅw��H\"��u��X�)���SwM�e��>���O?5:���f.i}q�?�!N<�F�"\-�5b�bו]K���� {-#o ^�0��� 0΅l�ARJ$���Mc����0�q���`�$<c�.%LZ]E�j]�4�,�tH�i-X�mv0H ����
�ՒH ���@];!�쨪A�����_�t5+@j�Z���!���Z��u���Z�f	�E��ERҋb�Pv-�ʵ���O�l�ǱIwT�]���ۿ�[Ǟ�mJ�M'8�(���X��(���D]����j0*c�`,Fwz�	������_z���C��}�˥��{��o�\yi]�ܺ8;z�Trvq����������˿z�ߙ���[�k�W��wn:o�_�g��w<�}k���k>/u�x����uO��9�P/~���9^|>��9��g�[�>>�֭��O����u{�������c_E�{9W��1�1���s���x��Zx^bf�I�u�.�qF�4c���b�W p�����#�C�`�F�!/	��͘�e!���$B���������1��:��C��t�D9KW�c؜h}��y���Fu������Ӻ��m\�J�9E�ݩ�"�!8ZV�C�.�V�Ĭ�*��ʐ�E�5�`Y5�qj�RF�T ��Y�@Q0�Ҡ�b���cw�㩒K�E�$�iۍ�ص,�Z3�H��� s9x��T:���ha�!\��B	֜��%1햆+�0	��hEh�sF]è�W�鍼(��2�c�Y`f��	��D���s��N����L�n ci8�5���W_������,>�k�������e���jh`��)@��� �Z� �B2f� P��L��#�<�>�@�b��ՅT'�%#�;1,�$� ���*x�=f��,�O*F`��Z�"e�)���(6�0�`�-$v��,�Ӌ��>�6�Bkw��>��$O�9�y7��-���^kg���������_�b燏���W��>�է�ӗ�����?}�?�_�?wc�ᗿ��������|�qx�|w�׶o���k�Ͽ��;�~�_~�շ���k����G�<6��>��OQsb����j��Y�O��p&��9Ӗs��t�d�ψ8�)�T����WPQt�f-���wVt@�L%`�8��"Wr$���D�^l��Hg��¢[�-�(I���̫Ɓ[��d���Q8�]���AW,��+��Yv!�`��V%�xF��-��� u)$�6
�LD'���%tL��l�f"�& B[�j��'C]`0œ��2݌q�ײ/IF3�Ų�,���J���`Yx<��_13�X�Q�,qvDT笇��B�B�vc�Zz[�a$�B'\Rҧ���!uy�)~R3����-��c K�L
�%/{��Նd���aӭZ��UKl�d�"٫�W 㬁;���-��6 ���rea$1�E˕�=�@�
g�Ԃ�a���%�z2�^a�4C�<��Na�C(�Y�+iFMe�Gh[���7�1 ���R�����J�%�$̮%����f(W�,��#��]��Ѕ@(�r�zqA��ç�ad�zlaXtks���M�����HV�x��!BR2��H��
 ����`H7�6��0��L��O=Ό媅ga�L��1h	<c��H��P�W�������y۱hY�ҒjK)5�_��(<�yY�O/�nB���
��]`��R<�:y��'s]!0� ]v�2,�I]v]0�H�d��I�z�{:� v<S���C��bg�fln ��e$[R�Y���d�Ǝg�{���7�����r��!����R��!��g�µj�&��tѭ�J �� ���O0c#�,�V3҉��i�)P::AHD��������tT�(ye��6��@5�O�o0L�X�� x��k��*C��<��+KvJ��MN e3
��$�S�FC�ZQ^�{^"��;QfI\HT��&��X���LRUKĨ<��m�#��5��uqյ�2�^
F�͆X��ŗ+ /<@T�j�w��N�ؤ��%,�x7!7�"�o=.�����j5�n��;��O������ڞ+��V��ˋ~�r������nm�^om\�I����������̓��=�-u��ۛ�;�{��;�;����>V~u���������'R��]޺�v�p����-�Z��b�|��j���\�Yöv�`o{o�̷P.<��]3�u�ᖦ/��om�k���@�r���6���Xߦ�����t��h=�V:�d�_x�����~���	y~)���F}�a�控^�>��=Z�K?��n�^n\x���/u�ߠ���ڜw�b��UkE���#�����sY�i�N�>F�x���p T�Q�@T@���'��Z^�Ӂ���X^���+�t    IDAT��;!Kx:��Tt��Y;-	&��C�>�c(���.*{�Y�v���_ϱ�f =#$�̼R�f�\mB>��c��<��W�]Ht\���;n���'?y��u��te�'ץ�����f�qJx!]�q-�W"
Kש\ZqD�x%��R��NVvN�l�\UkDE�";���H��Bh��Z�n*�W�N�t�e����%����Bt򱋈���$�A�Z�c6�Y�z\��g�y'2�\A���(��jKI�Wݖ`�y���6�=E� �@,��!I��ץ<C�6`��eWzM�E7o��t k��F��֢�W	*�vk��W�VƺM�p��:��Jc_���ui&��F*�й���l9���_��,E���Xl6�03]Q43Dx��Nq,t3�1c�@��A�E5������OɄ��!�*�(H�nv4��25��^�,tH	�¢>���n|�gcs�K�����;�/���/Ύ�<��:�xI�� �qo�����ݽ[��Wk7�~���|�od�z8������웙=��9;9r�5y�Ɲ;��;��~��w��|��ï���ͩ/��k���x�>=[�P?�y'�`q�x�ܿ�w������������i����^=|����>�䱶�r�"��� �F�KI�F�o��y ��*@&;����DQq�%���3EQZ�+\�����T���)��DQq�W��^8��a�;�\��ilSA�㪃�3��9��
&�F8B�MTe`�`^H{�"�\6y�^T�I���,`8��"��4��;��a�� HZ ,*!t���%���u�$�W+P��0g�t��%��[Iɋ��%���*Q]��N�("i�H]lD�H�^����4�pm&1�	4X^$`������//�,�
m �h+F ��E��E i�����R��-��)V�g?��µ���(G���gS�ɒ����y們ڟ>>]���K���`*���������{������;L���΢*m��HR��L cvF�8[v���k)愾�Xw@Y�p��T�fɈ��j�[ʪ0>�5�6tv]��Kb�M�����,t-�"Z���3��y�ŗ̿�����q���'�x|��ˋ����5�����'�>�|r���]��~���?}��ᭃ{�}��w�6_�s���w�Ξ<�����Ƀo/OϷ��o�v��������G�^�<��b{o煗_z���>��_}���G��{>v��ֵ��Y�ZE�"�Fa ƛ0r���B��}���xR�믿n��s�I��%;���Gv�κ�����K'X����{�#y�5KMa$0Zx���겳�F;픢���2x��p���8��u6!tY[X���Z#�IrZb0����������6? �j)��
*�v�P�y�jv��T���`��X:���,d^8]$\�U@�Y�$!c�����qZb㥤�D���Z$e�Q��"��(����5-�rQ���~����E�FXx�@�"{���ri��*��^vH!�E)��!���.$��Qx]�0�[`]zR���$m?.��m,�U��+|��0�9���g�3�"56vQ�6�x�0S
���I���N!Ml-K5��H!� ��8;���)VI�YU���6plbyY ��I�X`ҵ��SvF¨�39-a�b���	#��z�S?K���X�(0.]�Et1̃L��0z��G�"����2]1�|KF- �Z��(i�Sm����Q"�Uz$1L*x5G`&
0� ST��.�1"���v�TU#�>�L���d/��*���es��a(Z�t^��Rl �s+�(^H�i>X���a��tu�buy)Dy��+��Ր�\����b�-����R�9��Ղ��5 d�:�� -�l���2jU�^yMQ�x2R�D�c�Td�i,P�*�.o�E/$�����	El-W^-��&M�V������k2Rrş%��ΐgua��H��tkY�u�&������D�Yr��5�!; d��v�H� ޙ=d)���Ws����RyY&'#���Kf�<� Vg	F� /A��KW��` Y*�t�fIPT�t
|Jm.<�8�j(L�,`�,�z�xk�UN.RRm�ͲY0h+�ⅉ��`�Xt��bO����CrME���\��{�/��(F!�UC.�k��s��AHRb��]�����Gk�E�������v��Iȣ�|��j���f���xۻd�ϵq���I�r��m�\/��A��K�{;����{�;�~psm{gsogw�wn�>��ۼp���s���7�o��9��ui�w(�o��~���ƞ��n����ئ�N�e_�\_?���]���_����ɓ3O������H?��6�f�=/�����v��{`&l����_5�����I������c�wַ^|���u�s�Y��s���^\�v�Y�K��8�;?9���/�u��d|s����O�G�^�/r���Z��Ŧ�R�K�*���Km����x��S@�.*:kG�-s[Z4�v/���Q`]4������*������I"K�I��D%,2N;��1�.J��>�%|��'�Q=�T9B�� 캫!�S��:
�M�W+U�,��5k��*E���*�7���?��kw.�������=�Ǒ��{�@� WI7Z@ \��.�V��f3��Z�t��ሢkC�,�Z3S+���Ʃ%��^�bz!�t�K�	P-<-}��Dn8�V����!��q *D��ʨ�4ɨ��Z]z�\�u�KD�6]��S��q����ez)�d*t�g��B�n�R�#~EV�0S�5]Z�x�����M��;��͖�eL�rP�I�=N"��]��mH[��gkTFc��
A�E�BF�7� �Z.^m"'�	f�qp����̐U�8Y2V?N[b�J�#���>�d���iqټ� ٨�����VFk��$��(	QvG�8?ʊ��b8�0S@����V�aH`$t^-=#L�^�ؔ�"��sc|����/}���8���@�@>/0>j�?���!���^x���z�?ٺ�gˎ����~��$[�mYmK��nL4~�y��O^�<BMn@��ql!�%ۺU���}��'�wWz�i+k�o��o�̙��\k���g��g��=�h拓�az����e�-ܽ�������ʽÃ��S��x�:���?[]����=�Z�����S�8;]���Сs��W�}����_9:z�������ƽ��~�ߓ�y��ER�l
���LͬM�9�U�ke��a�f�̵B�;
G_��F��eԳ�g^H᪊�04��G��!�W��e�jq"$�x�Z|=W[B�Z�c���я~��^�NF�����t<�=��q���G�ي���]���=�zR���^�y^��+[�-��z�����Hh���ۛ����x�'�2��g�+W��)���*U;M�h��l�-Z����sr�1���5T��V�R�nRE���BT���� G@��a!� �!M=j[g�k�g�h{`���e�Ԟ�;�[�B�&����Q�pG�rA�����3}L�8@���-.)��9�f�A���V�����~�ƒ�)�p��H����o�Mͻ��sIg�vm"�\z��yB��e�(P:4:@)�J�h�Je õ�2�G`�F!�z!���1����WX��	��RB�^Il-ev"Փ����/�R��ڜ�æj_��
3���{���K?$ ��/��~�z��G��,����۫�٩�i|l��z�uvzur�z���Ow������W���7���������'�>������>���q��Ӧ�i��~�o����{����;���v�.�p����{��n�?�>x����;/=�=q�ۭ5�KO�MM�-�P�����-&PkI3l$��,v��F�:����IJ �7�hh��x�%k�,T��V^P��v|�����Y!��c��gJup��/�v;S,�,@H�4I��2��l��E5Y �p�0p4C.d-oC��4lRz8����lY�S�Gc�g�S��uA [%��!��%bWcF��g�����s�)P+c^"��V��_z8&Dx|�, ��P՜&`
f��uM�x�`&)�a��jp��n'.DF�b�i�U^��`�(�UB����[wѤ�	�g �b��	S,;$EEf뵒2�M����0kkjֶDR �'h(K��V�2G8�z
��>���� �#�+o��}jV'��T� �h�Տ�8���9Ad��L[C�xHd}:��Bf"^`ErE��D͈T�i�g؜8�줐!�'��g( 4��f��00='��9cfg�Oaf,Đ�5���(�a��	�!5� �9�G`���k�V!zρ�B�)�!i���B��Iy�UÜ�z,���Aa�X=�q\�)'��T�x�'�X��7LӬK*�B�W��*fR!S�!�&�NI��\Br�(��KT�%讃#��HG/$>�+�hS\l|�B"OAC�X}���e��4�o�r���	������t@-&���!q l�,
�ig���$��=U!�l�h��Y��5Ga�:���Кl+� Q��Sl���Ő1P�Eu�#�DN����*oEΨr�ǁ�F����Ԑ�h��@�Dm�%bh�3j�t���bWCQ�:�JͰS��Fռ�
o��XC�+����+->�����S����� \e������>�.H�05F"U˛K��@!2�ʞ�M�9�v���p��������/�.�4J��3P�$[�(G����B
����Ԓj.�)Z(�)���l��p�!)[_a��C�!
�~�)�EɋHD�}��TƏ_&��xgg�:y{y軖�pެ6}�Qsg�]o�7/6\U��K�;��R�8����O4n{{s������O����A�8��'�*�%R�RWW~��:l�]\�����<{r��0�:&���ɥ���q���ĺx:0�M�o�8��i�%��-��\�;.��Q�e���v6���5��tLw|!�j�����E�I ����]��P:f&�gD?Jv�
S�����{<:L�f���k�i��8����˝_�'�;�ռ��+�I	^��g#���I����5�G`�%��5Q�D���65����z,8���;��;E��I Wp�{�=�5���cnRhz�8�svB���a���8�z|R�l��7d��Y���o'G�u�h�B��Y2DcT�,<�����������#gK~����?���t������������eq.E�^����Z���$	ʥw!�,Q{CR.%9C(#ܹ������� l���IFH�A��\jh8��jJ:���+�BT���L�n1S'�|[Îң�������Ξ9�Kܵ^�6�	W�t�ϙw}
�fAAH�j��v��"n���P�'Rlj�PT���U8t_<l�1��yŖ%C,N���w��-���p�8�%���E�J���3��t�ü<~�6ֶ����]���˿t��U��l"���)����a8�B���.�X=�%���-�!+Q���B�-H�H@-BGČ�^H��)\8�D�w���!���,���ۄzO�}GH�&�A'�Y�3�,!��Q2ř���+e��Wk�8�Aed�(}ޘ�dpƬ�����x om^~��oV�nM�w��*����@�˞No�n�������m-O7}�r廛W�~����o\�ߤ���NùM��ى���\���7����Γݛ�_x}�`�`�K�������3��q��׿�_[��~��3U�,�ݸ���'nw��~Y������+[����|��5KgM���1��ߑc��y5��ǪrY%�q�i�1����b;�zC=DH�j;���f���p6~���.��!b�S3d�K��Q\�U��+k{ԮS*�6�4����y��7]����c⤈�M
?�$��@�b�\=B�)�a�K��m�g��j�8�Yo��!0���I��lL�LR��h��M3d�&�D� .�
/;B!@LC"h��!N+��-�_\å���r���WI��)ę�5�$��A#�К@z�@(;Ò
4�E�I�d=O9�� ��Z4!-u�،�&a� ����i�4��S�gTLht�55{�5�o|�^��;r�L���y�w�^�\���ou�r!�۫�w4)t\�cp)��!he��h�*�5�^��I�h���n8b^l�8e+E�8�f��@�!$rvY�so̼b�X�^�>0qC�z l-o/�v};D�z��A��~�M�*�����˫g�g{��}`��/�7���;�=}���Rw��?�l���Y�{���I������	�]����~��4���?;ٸ��ʝ	.�P���>���7?���~�����I��`�e?�|tr�q����8�}���Ӎ�3�9�� ~D�,m��m4��l\ZGV�\g�&���&�3��C7�5q:pkX��l�-j���9�P�@�VOx.qk^%zL��(d��\���B&��c>�՜�s:e�B֧V`�e)��me������kI��~�D�������J=�ymřwV���bj���LA�S�'@���kG?��6�+Ψ�4�Jj���ew첁\y'A8�
@����6%š<+�h��h�r���#���!��j*gğ&�*d�VLYRӇ���f�Fy]6>52f䲘Q�>NHC}̞���K�� �ɶ��%\#d�Y�
���\h��ek��Eeg�i&R�!0D`P3��G@�*o.��:
z�TY���Fn^s
pL��lm�8�JL0�z^6>o�jhX o�j@� 8s�r�Q�&n�U��*R�\�rycN�Y�,5�@MµY�!|1���� j��,ʲ����M����Rx��sɂo��ql3�Z��睕�jj@^Xwcr��+@^_v���2�! ��N0�7�p"W'А�� $0|]�(�|�G���-����	�˫���>k|�b�`�q����A�P/�Q1e����,i�UihՖ��pf4Af��Sgf��p3�8� )�����K�!�ā�2*��B2���ĥaj\��1��+)_k8r�=���2���'��&�R��=	hl/�ӱ�)���ZI�d�g4�95HYB�L�Ֆ+}5	g7�V�
V Z��A���]�X�����55�/$��\�B �8x6<�el
3���V5. İ�!���%ꙍ+�,riw�5�f��k���BL3B�\��ѯr�+O:�����cRnF�Z��f��(�h(\�i�4�X:���`v��g)ijsj�bė�,đ�E�0�8�sAN��s����"�gN��'�6/� ���YZ�D��
���!PI4�O��jyS�����Bci��ć�ٖKX�ؕ�P�x�1����"�Z�Y�>y~q}����\�-߈D� u����R����G���{�c��`nK|�ow���n_���������3�)�Nookw�?v�z|�s{��U.��o}�x�h�������f�	�������;�6��ťogn�������-�t��.�7��3I?湡�qmq4�0���57�b�.u�Z_��K2��^��M�PvG^7|���8�wt�����hʴ��}��:��rZ����Ү��a���ʷ[�7���e�>D�,���z�eO�D�`��9L�:V�XMv�!�;��y��Ds2ӟ��;���|����;�%�v�SI������}φ�p���~!d5y��*^1etd�YT��@Lӄ�,�Z%����>���J��b�%%��s��B"���w3���׫��5�W�#���'?�ɿ���;a����گ��U�sQN�Y�>,���eh=�s��lGm�m���YsJe���\D�r��1��J���gS���{"�5�W��Z�J�cfd�T:�)8�n��V�[Ό�7�*
q�	�>�}_'B-�]�?��O�v��iY5����t�E�(3�4�I�@@��\���k\I���&q.��3r��*8ðj'8�d�"�3*@"��(�	���J��S��cmݬ�ǻ�uz���UM|    IDAT�]ל�\���fW�~��������@�2͔�L�����b)����l�4^"��v��(DvX �e�����pdY4dB�qzn�2ԬL�a�'%���T��cj���Q��RX1�C�2"�b�v<n}������Hl����	q�����ԁ��Ͱ�L���T��vu�=����2�C�Zs��맭�=6}0����2������������������������7�v�5n��q��K��`����jʾ�����<w�t���W�?��::���Ã��׏���֦������k��w^~�k�8~�wq����s��������������;���ܯ.z����1Wb�V܂����h3e7}� �s���P8�Q�Ş��JB�\�/J?3���#�ώ����T^j넊i�!s��Ϋ��ve�m/Q�
�\Z<lO�{ګ��*�b��A2d�w1�يo���˟�[�4�p�(����w��̩�V��zH/}��,�81[�l.�7�D�����+!q�2�
�(�&�~��ϥ�"��c��D���0�4�'�5x��R ��Y�jR��(�6���.� ��)�M���aG���U�E������C�8���6*[�)�$UIir�m(�-m�^�����n2/���
L\���݆�T鋕p���c��-����]7�v��Y��j �B�]㷇�K���R��,z�6&�<��5�����<<{��=4M
�
�3c�1�h�:�F�J��h�F�,�W:ygF^8��e!�@8���V���G��!� ����8�8��?{6^ǻ��}w��\]���؜��ݹ?�����i��������qW���#?��1��������O������ޜo�^���$W�W�Rs��'9��/�}�s���ճ����ŧ�7w��e���䓓�㣗�=|��������?���~yq����mR��r���q+��6q�j���ĹL����L�Y.!� �,�_��_<�0EA�Z҆�.xcZH�lTjv�(/Y�Z��e�5A�+/WI�RjVCI�����&�_1��'��p�e��8kL�R�Fh��[���].Qb� ��OV���S�j�_��"�F*AF��a��&�:*&İ��I�T5�6��+�!���zd�9�l� 4MQ�X2ҧ�+p6L�P��P0rS�%�k�LSK_Hy���㤙8\1��jb�s%l��k�M��@��k��\ZY��!YY�L�^�&6Z��	zĕBs>�q���)�5Q5	�``%���(u��3��hي��p$�H� ;|H.�rM������0l%�+�"��"#����gkU%�ؖ��`Ax��d@f�a6�,���MNG����1f�^
��O�g��Ƒ�PC���b��*�JJʕ#x"p|CmH,�� +�>�#e
!D3Պy�5/:q��O���:�K������4�
Ξ�Σ�Uv
8���	�T6�b���&ȨB"l�R+���G���<&�S^(#]�lM�w�bZ1�����V�T�ِ+�rEV�U��!RÇ�O�߃:�j�΂���֚���U���!pVȮ���2�C�(ܰ&�(����zf���ZBGǶt&-D�k����L����r������M-OBR�*���o�yUU�)H����!���o�tL�P��Z��٣ieY��Bd�����gHT�ć�"�����g���j@��m�V�\��R���������*0�55#��Ѱ��D�Я�D�4��MM8�&��G��-D�s5" GK�b���6�N�U�gOm��2�8d�X���HU$oƌ-���DO'A}ê�6A��d }d���N9�P�д��,��qѲ͚�2zffj�56_/��
 �t���򍜖�&���8��Ԅh)�%�
4�DȆ-�P���@:p �b�be�y{}5��LdL�p�7.n.�\$�/a�����w���d���e��q�ѷ"�w���������qjxsc�ӫ�����uɛ?�r0n�{�L��t����I�g[۾��뾸꾖{w��_
���ݺ���7�U���������3+�������X:Ga���z��8�o{\�Tɵk�"��罈+|ss��ې�hg�/���o������͔�W�ϟ>�Y���!>�t[�ͺ�{���k��vo��O��c�ӕ���T�=�t�f?��!\b�{NY ��쥿���j:}E�'?�����ߋE�ɰ̈́����'�7~�7���ȹ~gMw�� ���./�?j\_��`e����FG��e���o�K��?��h�����1�����eȨ�U�!��aj@�!8�8��CYK
�a���/�$��%. �B���|�;��[�ey]v~	�j
AQ��%ʧƭ�uZjQ\��Pv��xC.Q�=�	�Wg;JH��0�hD�Z�N�P��z!�d������y+h�)�>�P�?�Е$W��u.jvJF�T.�=����۫��'�͹��iȮUa�44G�'Ͱ��F<\��d�C����/d=v�3�Mm�&5̞:V�t��&b��T�=���7V���ow�ű�I�#��aKj�=�}w����\�<��i�(�t��mf�qᎈ�i@͡4T��4pw�Z8�:Ei�66�c^l�A
��.P�C /e��pj-B�1w��VF�9Z��?�ƅ��^�Yc�$�G��[Q:��t7�݉a	�!��Ahh��T�L*0,���l��扼4?O=>o�|��/l�f�u��MƂ����U��M{s~����s���nWg7�~S���<>y�t����?W��fu}v~�v�^#�6/��#칓�������]�q���#����j�������4~x���G����'g'�7W'{��W�����\���n�iM_�|zv|��d5nG��C�cW��iM,��vyk�om��%���/{����a}�lA} ��z�D�;^ʘC��p�U$�����G�G`k45s�es��bh�d6�jHʅ�O���Ft���c��u� W==��C�\1v��GO�]kb[�>��\�^=n��T���`4�zV�u��`G���\,��ȋ�<-����BS.�Jت�#���`�F_��uX��g<���h\��<�u[=*G�eN�AY��BYf/���G&�B.�9��R.!��@����V@1z���P*>��}j��W��V^�(�jJMV8��S��n���m��@��^�ME��ϕ>�{�+=�JW^s.����b�����S-We��(�"�c]/ħo<L���z�
cW^���T�l�,GkXT���!B�5�h���5�b���I�Z�b!�w�W�p��(�i�!�/(w)��!Ô5v�heq�]6�%�S&���Ⱦ<?sd^#�3Ǐj��*�Ww���;�3=��[�\m<y|v���;��|����L���r9�	}qӫ�ם����7���׿�~cI��o�o����jk�������?8x�����·�v{�dk�����?}����GWgon}�՛[���Х���CN;d�.� aˮ� [�6�av�*��9��Y��B�X�t��\��r�8B��&
1�pL��^a�|6��y�Ӭ<�L4mH^!�y�F��^3*iQl(��HY��g!޽�2�Y�r�ח����LY
���#�J����d�yJM��ՌlH���,o�B�%���������x1��q"�e�[�!����2��y���S�EʎY�p�33AN������s���ہ�p^�dx��*�㒍9	K���S��P2D�GӪA"j���®K�]x5QD?C��\p��ټIM6/��3�p�p"Ryl qx�,M.Sk^�\�C<��Ѫ�]ѐ�d�qt��R��@=�l�4`:�*d�5��P�l�/A���g&B�m�QO ;׬0/�\)O^�b��5�z�@j�l���n�>�8�'+�ެ�b��������Y�"!�&5ժA,;qC"\x��,�����0�;+)>W C�^��2H��-q���L����k1�B���_<�B����-�M/��s�DX���dTR=��Y}4�eDf`2�
A�J�jMDA�uIm�:^�a �2d�d3��B`TҬ*N���5C��6�AnF���a�R_v�V�RC��M�0<M}�r��d(iV���	/�P�G��sUv`Q�r�NB��U_�P�&P?�L�7>\�@���������� �T8\
!�t<�p���es!����"��~�uM�z�0�h\��2���,��23�Μ0��E +\���F�����K�!�����y��ϖe�lj�� ����9�j�G+�������j�Y�tҟ�i��,��P�jz F0��	6SC����7d.���zr"���]�^R=�^�v�D�U^�gБ4M^���ߗ5m~�{P:�ҕw*Ԁz��Bh~�;���C�n��a�@*>�Zd/���2ʘm������r͞p�j%�y�*��y��<l_:��=�?��:t��w}���oLz�9k��{�^v���w?|���'u�]��e�q��c��K��7g��wv��븿�g:Y7�Ժ�3�.?�{vy�w�b2n��;%N�9�,����`W����{,��"w�sk��j��/P�[м���!�[7�&4[��-*y�1߸��a�u����d�}��k��/�������ǻ�U�R��>\�l��0�)��;�)R�qs,�rN`�g>�>�o� ��r6��vl �#x�z��$��L���G����:���и�a�w����4�y���lqI����(p����mQ
���9)�m�q�Ґ�e�ٚ���0��q&��B4R*�̮ADe.ּ
����2�1d�>&C+;N6W!E�4.6;�d6�`e؊gX��@�]����Gk�Ĳ�h���j���U��K�U�G\�R�'�-�������E%����l���5��Q���ф�Z4�,ͱ�y�3NK�I�3����C�t0y5C
8=��7�W��e���z�L�?��?h:?O�/��/�z�-+��3��E��ѓ��Ԧ�lj����\����'�2�(�Pc#LB�ρ�f�W?��4��+Z逼������~F��W������}d��}��y�n0Z@[�
��l�YpWF��o���r�[gJ!�dRzK
��8v�eS�^mh��\�R�� "75���Ѭ5�B�MG�)끓Y�@����%"0\��q�P�+G~������<<=l��#ъ��ҟ�ٟ���FzO��5�$4�������5�f�S}<M��Q�2~��7�-�O�x��:�w����w����Ǜ�$r/���s����[�z�8�tem�����'כ��{7/��[&xָp�֙����#ߜ�w�t����w./�?{���O��/V��>{|{�_ٴBO}c\%;7'�Ч�����{�U�p����/���^���?:?����ű*&+��{8�V ��׫�,�D��>���	!�#�0q�b��@����^#ײ�x����p�P��C�;�t�b#��(R�8�����ұ�z`�5����p�Hd��A���ċ��ׇ�fR��ǰ�i�R���7�|���\%"��Æ�lEW�m-�-j�k���lE�t���0[���a4}Z�R�1��^��	�!m�I*��>Y�!C�rQf�q�[�j+Q��\�����8h��A�h�D��MĔegk��z�@��b��%e3/��)p+i�!e.LK�&���#�ဧ�g�T�1[1���\4�f�V�H�pd�՛����뎚g?ȿ��Fh�Ѥ���Ϟ?�g�oz�#}����Wd�{ꭒ�d�4j���U���`��)ÅDn� M
�	�cA�SӸ;
l��ɖ%��z!��g�>M}H"��7�ȴl�bs�gC֦x!�*	�o��:q5{�����V*e��põ���Ww\����[�{~����'�W~a���Ư>�Mh7p[���vḟ/?0�����o��ʃ�[�|��o}�ۯ����������g��?��U?rt��k���e��������'�������_��З�~�����O����/��}��ڱ�P�o�+�j�jk��=(�@Km:�\�vr��ۺa2,��)г�!#����6dc�0�xN�ƈ�U�����S��[Uň-�<p{^=��2֐��5}�ѱ�^�.V"���.�WH�1�g��RTy��R	B�BR8qC3��B �M �RV@R�@��2Byc�~fO���>�P@ ��V^�9�V�zj�K���d�z���ɎdKW�@
�b�9M���C���b�/��7�Μ�QX�S��XjC�+ٙ]`|�*,���蓝!��RD����m�T.=���ǚ��{LA����Rdӡ Dc@�$�Ԁ��X ��ҁ�"�X�M3ע7�"�2�������aFHg�t�,B�EEƯ��6�����q�5��
�Eq���A��2���<���!�GC��٤Zj�uN��I�k��l^�DiH�+o%���);��g�T+iv�j벅������M�7�lx�
�ڲ�E1p�3Q�-N`����`s�6eV�!#�D�&N��
$�9����qU���E��P��|	ָ4 5������0��N��ԑK�a �eؼR��0�%J*�#�P���q*x"b#G�m����)���Y�
�	I��tӋP�8�
IP����8k��ZILv��y���Ǝ��8�Yd��-P�z4�˥7�b�h���4
�<D��©=�w��C��y/Q�駦/���/�c��0R�4C
��4e�C�k\!����:"15^��,o8p��uy�͈`�
K|�h\� ��N�@�ԙ�!�L6N!Eńh��!E5#��l.z̙=MYֽb�5�h��	��-�z^��ˈ鸗%�bqZ��ΫU@�(����N'|)g,c�6Ĥ��ay������)�.;e�8����a%�� ��p^+���7M�l�i��-(�Xjن���&��j��t4:��\�W��3u,>>�ī�P����?6�t2/�׌"��qwr��T[��q���Ζ���&
�,��5Rz�|2�풤ߕt��%@��2��`.&�҇���g��C�;�'>x�|��:���zy���#�~��9���Q�G��>2���k�l��*�����n�s�_�t��W>�]t�q�c��K�{)���zU������m�|���kwwV��Z]_��芪�򷺣�,�8��Ⲩ?ީ9D���l��{�o��s}�$�x��|���$6�{\���W��G�������lm����3?�v��q��{���������2��w2�-7�.ƍ|ǒ����G��\�V��J����;��s�l;Й
�M��m�|=��k����G=Rp������&��OC�� N%�N.u����xi���N~*R1��Ȥ���H,M"y�pC
zMa���Z����t(k\y3�j�ɋI�W/v�g�1����-���l�e�-��@��W�W�9�b������AM�%�%N�F�t��VBv4�1�egЉ���z3���3 ZU!�qU���P����F�i�*�谚�����њ�������P�
y�_"�c����������t�:�-g�q�q��n��j��##Y���q�48���^��`Ø��TLù8F�֣�ʨ��qf�R��KZm���q��ֲ�*�����X"GM�J�nay;g�0E�-WC\6��?�sQ�q�c���ٜv�A6&�=�k��6SI2���[o�
�aҺJM��瓾6f(���7L�3 t�JeK͕����`�HJ:a�6W�elX�r��g��S@��������|MO_:�r���"e���.��R��a21���݆��KaH����X�(xsV�˙5t?$m[m�����/������^ �#?^[�o�o�ݸ�����B�G.Nn]o{���s{�:�ã]� �� �㜳�s^X����C�W�Z{�CE���}yq}�N���    IDAT�F�����n�^��|pp|{���~G>���.v�<�Y��@�����?8:�}���_�ٿ���֑'t7	�&w�����,�T3\��Pd�u�ge,K�����G��B���M��̋@��m��0�)ܰ��2
dhe��j��r͹L���"sY!�b3�=���o����bk��������،o~�8.X"�K����˧�z]wg ��d{|*	�v�{��xټ*��
$k����B:O�h��!А����BY��t��
I��������A��b9!ry����f��bv���@��[48�!�\R�R�W2}C�c��s\���XQ�V�D	����B�bX���T6�MIz���\�26�X���ZY���;�\^N<1��LP�Z�C�(�Ѽƻ�i�z'��fS������^�4�ߛ�0�5!H6�2���) p�&�hMM1
�����^ٌ��q41KRF
��ע�ɞ���q����7;���h��,�uwi^<�����i+��- |�@�~_�j5���3�^)v������ͣ�r�_��^]8��^O�������^y��og������������ۯ~��W���K����'����~���?���΃�_{��{�?8�8�|�O>ػ��˯\�_����͇^�.>[]��7�n6>Z�l�l<?��:?��;>P�I�ۊ�Y�P3�����[H�΀d����zb����V@�X���څ�h����wQ�T�D�>7�G��S��.4"z�Z�+{��6�r z☢�qb�Ic��H"0���S_IM9N.!3�1��Њ
�k�qE���(5�1G�/�^�zH�d��e�Bf:��)~Ê�x�D�0���n�����C��%.����ϣ�١��VcC��jy����b2Z���_,B��@�MG�F����Th���+�����0E5�R&�.;Zᔛ�&�KkȨf�h���\U�xƇQ(���2,{�Db��aL�J�� E��T̒��� {�4%��c�&2��n��g�:!�A!e=$}`%��O����VR!xyM��򒊟2�!e��P+d�/�N��!E6}`�Y
.����G��e�/���@���⤳n�I��_x� M'e^:m��`i�����Ҕ����(
m:!@��^aC�,�@'Cjj���2b"T9�� D-N�U�6���-;���P^�Dz��R2��2p��Q�z?�B4l��-62YFvK!0eC�J�j�Y�(��K�;\/�ݰDq�RӇ���i[^��솢��{��Wj�P�,;�!J"�,	�x��S�Z�Z�@��1���bȂVHC=D�fD��!:�ڲS�7^+�>pz�W�
V!C��2�&MZ���F��G%���iȂ\Czi�dD����Df1���Ȕ�r�h�s�`~�`C8�pMl�)XpFG�a����S��jN���G+�`�^�a�q�b��^N�@Q�+8d���͹�Z��4_6�&���lFLv4uE!C4��[Wy[�l����s	_�L�2
$��Wg���Kl8[��~������T`D���I�X�VjŨ���"�={L^��D4�����ֈ����L��)��H=���&3 �)"^/��,�f�N}�!&�|�%U�3Z�����
7�8� ����t��5:鸈'��UUʞCd`�J�v;�����ۼz
t�V�\������q+�=�^��-~���Z�S�����.Y\����ŭ����ŭ_�t�p���!���v�۷�[�>��G�m���v��6��+~scϗ*�i�&I���{;�����hC�����ۘ����W6�������.w�]~���]WBw��n��H7�˦c������G�Q���c�w@w�㳓�xO���?I�ҭ7��v.�ǽnǪ[H��Q����8׻��+?K3��=��>���9vT�=5G��rTGsb(D�G�K�h� 	4�s\����m��X�^R@�]�?ù�7�?�)S��qyeqjԃE�v����P/��1�p��\m�.��K8�le��J
��Py�aˋ�^fj@��FR\� ���$�Z"z��z��qu����݁�B9������g��%ur���#3rYHCs,fOǁ�B�:y2.KZ/�&���(��j0����୕i2�|^��Υ�^��(
��(e�@B��ѫJ,���\�B�[Y��%"b�9S���=�=r���2e:d�,f�V@�N����p���-
��E�gH,�@+6�avxe�-Wʌ�21Iя��#�,�$�>)�e�.�!�b�_'�8��a_!�t�p+�	��Po}�^�X�!f���ͳa�R��,8�N/;��8>A�Qs�C�!���"h�,)Po���iF�ag hl�r	oa '�L�D:L@`sI�=)<&c&�Q�e�����W��W���ѥ"_�V����S���j�(����>����s&
b�� ��Õ����M�y~;z�..o�����ך���d#�����|:��h�v������8���u�M.��^~ɱ�w���y>���l���׷��c���t7��˓��{�P���ON?~���׏�?~��O>~��ۯ�������|����v���֨���x�[>(�ˣ^�w�����/>�������/{����^�m���ܲ�:Ns��q`��D�2�`}'+�A�q�p���@ez@}��
N*#Y��Yw�0c�B��P����"b���.C�zpjZv4C�GF'^����,7Up��mS�6�WO�ɞ+}u�C<,q<z�t�+	��%��lK����vo$.�N��V5�NO�*� ��6ك�-\T`�����_/�Dp�T�!/XwO߭9�,t*�a�(p
�p����).P��O-����!!I�AA���G�W�o'4�D����p4+�nI˨/��D��Aa#��
�!���petP��[^^���ٳheH�J�݅fq\����K��pJ�j&B��L��[��ZK�Y(7[mbjp�l=�X��k�6���C�y����VRGa��qU甥�
C�NIk�e��+#����4�.�2�yE�)X�.[U�!{���(;�^`������}sx��>j�#�~a�������}w�Ҳ��ع�E��ˡ�[�_����W��x�׿������W�N>;���7�I������~����n/�vn�}6�����{G��W�����������n~���q�����//W[��o|�˧�ǧOw�<v������o5���{��e��h���[.�{L���Z+[��e�������n�3��e��h�Q/��wg��J�ŐH�9���в3RP�av=~3���đ��H�K=�R.�%�9�!� ��&Pc���(7��gFH�@����1���l`��%AG��g \IϞ� ��c�g`Y�"�LWTjz^)��
�A�{�@Ц`��֧P`��ͨ�R1t�pfkY�4��e�ݒT:)�!�/v"h9is��D�I9� 9@ƿ(J[�P��e��(<<5/M�3
"�!��WO�\1��0r^�d�&5	�jC�-f��N�2S�62p�6'[�d���%琪�)�	4d�0Kg��3s�KDj/|fO6����d��6���d���\�a��Z��U�Ӥf=8�M�W�5ްY����Q�j�u���և~�y�5v�:�Z^��c��0J'�h3�"1!56P�>�j���0g��!�,��=�VI��@4M�bq�s���Z�h�-�z�t1!�u�J��Ԑݐ��t	gcj��٘|�8�B�^y�\씋E�����Ф��P�>��3��p��YAy�/e[�b���I�(��t�H�����Y P8>D�F��y�W�� ��=�ǜ^R�Y����??:��:��5l�d�+�JD1���#ϼK���4g1�f%��\���啨"�B?|�����z!z%1��򖑫�K�����8�8-{
���"���7�NP3�%�&A��5���dh�fg��ak�hlx!p�7J�`�U@v����s��T"�S���ٽ�U��b �-�s}s�А���)�QVv �ӗb2��s��x��j�"@-�b�'��%�Yf�;�� �f*������q%��2�54-e [�bB©E�Cx������4�?� %M����li��)ȥ���_F�DU�@��'?P\�x��aR�Ef�iQ	r�?�*@��	0,�޳Mk��_��)� DdL�'����ړ���R�����o7�	���"oܬ|���nk崫/[nl^�II�o7\w���ɽq��\W�nhw��{%.v��QG||�Ӆǣ�m_���<���!�ۖ��1W{;.���mn�
�{ɺ�����]��霭��^���=�q��bu�g^��6�6����P_�t�ZW}�tsg��j\kuD�J��ۮ����Mw���VV�8���ظ�^��祫��n6;��y���|����K?'������八�7���w����`�����c�3;�1�p��D|�$����1���m��|����ks�@:�PG�u�����;��ow���ǡ �~+��<�s�v2Öp��퍣�ќ�O^mv#��ޟ�[�1N5�L�4q���x�3�+а�p�-�^I8ڔB��0W=\�u��`+3FE�j�&�K^=����?��ꢦ�w��{���;����	Dky=? {)����JZ^K-h�=��4�,8R���tPD5}.Y�b͈���B�c����G5�8lm�0��'7)ȪS����u/���sF�����~�u5'3�:��(�?��?	|k��iR�E^�t�4�S���ҳ#3�������hh�Z���J���+$;oQ���
aL����75Q�������^L�ɝa�b��X?��дU�?Pa�=x���!-5qW"��p�1m'�φ8�N�IG��G�wo�������7Q�pC=q�5�W ~ǎwN��3��pC�R0�8ͅx�3/��0A.��Z���	R0#�D���ۿ����������i���Rl��������W�Z��Q����4>���%�,)��!_�`^�p��Y�^P��[W�ƫ�p��e�q���xv�=v��W~*��j�}��ڝ }&h�
������K�}��_�����7�+�=�8�-v�=:}��K���Ϟ<���=�wt������^�͸�w|z=�,�CZ��i>羀���ƵO2,ϸ^�ն�wx�U�]?�t�tur�&.�n�P�W=i,w����[
=�"X_�2�x�	��=جD��̵�e3���F!�����u%�x��&�6ʮq1�䪤8ea��Cj��9�q��^��p�f|ކS P��/^����֡����c1OZ϶v`RՌ�lh��e4ĔH`	u6.�!�HF��5��q�*_����o
B���B<�=1 Rs��d�HFj)T-�z��fjӅ93�$n������~D�Z6�V���Zyv(���\.ΐ���*K+	�Q\E1�d34��D��U
X^=�&�2�EAZ@x�˨�ɝNO��2�,���V�i����b� ����>�ov^K�{tR��덂�D�̈;��)���=�����W��U�h�R��e�2�-�u��t�k�B��tDe�2���MH��S�O����`4�u�0g�"р���2��@�e!Ԭ'��Z;�z
�M!\�Ԏ��矹��������/��ꗾ�/I޺�����+�������[��5)j��SxG>f�S6/}���_|uw�K�W}r����7W�_~�O?���G�=���O����΃{}p{w�`o�c~]�?��ݳ͝�/�K�����ǟ<;��v�uo�=�ON?��/���v[c�[1��&�%�+�f3��1�͛��3��o�|@��7RV@���)JO�;'���h�Z]m�[�v�2ZUǈ8�!�G�^l�& �D�\�iȮ`FC�}.�^S�I��B���Ϲ�T0���^3���ȥ�^�T�L��Y9B�z-��i(v�3�H�r�T��+aYI���z'��P?W&�dZޤD��K$����B+X1�
2�'�����0ә.��$⊜�������!�R�Ւ�cR�^1�#�������+�z�2P�(u8����I���gq"��q���E&^����P��q�PeLD�p�R�Y��eT W�s8Ss)UchB�z|}4��0�Xr�go:Ȥ
.�]���D�͗����3��H
�嚂�!s.Bz�t8��fF�g弖A �ְ����-�6���\��R����^�,i����ټ��,k�@CR�h\����W�,���yzUUl�2J�06����Ii�p-[�
��g6�!�
�e�s�'�VC��׀��h����ٓY\�^`�)�3]lE��d/���.���P���GV*C[�"L�\�ˋ`,\KmAC o8�d�؆�)�����M�a�Iዂ��I���a���&�n!qK�J=kf��ZJ],2�Ql���lQ�����#ً��\<cM�^6�r�lu�'Sl���!o�T��22p�_�Hٓ�MW�R�
�0L*�0f�\����jٕǦ���\_I\��z��h���=g��y�E.�^;��g�K�/|rb�)�.WC�%�Ψ�?���9N&C�I��\J�x�%�)u^4^H��fw	�70����>9�����\=�Q��S��"s2�JAs΢X^�R�A�h6�a�#����;�Y�m�BE�.�>�z�����>^�1[g��'˰�=e��I���o��9�%K����1��)@��R�
5���f�LA�Y;i���~Q��13V�3[��ڏW�o���7�V�/7ZT{_��sj�_�~t�W5}A�=�\�mK;H����>������߳T��z��/F�|���v�<_q�>�2򛁋�������N����k*���3���<�5��w�"���W��>Z�����^���J��y�P6����Q��uXd����N�#���@A�ݖ֯��/k������ݫ�g�/��r��������὇/=8:���=<y����턳�ե�q���go�N/W~Yӭwk���-�4��l��e=�::�#d9�zL�bc��8��c��A�Ɛ%��@�A�fs�ʧ�����@!�4^�;%�B*�EM��
���akl�u�4���>7�H=�^�R��&;ԗi�"���E���=���7��VF��h��{$j�p������O��eb�7�i:g<\�t�E���0�Qa����BY��	eD/�@�����]�Z �������At!�hӯ���#��"������d�����,�X����J�X}!΅�&��&�-g�h*��<A�-�JL��_�H����B���@�8��!AC
BL9�>���!���y��O�W��_�z���.���eT�����ǲ|���wg9)g贛�n`��%\�@+ ��8�Ԛk��Ȁ�,~kn�qp�F!mWd 2P� ʐZ��pF�i��!ל;��j5�6Y6_���#p�:=DU&n��YjS$�И����˷��iyk������ѣ�lH�ZmJ2����,ITJH�B`T1��`��*� �&X��K�p�����s�͞�g?]��k�����������͝cw�8=��}�t�X?q�.������{������_��W����������+��y�G:?�ċ���������ٍ[�{���8ؼ��Bn�l_�|��/w�p)���ˏ�Q������`���Wm�`v��֚��2܊��1�-EHd���ɕ20�ZM2�l@�Q {=ELjy=�hԳB�\�e;:pSӪg�x�ri�(��(�#���B0���l-4;ҾD#hCJ�1�	I�5$�I��<�;�O�F"�M_ٞ�e�-�A����1�*AV'q:\�V���h�p���җ�-�D�G�,�-vxk�)0WR���k}5���2���ӯB80Y���R��l�<e�hp��1�oq��1/d=��^�E�W������4�)�E�2,���z�&B���Re��륣��B�tZo�|?#��    IDAT���A/��ٓ2�1��S]J�OT�L��n��{?�j��B������(����w=����JК#��"4�l��Ԡ�����)°����w��Q�ZL��T�Ǳ`�dwP �D
�6T�MR��b�����gX"	�=��Aֽ�J�]e�?�<ת�mڷ�f̌a���O?��K�/@�%B�B��Hc@��v�����%ϙώo��fK�k�g=�Yk<�	���!��ͥU b��D�o):(������G|�>::8\a{y�}}�=<�L�m?/r{���s�D���\�ҩG�l��//܎�A<;�Ǟ�p��g�������_��������{v�+�}��C�R����S�뜻��y~��Sm���[?���l������o=}��W-}������o?}��ci|���B���=�*�
�v93j�Z.C;��:�>CR=W+��X4�8>��S�rH���M����V����\^�
�9D�eIX:C�_8#��x5�V8��م��1{,^�	"�,�s*p�+c�2��Z�f8k�$ $��f�E5SfSf��l8e������0"D3,J�r��/6>0��I��VM.^�Tn�m;C�q6�i�xP%l�V��ÅT^I�yF�Y�j�WC�
�ո�Mc��8Z"�V�g�t�]u"�]�u�[��'�IA�g.�F��a����d�$��aTfv�BBhb�z͆���*W=W�	Ԓ����$6r�ö���T��C�Ȣ:V����>�	,u:l�iW�\-ee�A��I��q�n� si�#��$�`=&�|c��iX��'�U^��y�Dq�Aa���x[۔3���2����'y�H�\�)04�Ճ ��\�D�Ac�hEe�+�pa����2��{곉��B��3���-`�T��[1)�!U�ƴER�QZ�q�9`�0&�V K��dÑ�A���%��_U4!ZdCd�%hl�2�?�K�W/v��b���x)�h�D�D���;.ᆢ ن�a�'C���9_WQ�q6E
��Z����Fk�*{20Ն�IW�Rs����ĿDFS0&����@}�9����ZReWȦl!Ml[ꇧ��c���.Տ�Z�i��U��
Z�z ¬$W!�Ҟ#��E�� h�Y*B�j+�!���=��\���d4D�L�\����7dk�8Bؖk�ƖJ!2�|}aN��Q��rҁ�D����X�~&�P+jʶ�8ӠY�ʀO�Xx{~5L5�/M�X|̩��V ����M<[O'��1�1�b�'���h��7,P����Y�H���!�B��>����࣍@:��U9>/5�Z�Wd�|�!蓜^S-}�d�Ϫ2�$R�\I����ۉ�a�+MH�a�j�W
�����c�(��ajh8����Q#�}����v��f�����,w��;�����wP�}���%E���7Yn�o�N�{TƇ?gcƵ̕��z�76:�*�gʺ`�K?����{K�
̎�3^�y������+��˻�q1o\j��Z�1������� �Q���
a9�c����N��`��C���nW?E�,�_%�ҧ뇴�e��nܦy{q�5�Y��h�F%;�7n[�>�{��u�֯��{F�z�~<�ˮ�Z�X�����۠�5(�����(��F�!�j�eӍ������mq[�Kυ�e/M�����|�~��@)ʞ�@Mj�Lz #���5!���� B/�A�Vx����*���˘>Y ��Vxd�����Rc W�1��6�Dp�S�P��9��������N�ɟ���{�'�h�:����G��s*�K�N���B��Y؋�&�hi�U˅i�A��ʫB�"!t��'b��e3�7�E
�傓B�K��bx���t��%%]|H����K�B<N�|��GJ��c�@\�˳|]�LVU��8Bd�g���͘^�(}
-rL��Cjh�z4=p���ҟ��YT[��UE��ed[��64Z�.�[K
w�Υ����a%�155Xa./m'�E�S�D`h�a�$�S�{�@����ͭ�*G����)�!&c֌#D��J�X����h���VH兓me�-�b*f��٘��f�|!�����- [�*��e E��E�L BR24B|���2Tf�X�Ĭ�p��;�8��;֗Bتwe��;�x��h�[n���Z�����#�s��v=��,�����^�������V�qQ�ΡEm&��7�����{_y��������?������g�=^���݇��#�޽]>�lݞ<:�X��j;���g~z�xgou����7^�?����OL��*ƏY�:���f�n��E0���g���j-#r�/j���!�d�!b����Є�H��A�t4Q�!m,!R@S��Ѐb��DB�~��@���z AጱK<<x���a��p�pI��@|�>��"ĆꝬ�,�(��H�	Q �9}�p.C�+ն��H�W��d�j��'��oF�4�4ʚ!e."�3)�a^/�4�*ė�(
"�����'�-$}^����+#�>>���CT`
���Ճ(�fd���3Ae�R,;�m�2*��lj��65���#�hb5+�ق[:�,���Փ��L��Jݹ����/�K��\2Z�kvT�%)W=�{���7 C=BLJ�[���9�
�^���Z�zH��P1�z�jhȆ�6C���+�!P:)-C� 3�P#��HRb�*�(4�y��Ij�`����+&8SChbjR�se�JaD��!#��vHT_���O�y��7������������������]��q�ڥ����x���ފV�c'/��ۇ����������~����Wg��7�_}�>��w�������~z���?��'o����'*y����f���������ӛ���?{���r�Q�#�v�=~�;��OoN\]��}�a0��c���e���X�l��g[.����m ��uxa؇�����9~-{.D�d�[��?����j�,ְ��ͅL�t��	jH\������.oR�@=P�)pz�Cb�!��M����W�/���3��*��!�r�S�0=���ǡ���N^HK��V�4�	�������1�H�)U:&P�dG�68q:�)�ڇfMȌ��|˶�06�L��B��s~U�̘��*�4�dTFC"8"CJa�&�K���ci��cZy�v�:B��+�W�$�C�a���5�H_+\�!o���>W�t�lD|��P��������gأ��d�/W�xuZ4��"�ed�S+E+�WCK�YO-0}�DZ=6�/c����!D������
���\���ְa4}���.d�CF�1�W��
Â7�ְa
��;5�LM\�,���Z��@!!�sC��<C�C�Y3�J�����a8��z�l
�z
zmf�C
�%����䂔�M�X8D��٢6is���pF!)�g�hl"M0�^�n֓�D$2����6�͋k�HV��~�끅ó�K��+����b�ZK�>[�tC�ܠ��6j�����(F�C
�N�-�
fE���
���3���.M6PF4��2�s�79b��S�ђ-]᝹�9/����!� FQ��VodY4U!p��9	i�dO�2�!&��@}HFًu`Ǭ¹�� ���\U�\z �tl�]��kā�!c������e�E,>B�p
���f^
1K���7�D2�K�R�b��Y4ߦCG8/��0��cOc�I� �l��e�����e�W�^�^�S8�6"�VR^4C�M��k!�ڋ�TX.�)��gp�D���V�VZ�Z|x\�������T�^��{>S�Ig�0�D��-�r�U�T����Bp��h� ��n�	^�H����㒳OB�S�] WEV/DoŲ�D��@������Z��b�)��S�!+���g&��)Uǒ��¸Is���%=�u����Z��<L�f�W=��G��q:ׇe�P?�3�7{�Ѱr��g�����ͭ#�f��H@�q���Pઐ�ֻ~A����h������x��:�핻��;ɻq-s\!{�s�����9yA[�w�x ���y<��{�U��.q"<xv���j�!3_�.V�g9��2+����4y������1#���|��������[����)ۓji�u+��×Z��(yYy�X�����es��L����vh�}�3�X:['�B�!cB�4�s�N}V2cV��YU���!��g��Y�ȴ�3/�"�J'�!��p ��*H|�f5hj�@p�ђ�*M�0�����W�����fV�謡{lܱ�낓SI���i�D��#Oe{�sI�����d���Z�B^���KKT�z��m�٬���Ȫ���)K���M.^�2�A����7�*I.;)C����&S��|�FV��b����%#M��u�I��F<���)kp��B��U`���8ZFjlF=פ	'��1WdL�z�p}۱�,�t�Is�b�#$N���fmm]�N��[RS�f٢�j�5�~;}K
Mv͆ʮ'%�!�M����U\�t�l-\T�h���KAa�� \Z�Z^.�D0����gf�&b�\�p�:��5�檹��I�������=Wםʗ�2�����!6��KM$ؒU�^+e�X5e(%�Q�;��Rse�w0��<�ݽ����/oT�яN;����(�e��ҽ�������l�q3��� �:�V�j����Or�@�,���PX��}�����������;)}q}~zyqvz��~�Mg��ҵԞ]�ک�4��m~���?	}�+I�e���g�g/]I�z��������v�Ŭ�<��3��I���|G����y��
�#8�pni�Ѹ�'&Y)��!d3(�,z_��Lps"�r͡��*�+��
�y�@��l�W��ؑx5����7�1�����Tuצ������ַ�|�{�����?�ۏ	
q^��zd��k�K���p��&d()��R8w�0l"��KD/#Ye0"�N ���+��g�x���9�2�*����8��R6�B)\8!�f骊 B�����l���(P/V��jg���l���dL�HC��ʋ�cR6�(R�[�B��>���-B.�i�x��T${V���$BA`�ު]������r�W��@�T>Gyw����0��l{�\s,0qW=���HQIj���bV����V�j!\� ��B5�6��p���Gf����H-��ZR�Je�B�����z:�s�s�h�����nJmHp2g%��%Yߐ/���+�&��Dw����'�+�c��wvϯ��U���%�?��3��+<NǓ��.]Ͼ�~|�V�CC���>�z�|������o�����7�~t�����O�.����ڷ~���~���g��<�?~�����ϟ~r��>Z�����.���o?����x�ŧ�?��={�[����{a�/��'�X+СC͚��8Z+֬۬-�iZ�f���}��*�LV��Бʺٷ�c^�^b@d��䤖�_|J)v�mxL}eC�˭�]z}���Zjzvk���ʢ�^^F�5C=\[��5#�!Ų�����tBIG��G�lX.|H�(��V8@������FNb�2�5x�����k���ײm\�f:�9/r�p�r-C�f(\c Df8����1��I���	"44SM~y��4l[O|j� 2�`�ы��oX�l�Dx��17Gy�l��X��@S`L��7oێWDK�y�_e�,��8K1�7�f:E1�åYX`S 2��3(e�z`|.�؁8R\�"Wd|���h��`"�By�f)C��p���Kä�'Gj�aS���
P2���q��BV ��lL�9�9�%�xe9#R�^"�p+��H�c�����z&_�����RL��eTX��b"�f]Us��W@�zR�M)H+�WTS(�!���E	�!r��Y3;rs�<�)��GPK����`�eX�!�0�JN�!|

���Z��Gcd�7dk�3�*�����H�jŦi���Sȕm꤬���i�Sȫ7)v�d�ұ[���^ �e��A����\ђUvF��C�����WZj��Zy�ل�)�y�s:�W~!X^=�㉙J
ie"ȋ3Efve��XRSЧ��t �¹�ˢ'RCH�2u�MR����;�)�n��b%-6�4,�^��y��b�b��CY���b����7��G�%�,�ىj���k����u��@[��0���`�Bx��V	�nȎ'����uj��K?0ي� >�����A�iU�1�pù �p ;����!��TO^��NQz�U�,{J��0գ�h�nqgu q�3PH5��M����G͐�J�6h�Hb'��5e��C��{�ᅷ{l
V��I�� d�i��畑 }�y�¹BА=��V�F3u�r�"x�Z�+�_�I��vt�S��[N��:��u��[W	�/��et_��s�~��`����ѡ�(}�v�yw|��y���������c?h���{/��u����y1?8v �_�[]q~�/i��H��<��~o,����h�TUo/{��Є��`|fsGX�?\��:��S�nI�q~�����O�G'�.O/�.���!z�a�����^���連�w{z��'�Z(���^�XL���[J��(#�rXh�5EtA�PT��-"��1�����6�ײ�&��:Hч��)���@��!z����r�)�0Z��l8Æh�/)<�٥^>C��4�͞�I�#���ǜv�&%I��/��B�&ȥ���͋�FӲ�-�������o��t��8��?�3��e����ĉ;��q�O��g�;7R@Y�[:}�LM����e�ضZd|��5�+�l�4����tZ���h��Rp�	N�%A)L�)h��2�w�=�l��cS#+�r٩\grq�yQg�M�P#����N�5q+�Ѭ*6�>0<c!~�сL�����R�3�Ų!�ٳ�KT"�UbX̙+CWL�!Z����*<[?���9�w�w�%�a߰��ܖ-��Aa�z�5��M�W}�h[+@I!c;�����m�ć#�Rj� �
��w%Ul�ɂ,��P�A��i���f���C���-���RHp�n"f�K��4���5��k5�kzѢ�G4�\�ۋg/'GB�by��ˤ��2Z�4�����`a_�v��a�-��3���ذ�G�V�Vps}��MRw��>�@d�훾�G�׫�m���X=;�u=�	裃��cǎ���f�N<x�����������xqzv��{޽;`�m׳�<Z֞�����do���ǻo�<6�s�}+�`���S��]y��_yD�ξi(h�/0���{�6����Vò ��!V;\O�E����6��E��R�7����+I/6Y�4hN�3E�)���>2�zT�U	�k����bK��U�Hj:.�؝\���A�!�ʳ����D�����q�NW��A�.&9�ry߲���G�Rإݐ��Y�R��DPm�"�*C`^+���"���琁��U1h��v�B4.)��M�p��(�5,c�
�&��Eͼ������P�R(�B����m��
��z� �04xu�>�$��h�D�V'N�F�l�@��[E�@�M
�0d p�J�lRz�"��%2�ZhJ�����8v*���X��Y1.������Qޖ�B�Dz��B��!.����(��[��Y�-#D;���
��R�i:�M6�4˫�5D`#�D&�#P`��ad�yf)f)�4L}��DCt) n%-��65H�x�����I<$�X�)�E��r��?��mz�<uf|\���c�/�C�����d>_�o/�g�W~c��do�����ݓG;~#��['GO?������g/��W;�x�o������ʫ������=�??�������x�?����)������ŞG�?vǯs����'�>x�ν'x+��k�[�ω�#�M�1A�����XC�a�ml�V�:�!�A�4{�    IDATn�����sy3,�C+fu��#JR)�l8�@.�5Q�^.Sc�mFۋ7<ACx�ç�fÉ��Gp0�6=��2Ģ������ �`C:��y�gF46=�!CꪭoR��C/|�p�f��D4ىVL8B�B
x�����E*W��&�u�ɨrF�֚��Bx���ጹ��1p��->�j�9#��^��
���%o��˫�*d�0�P�ȅ�k#ʰp�\�l�LSHR�.)�!z4�^�J���a3�c�y�k8ER�*�e4$�[�bg�� /�u���A��tz4�k��eώ�È̖��!�yI�SҐl�l�����!8\�\y��������P �ьrs����%�1��3Ԭ�אB^C�j��p|F��lHdCF޲4�)0��D�<�Ɩ+���ZŜ`.Cy�d 5�z���RR�Ε���o�l��@L�E1����P
��]5S�}�OG��B�
cc���yф�J*�@�6e�%/�B]C�r��)P�A��в+@x���]aCz7�h&�]1qd���]+P�2�1[y�錂^�)EeW��/i����
h�!U.D /���քOe��l�M�Dl"bd�'"���j� ��T�NV��>$)!��F������0�z��̂CdJ!��a�)p��G��NyJ�?�(����!M��!Wy�NML�)"L�YL
�@��)U? �Y�z����s�6rA4!5!zC���=͙N���=��(!�,4!U�5FSF`�T�7��3
M������9;�Փx!�7/6��cr�I
��$�S��" E�b�1���� ri������0;^��5,�~"Ȇ/}�"W�aL��[.-&W��b��!£��Lpr�6}v��h�Q�z^�������`k6�,�>�\��aR��ӢI��d�c��n !�6!WgQ��Z��\����/�(4=W۫2��Do��AP�(��83����	ǿ�{/E��Y����z�Z[�U@'f}~����u�����ys����IQ�ew�X��U֫m�)m�mτ}ع�w�s�n�ȑ�Y��������a��:�U:�jr���j��셛<]b\���put ��~_��|�sy��>����W����8N��GǑ�Y�� ��a}�φ��:���#*��V�͕�?��rK��r��M(\'>�^]��^��'}5�e�<�[no�Mv�:���\�]~1t��2�h�`ew���肥K�PІ��6��}&�-27%��0r�!6b}�5�ā�����s�Z�j��Π�K]l6�E�H�����!�I9
�׫V���`�ҕ.&�W3��Z[$�d"����`3���Q�͝�����O������ΐx����$��~�3_�v��Jڠ�i�񫟸f�������(hh�8Fٚh�r�1]Xu�P1��k�R��~I�\�͔�!>W���V�P0Ei�� ��H	��(@�Q�0�.�U!5^S��y [�թ�����-�b����aY���&�����!2V6����8�iȻ)�	Ԁ�8�U�׻D
��Bʅ,K[1��V�@�8���Vg-W�g����� Bf���FH���)n8	4ۂ�Q�ڸ��
�l=$���)R��L1�c��0�n�ً�(^Y�`h1)ۅ��-8�V��'��v�K���D���W�رZV��n�\>T��ө1%�UJ�W�&�-��wA(���Ψ�ۏוE������o���p����:={7~��׆Ɲ.��su}�h<����[NG��;}�vϓ�����������ӷ�~ϻ����/>����>���x��sr�2ծ�ң㽓����˻���|�ݶKn�m�ۦ�/�k��z�u���n��lS������������_(r��z���Z
Sc�!�OH:K�8�i�{d�V8o{^��8em&�Łh����ja36�����
�R8/p�F�|d����^-���X���k��m�� w��5H;X3��:J�뀔�G����X�h���w�]^�C��u�ڟ�����������YI��i�<_mrA4�6��Q��m���e3���(�-���8�l8���d1T��>�ea�8\3i5�%XT��L�����G�UUl���H��fS�$S+*BӑHܐ�Fы�eƌSyl�ZYp�@F�RФH�8�s��j6�^�f^	(#5�F��j������]�E�n�%�	�`���cb�����;GB\ GV�(|jՌ���&]Z�E��ןK�BE�oUIM�VLC�Z�=)!���M�a�\R���RD��E��h���d��j���jX[L�zM,����D�٫A?���E!~�g�HS��B�bD����n�WEﶮ�_z>�8��G�x�����[5}\�_�b�x|�?I-���6/�Ow�wN?�����^<߽<;�_����>�^�~���G���7������������/�>rx��|v�V��#�p��j��`�r��=7��s|�sp�������w�?:<���<ؿ���[;���W�њ�ǚ�=��25�6������z�\��}��a�����m�X��Ľ�n�)���Zm�t��o���p6�ض/p�0��	�,qrM��B)V��ͫzؐ���2�a��+g�<�Rc��N(��,��TH��	LDxU�1)TL��g���X!�5C�z��B�������M�a6pPoH�T�Ş���WP�a�zCr�e�*	A�8Ь�A��ى#h��|�4ӗ�m0�)"0���� ���8�&>����h��:��a�8C5�!
Hʰa �̫Ø�4q[H�Dئ/$>��S�2bF+��!4q^x�3�L�����JDfl��6�pEJ���A�H��q̐1�2&�P-}���+���ڐ5���(ʧ^CMU���ї:�p|6\�O�cX���*4d�Wv�t�J�_"�b��k�/�����-�p���b�Z)L�[�����h�̂����\e$)EU��*���b�S���tbt�	�i� $���a���h�gC̫p���U����Ѫ���R��'�|�n(#[���Ӊ��O��Q5ʼRWdF.=�R�S�����D�G慧fXC�kL
(аX+PF���}f�*5D��zL�62��=���
��g h���VO��'��P,���\�p�������P���u͹
$���>��0p4d.�͙� �e���+�Լ0����.Q5�8�i�H������1$ΎM�%�B�.S�d�G:�
��K}�����v�؊��������3��K��-0���*	P^��� ���f��Z�ʣ�9G�m"���-c�(d�bj�V�ܔ%�x�vj�1�UȠ_j6�\ު��l�=s�dx5�/J��ְYh��W��Τ�V�l��@Jb��n^�>�s�15S���g@�����Y��}°um#���В+����Ά�VUs@o�@DϖEl�l�^��Y�LT�pl�\m5ErA($�V	�,Yor{�s*ӷg퉅 �a}��>4Y� }����V㳧�۝��������L�� >@��Y�wz�;9�OY���`��ou�:O+�+;�����N�9�z�u�~����j}����Z������������ܺ�ٹ���='zw�?r���Q��7���!{�%[^�Hn���ꚩK��S�\��H�ٝ���K��:U;���y�;o���`���`���+_�\������kZ?ܸ��.�l/��]������^J3��W�W7�o�y<4�}GI��z�-�'�d�eoW�l�H�aWA�^dk.�TC�2}�(ż��]K��@�Ĳ��"�Cg��EQl-P���U�i�Ȼ)��Yx�~r�O�R�UN�#̤\��zR	�O������*9�����g�=(շ�����Hx߉w�����WF-R�N�9���p�pU+аu@��8�����RI9E���7�ey��z%���lq�p �3hl�S�h�4)4.6�&�(�Ƿ���[�Y���)�R�#��$
ΥK݁��N��*J�
��A�;_J͉w�uΙ6��������z�Z����
�'p�qͶ��(�[O ��\�b�l�VO�%*i�!�^�ɦ���ɚ�a5XI�@�O�4"#�͐d+ o�!l��6��%۞����ٚ(����zC��(vR��[R^��B}5� ��	��\����$r��O>q�"q�l^��^,^���4Qv$4CA�P��7��`�]��ԧ����O<n�l�oV�D/��I�l)MJ�K�B1�]����@��	�a~bs�H<��~}��b.I���>�wa_�����z���gk���!�^�n��u?J�������o��߸�����ן���η��N�{E_�I������;�6�n��7���W�����˫3?{{}u�	w��g#�W�x'P�y���_״�F�o��"ʙ� ZL룱�ٌ���e���� Z.4X���ೆB��1әvd�!5sy-�ꅍ����A:��Zv}����0D!����c[#�x4T�7��O���	�;J�����m��#���k_'B�˘��ogv�Ig��1m|L/���z�͎MS�V�������$%��~�����D���{���+���(|)��Z�*p�l."ZG�f���-i�ŗW�;�+��}Fyi�`c.��[���:����%�^�6�-� �~|�5�U���Y1>����Ԭ��^)���2�U�U�>A�.�?b�l*k7P���}�M���@�_��a"��?��\#��V�~�\�	z%�������o��SS���V�>I�Z���B��2r�L�a��0���2�"���ajhI�[%�^��H1*h(<0�K�o��Fz ���8[=l�l��!����s���m�*q��hW9\y+o#>z���j���o�[�w�z�3���S�zx��ۗ''��{��zv���~du�u������������o������_]����7ߺzt�t}wu����{}�����o�������uM�}��dO������ۗ�/���tX�����}�?�9�>����3�fdWd�H
���:���f�E�W�%j�~����~�V��"�@�K3�Ν�����3�Qղ�m�I�/��21+O���N_/����#�����VjiFC�ڋ��,��]�+�^R���-�@��72C�@-o}�E��E75�D�JbX%���\-{���JJj���J�G�d�׷4!�a����s�	�1'��k\s+�Sf �S�0��;H
����(*��(v5Ͼt��%Z�f^v��ĩN`�E�E(/��i)�*Uyqqb�24�6���g�5|��d�7i2�iR��
l}��m�a�Z�\7'������dy���)����2�Z4�U5]�35Ak5�7L89��rI�czZ�yg,��)�D)lrR�L!��o��J��bFӓ���]k^lL�=|�Sd2�Yv��GfG�3���pQ�1��WLv���N"�H�$��H���pC���S@�e���)�P[{s"\5;d����]"�z��55.E窰.WQ����5."hq���Qj���M��/o�t��h�5,o�%�ˈ�S�%���H0��CN�~J%�#Y"H �(CY��-�ye�F����A'WY)�Y�"�j��Z��N�y�D�����hB0�O�N�t"H��BQ�����ԋ��
�������+��ʎɕN�t6W[T�<B%��R?B.}�ȼ�hͮ�Dp�S�*޲��� �N5C�f�C��a ��9��I!@���&�B�ɟ��E��\" -u�s?R.^��L���J��!d��^��!�ؖ��@�����K���k����f�lҬ�����_��DӦ�S���9d���GckD&Θ�\
��nͥ`7�,R8&�9o��]�qx%��k�aҩx�8�m�9�V)&�'�9�q��^�̀L�Z)d�!�K,#~3��P1� ��+� Ef7#!����<�9Z�%����Y��ʨ6RpMZK�l�v�ݥ��{9ݩ9� �&�Ʋ<)����xN��hk��F�j����<Ϯ��=�N�O��}�������@���Iӥ�Վ��;�'�O�.o>?�;�8��$O����=<�D�Ջ�+o`�ٴ���9n�R_L^{.���ݛ�~���1}w�y������u����]���Q�s�^�,�5s���{��N�=��3J�=pRΑ�؍s���F�/�_�U���}i��qj9u9nryX�4O�G����V���� H�b���>�&�G^�Ϋ#�}���8ɦ@���� �'86��
bȅ�U=���Cf��!����P%\�I��s�l�K�h�e�ϩ!�D�YT�&�ƥ�&ȀpB!Z�L_s~úY4�0��/��yE/�?��?�������?t��"&N2;-�Q�uSp��H���q�Z[Dj|���֬9M���eȥl��PƪU[{B��l�B��ռ�
LP�LD1�\�շq��wԱ� ��r	�\,\3���I!"#X%ʆ@5���:��J���δ;Wov���'?�g"���IIT����ް�P�h8i�gsi���]��ye��ֳ79рU� r�I�5�SH���H�1���K^�B��^U!��W/��	lI'�E^����P3�WR=�( ��g���K�kcE#n�$A�
AӪ2+4d��Ӿ!�xFG\S�K��)C�^/6�hjzaJ��:�]�>p��>i%�u�oqM� ���	a@{���|�\����[�����=�`��Q�%��e/���4//OVwW供%{����{[��^/?;}�_$�>!�G�{ON���N��n��y���띋-_)8>ٿ����]��jur��*��{h�_�;xt��w}{���7�=
�a��������mo��뛳�g�k3�w�_g|kiu���:��{8�wm7�����;�1?�O�$��	i%�����cp�>h-~| ��)�!<5^C��Ky�ep�
R�Ȉ#�vl��qs�Bh�ϐTyt�����h��
�B)��H����yM�f�lj1=�[鱱�ҹ���K�q��g�u��ya�H��*��P?���}�{��{�|m���`*�YK�Ȩ�W��w��-�) 0�f��H�
6GH�/�!o"8�8��+2[c�C0�Ev=&�@Ǹ�1�l}�J�:� P+{ↅL��&�E�BJ �]B���pF����ցA_#h�Ya re�7D�K��^�ȵ>�� �I#^ C����Q����cpX��k����`s��2z�T��.�}�����iە� �,�k���R8
�k�.Ԭ	V��b0��3��K��Bq.�WF)0� 9AdN�!���0�Os��G��?z�5C��cB�wQ��T85!UU�^azk��b���ټ��B�S�pf�ğ�+��$^=^%@�+Y�E��]�~���r���{Ǐ�W[�>�l���w]���v������_�ֳrƳϽvw��y��[{�q��X{8������D�_lߟ^�����{�߮�n.}It��r������{o��x�����W�|����|�3��g�W��Ƚ�wW7O?��O�=���a�f�Ǧ��=O�ݹZ{�����f�M�h�lͼ�Nui^h��LpG?��?4�Lz[Ao)�{�g�!Bbz�@^���^�mG��;�(_ ��q�d4��o�����U�/㦔��%��GI�ZRl^�a
4��ª�0>�0$<�hp���8~ʁ���h�/��h&;3)��0ߙː7�p����&��:�-�(����X�H�H��P��@�
)�	�Ԛo�����#�y;�V�>Gc{S`+]v�&����ŋ7#CM:/j�`�:�UFQ��*LN!/��V ��狽�B�[�h�5njVO���,А �ސ�J���k8I��c
�������2�V��K$5ީ )])�����"[�p�a6��"VՐ�XF�!���!�Jd�/���܌p�d���a�ŖN�8��N�٥� "�pC��s��h�N\�p�r�z�k����v-�    IDATU�o�F����Y�J��F+�����`�o� �\�����!����W`�(3�jBq�O�����e�
��Ǆ0�H���B�>4�XO�@8#ފ�XF|��*8')Q����f%E��$rA�E%۰>5^���N�@�&K��3
\R�@����Ŗ���g��:f�*R����̛�!PlY
��&M���A�5A��S�:���!3;\ B�� ���9�l���N�'q�L�ԛ���U�9"�W8����35^
� ω��
A�k�b���O��1�+�M�J���k���n�G�lV�+</e=8�9�3��R��H.����T9��oe�4Q�lR�&�	���=��9B4�z���xS��')Ws)�X�!/[��48Z3el�ϫ�l�M�M�ά$�MK���k�Z��ɄT!5U��K���A-;5C:�Ϙ�i2"��)��.H4���>�X����ܠ�
׳E���m_�
�5���R���2�B$�(h���� ��ٞ����.�PT`6\1�H���5������:��k�Γ������T9�4m�q^��M�4}hu����V���ˋm?i�޽�W#yv]�|�s�%�K�{+�5���Ⱥ��3�g��C�$��;X�=l]_�>������%��R�;/����;���\=���zx>N׭�⥙�mq�'ƶֻ�w[��X��Z�~l˝+k;�䉷ξ�8.�:/삣�;N�-?s�j�f=�S���\'�W~��!ʹ������������8��(�'�=�Co�.����~��j������z�.��f�8ŧ.'<~pmZ����W�"���ٚ[p�6+��M��2��p�4�j�ȶi�l}`4�n�P�4ò�� �\.FR��@�5'�)ps�ЇBdƴK�ooL�D��hIaB���씛�u`���>pG��^N#��_���R�Y����4]��w�D�%���DֹV��� ��֋R.}g�2"��\j�ZLMl[�����6��P�3�jC�����*5S��XFe���Q9L���+ʰ"Ѭ�Ճ+�+Wj@G��*[a��2u8�2����#N�{|][��C7^�h�>��pRR�l@UNNF5�����S-�Lİ�0�hJ2)J���ͤħ�a������V�լ��_
^�aIea������fH��lwbW�싵��b�zzL���m�l �!�l�1m2�,�v
*��a_j"�H"�4�)�͉�Z8�N�#P/Ď�M
�H,}�ש��^h��
�M����g�s
�P1em�HЋ�%�VJ��
��f��������q	ӟbc���{,w^�%X�M�sn��W�+s�N�k����]� Ư�ۺs�s�.ʷ�9y�+�'�>�Y�~tu|�����a���x�&Z��=�WW�ޮ����/Q{���ՅG�n�����ĝx���z��=`v,��y���x���/���[�ã뽗�O��;A���e.c�1)׀���^�[=�`[j��MG���V�����Y7�)��9�(L�F���JGOG�[�C�!l���k�\h1᪪�#�f�joQ	CS6'�"���:�]Fd{�t�L���Cz&�Gx��k�B��Tk�MHo'jpiӶ��f8����Z�W�:�C\�b#��J�%Qj���Hj���G��(\���&�j��^�E!lS�w'&��DFX,\C���6Ԅ1�(����,o/IL�h2���W��&�,B=��m����d��J
���5"��+�"�d�&�t�nSj�����2~Q��i@L�p8��S�����D.7J�]�n��l��>�ohR���[a6�?�|G��.��ʂ϶i|#I��|�;~�U��*��fT����Z����,��5&А��'�L㤉�+2�L�>��F\�O�YX`��\�Z@v�f^`���i�ⴽү�٫as�6U^˖]`M�p���nn/����u���i�7۷��'Ǉ���˳ӛ����}�ҷZ�_�����磣��O��O������o�����W��sv�o�����������A�n�;��쭎����t����������'o?���ͯ>����<���������������~��~������~{�x�p�|_�n�#�8�i�6���i���9�l�!ZȀtK���@4G9�r����M��i��S����^p�ʓ"®0���`i�)�b���)Kdz�D&�
�'CD�eQ�J�D�����5����	2����1ʹ��C��qdфke1d�#��6_R��7C�I����@�k�oH��ʁ���!
CX
�Oar��8B��D���������Ux��T���a��G(���5�Sކ��hm������*a���2T�-��k�P`LY�;f�f`��ٌf�@�3[�����2_6oyŔ���h\@M������ϥ�k�2�#3�PRC���!Ǘ�{�.���
I_ߤ�@aj���S�<d��j�I["|�$���H:�<�����z�y����ij�Rj����!C�Eг�~��v��L>�M���Йd�\�@�}���5�L-CU��6��7	�2#ע=�)c��	�sa�����2�qRƌ���b��7,j�2ʫ�]��ú�PH�����_�0��U��n�TQ�l\!(�2$
��,�72�N��n�f��@�x�Q�eMφ�eW��hs8��T�:��!�@��l���劶8_�\���� t(cC�Q�8SgX��>#[Ͱş%����^��0.|^%E���1/E�h�����Yć�An�	�2������!<�t�z�(�f��@4☦� �By�w�,��1�R,�fdCƦ>����yhSd&�Ф�S3�t3v3Q�f��KSM`C��Z�8M:`F��S.o�Df:Q�q��(��F����x���iwbT||[
�����ZY�h)�V^db�E��ah(�2ح$�@��1���(��KR@�p6��D#f�����9iᅰ+69��U�R���N�������Z��ң��8"�f3�|Vb7D>_�e��"�jSYvC�'(��a��)��Қ�t���QK�~I5^����t̅�%�'Π�j��M �M��<z�oi�������s��|6�7�g�>\�ZI�]v�$�����ː{߹8��q���]����+�Q9��]��~����/}�������j��t�fl��]�+�yv��1�CQoo�'�ݣ�?�n�=�`;%��n,�4Y�:l�)wW���1~��G#/x0�ci����;.�;~��w��Ѷ�E��//w�ػ\_�'�g���o�me�Mve��������5WG�[�o{��(�b���n�$������V�E��ld��4�f�*��l#��Z[G���Oj,��
��)�����&�f�����q�yN����g�D�T�^+u|伆!3�j��+�i��I��Vl�!�g��%��!M�(�DljN�������y6G5��%�[.k��E��$����;�� ���������Q��*^t�H�ɢ�d(�֓e8���^��v*}���9�dV[�
��6�r� �@��h
��Ra4��1#�� 5MUѸi
�U�up R����B\��-�Ω���YV�:�Ⱥ��!	�8=��~�i���)��CY��֜�&�������I�C��#K&�,�h�h?����vL�62��1��4q2�t�2�+�75=NQ�՞L��)�E) $��+C��ܼ 5���ڲ.�Vf� !z�����eΨ`F�UF�u{�=���:�i�Bp�5�������9AT��DBJF/';k�F�hy�F���-+��'��"ME#Hl�]u0��)�R��r���ݵ-0P���(ǆ_��kOS��O*��^��������{|y�B�ݭ�7��|��])�׷��?�����ϗ:{�^=�x|r���v�_�^�}��]�W���w�z�ݯ��B�~�n~�	w�f�ͼм���ˬ<$86��XS��{o��d�tǿ�߲��,�f���l�Z!`B�&bq���,��${�34!��c�-/�)�+}�,/Ya鰋�HGmE�O$\����EZ"��`)�2��p�)`/�R#�������nKj�@.��+�=���K­��ݔ�%>�۶��ʓ���-{G�lg��/	q��¤�B��tfvd�^T�]��$�*aC� k!�+;e�)Dï��AYPx�j�@G���&������B���9��D���bB(Д����h3��N.�R@�Z�[*��BR��'�P�l�hԸ��A��jX(�*^����5��I����}@����1�)�*�r�&�[�?e��%�iv]��J���c���������f3��r����[�A�uS5�r���Z
�������i�M�7~�9):����Im��5�Bg&�Ӱ,�h�z�r��Z1�69���l
�����0�#gW����+�a�����@�i�_�8�]QO����;���������'�x�͇~���v�%�gOO�|��9<�E��������g�����R�.:����������7������_��ͽ�q~��pptx�w��,�=�����|��/�w��ߜ�������}rr����������9���?��?�/�ίO�vO��ݞ�=r�Ռ��|�B&hj��'�l.G-��'�1}��]�vu��|{5A��1�j���Z��EƄh�Gk�Sj�ᢴ��%ի�E�b�=Pc�����1�
�&��0��R�"D�/<}�����Q3[��"t�����^jC�LH�@)�x+u(.����_K�(4.@��fZ�5i��k�5�8�*�&�,��4e���h����eg�'�К�, �Z������z�^�;ɦ`ض���L��Fan#5� 3��&>�,B����^=����ON�!�BO�0Zjm&�f,�V��B0Ρ:�����]�Ĺ46��7�ҩgp�O������p�_����=Ipf���'͖�-�ѣ��p��?���þV�nXq�fuKꡪ�������g��~nFw�ε�^{g�@�� �p�"@�� Z��p�Bxg��%�jK����@�$���vށ�C��yS+�z��`A��0D[&���RϘHx��5L=m�5��_� �IF,���r!��S�6LC�g�ڲ�pd��=�!ߘW��W[�~#�E�e��_�FA�G���r�6a�+r|��4$�	�=�C��_���Ƌ�H���px�XxsI_lCF^��o��;L8�g�B����+�ʋ��lRb)���#)N�A�p�ѷ�!ͫ�A6NC}�z4�K]����-/~Π)u^��pRN�є1�Ik�H��Z+�RT�X"�lj���)D����#���5��0�-\yz��7�P��fp���f�M
`8��C��*�A.�^��[��"1���R�Z�z��ر��=O����1�5�4��N�![�N���L�������@��a_�1�)���/[_�i5���z��@�@�6�-&�HWv!���e�7�ڰy�c�Z����mrR��T�D��%e�mg�["=��n(p��n�2�W#˖w0q4$�0r �nѼ�������vC}���1�̥��1����Krl�枬��t�4�4^�k��0��:W��
��5�)![���Ď�<��@�j�-E���!.��Tֻ�%_2�;&���⪟VY�����/e�v\�\��X��M�{���p������9�{��뇥�t�V4}8��O��{�w�Ș�����k_���]�Ow)ƕ��7�����n��¤��t:�w`,�k�N�=�N)�t5ӓ���t�~7�eX��'E�o�,����O�L�6/�4ki��z�������y9]?���t��O�<���r�3����+�˝���������K�t1}؞­��E��������%�����I��U�`�{J���az�Dv(�G�`yk��G��@`�d�KgH�o�Eqi���`W@>��_urU �px�ɨ��A�&[j�V
.C^�\���+N=Z3*DlLd�9~U���[s��{ b�8�N��������4���3��ׯ~�+��QpJY%��'���i��21�s!X^�&��Q|�\�V���lR�B��XH)TRD���Ɩ����b�/�F�N ��˴&��&�F�0q��jc��RS�jy5������ `���.�;�d�s�~h�y'�DQf�[j�T]�����f�m��j�ǐ�Ȟ)O80��x[���8�Ɛt�J��'��sA�~|4�,��M!��sY%�Ú����b1���@0���U�p�iv�""x.65�yU���h�� \M'��)7ܞoy�[�z���w)��Hh�!M��6�8�ţ�\ �f;�Z(W�1!���c���?�9����9=��CZ&n���J�5ԉ=�$���DQ�2=Ȯ�� �Q��g=}�̱�g�o����2n��5�����Nk�x��7�_?�ٛ~���w>>�����[�]^,�N}��a�7�;�����^�\����s�~��+��N=ן��{�p�z���ǫͩ�y�×C�V'W�S�������7�^�_}�O�뷗�}�hz��u��ỹ�Gx���)�]k�6q��i��m��*­U�c�+�eL��[��ɰ�m�d����o+����`� r.�]T6Z�����pȢ��2/0��8�◴UUv:��ྷnO��9���.ϕ
�� ^���E�=9Ld}���!W9����eN��'M�DhZ[
8���4���T0x��	r�,�@��k�
=^E�$��������z|��=�p[��&�'�

з2�hzKl5
jb��ф@��Q..�k�Z�ly��V�C�i&�StD���9� ���u�"3���E�MM#�1��&M.���]�澩�R�\B8�j(��6����~ɻ���o����M�"+���Y��~���~������j�ꯉe𦖡�����1Z1:���\�
�e�2
O�0d�u
�n��$�?p�x'�G�;J����hSֹ��h�Q-��Rc�r"Ss�Z.�&�/j�z���l�2��b���w��Ow����|��o�����/~��g^�W˫�Gx�s7���Gg�����?}��~v����v�w�]����x��ч�y�㏟�o������l�C��>}�e����{p����˳ӗNHܽ��Zz�-��������W�>.��ȋ�/��t�o���3�mS�[�\.g��K�2�+1-�(���[7=rF�l�rmi����y-�^v=|$[�y8`�B�L��p�@F0FaU�n�Eh��jKMIc}B�5��I���(ϐ�����C!oCv�3��Ha�fH�*�X���b��2�ۡ�ո:h�%�9�4�a�,ѨmWB�C�ˮT�ͫ�p�0�1#f��oK^|}�"��
ɥ�x)�y)��g�iVs|��
l{T>C� �AP��q" )k6#�Բ���j��c�q�W ���+��z^s�k�PS�]�LY_������-;0����۴&8�7}"p���(�!�ʅ Ǫ���b��i�p�,rE.cŌ�q*&�mf�2L0Bu�peP�\���R����rIV�&Ȁ�	L6�t"Sch@QM���ː>���k��� $��{|Շ�<z̑�ib�	��5�N��Q8����A��5��
T��_Kj�c�!��ER�U|Lh�`8f5#��+f�j��:ٖ�0��!���F[%�h�h&Pm���F��,��@�!�ʋ��x��FM�R�8q�D�"�� ����;d1KM��GM8N4:�+�aR�z��0�P�l鸀M-�p���T��J�`��MS�B� q��p
� /\ fx���)�\U���p���%�%��HpD�7�#�IBj��Z=�+��V�=�� ��)�M����4k`͐���3�������B��m'�Zʓ���У�f�)*e/���!��\>��nU��m��򊢦��d�
������z�h8���HZ`�t�&�n���%E    IDAT(�k pv��Ǧ v��&>j�$�+���@=�!2���ц+����%{R�F`5���'Ny$bht�B}��F��v2��%bM��2���YUi�-u"y��g��`L�KT�R���їEI�ǥ5[�0MQ�E5Q�����e���9#���Z04�s�i�Z������b��f7&ڬW�+?�⎲�iE]��r6���}�N��w��7����n}}�γ&���Z�����h��b:fs��rKYw֛�:���p��M�;�ǿj�����������~���V�N���z:���E����s�{����0~��[jߘ�e�ydRӗ'�.���*�y��ک1S��,�i�9,�_�Ae�Ѥ|rvz���w�v�B�V��e��W���gw������޵;��n�{�l�5s}��Mrww|��Ե��i�g���y��S���m��qW�))jtѴ�Ȇ�tpm����h�H�����P��͆��h�B�l:�ӑ�9 ��q�p�3ن#Q��C�lg ��粙��|.�Tm;��|����	�������|���j��������K>����C^m�\T5�E�m��Y�n��<�b�!P,N��ep��*$�hr����wThj�Z�eOJ1��M�?M�tNH�v��oj
hQ=Ye�i^h�yR@x��ќJ
�;�f�Kv^k�1��\p��+��z���,r�zM
�5
;Nޙ5u����!�VH|���$��p���\�\��xI'\_a��c�T��L��;��\�uq�7��M�b�U�!Sh=�l���,�!&\#����!؉tǥ
�z��+������cq�� �^!�p4�Y�6�\��e��$`����~�-$Щx"�oS�,]�b����
���,8�o_:�ϧ��$����C����,DV����2D������f8�����{?�^w|U��V�rbx�NW����<�W���g����Oz�����Ƨ����^޿�Y�o�������On[z�������g���;���m�7���KW5oެw���N��ݺ�[��oov^~���J��իK�p�W��L�c�^,�hv��v����|����e:�'�5K�[�i��m��Ŝ�b^+�hO�3�i���zrՐ���!�����K��w	��\��z.���h���qHE���&MI��#p��5�a��;av5�}j=�g֎kQ�(K
��p[W%v������{0��I�5d����G�ESO���VH�%r�<H<K-����hB�(:� K�,@�&�	�J/h�c�1��ӄ3���B�ȕ�F�Y���r1Ȏ�^]��Ģ	�����3����0�e�G�4��)7A�\�MY:���B�8�EM��vRz`�R�7ejڰi�J���F��R�=�@��J �5ѓ"�}*䳹!�h-�F�54_���G�����g��MD�&��ҩ�/5WLC�	2 -W��pC����O!}�c�m
)��D���U�b(�k1I�q��RF�g�Eв�2���-�y�űV8\Z.F"5C��M����������`���hs}燜���qc�_�<��/q����������?]����3�n��;�/>���|q~���Սj������C��1�����S�}�v��w�?ۿ雔~�����iN�{���9�D����o��_�{��Ã���ko���wq{��/~��p��_���;�?{����_�������}jv�ndX������ˑ5M��l{�ǢY��h����h��д\e�L6}|GA�W� |+l�fh����>���:����(H(
� ��eG�-�^A!��#���!ŢieIG���p���$�]�1�ݞ��<~��,�C"�@��BF��3B���5R�5�k\4y�W[��ë<���1������1���˰�\���#e{`FNd[?2e��4v���
ۮ��\S̻�3�-Wy��M3��`2��r鵊�k��h� 6��Bؐ�	~CJ`��i�R�W	CHQ§
�=�Q� "�����ؼ�~�M��^D�hX�P��
��Ւ��a�K�Ly�F+�4M6���
�p$bԪ�!��Mk���WH�^���� �-� ��A(�كîN�X1I!�2��B�l�pC��IUC4�@vRz��iF�ksIĐ�^�RTy��F6$2{,B�ŖT��1��0#�#3�BȪ�a�H�!�GTL�f��p�\@�����(i�~�^F�(`LH$#&���!q(��I!�P�RC���>Zd��v'�oq�:������D�Ȟ�MH�|E��mW|C6�dh��fO2*��);D[�l�a�E��,$�j�20�-�f���8��-V����,��������-);�٦�BZF6�,2�2&�VFFj�2X���K�7~ʃW��E@֓R�s�[`��Gm��u�(_cg�5��06���URI�ȼh-N�.:�0[�@�tx��Rc�#0�V$���pQ>[R�>c��
l�\�	�̦�QP1����;nv-v�$���m�Ѫ<\�&�UbL��J�S:���ү�RC�r! �-i	i�W[l�Sc�%�(2��V,��6jޖm
�Iq�1� �:KT^.m���T"\`����оMs��
 �����N��#x��]����$śxu6G�([ �	�s5"!8t
�h\�)�ǳ���,�8NG���a=�!(\�<�I�,�d�2������s�Ho�⥹�Z�������;u��}�'�5������7,=m���L�?�)����qÄ\��e}�c®o>N�_	;8�	bs_yK�9:�~2}E����c�'���}��U��ao�:Q���̰��s�FӷN�^:���'1y���na�1��F�x����+�j��].o���������.}�eg��������ή���
�ژ�{N���v��Z�iu}Mh�26�e�0u�,5A�i��g'��a7ꩤ��>C�G߁N�(�6�=���$U�D�6�"�.���"F.��Zj��I��Z!�EC8}���F��·6fle��f�rAj���~�e�eD&"G�1k��|Y��6ז���ї�\���t���3�N�Vm^|�b�ҥ��NA�ӂ4��["s4d�j(�����E`���޼l'�&K!k"�/f c
�x�q%[:�����!�fv�.�T�D��\pU)Co548��S+)4��@3$+�R���)C�O[7QcDpB.���`�ae�#QQ�+M65�@��!n)�
ɕ].�Vx�)��E�����s�O�\���h~h�����caۢs�t�C����ޚ["�MUD�%�7���=O�'k/�;"�:&PO�\*q*n
tdq�m���n?@EA�&oj@Q����*�Jx�I���L���u��>�=`��[7�ʅR����ܻ�*d�K]��������K�t���YQ\R2�ٝ�K�&ي�դW.D,[�P���9)x1�V�����L��f��)��>�^C�~�����N�p���/5�u�o�|���o?�SdV����=;~�����g���^��o�����{�'|��?���>>8Z�R���3�D݁�+ӳ#B Y@�����}t�⽳���ic.NN��7hv�w~���d��uӧ��vw��/�z��<|��W9���}ȇvLm~A���o�Fk�R4O�i��ֶŌ�3�����8��!X��ҳ)�m^�iw��D �#���8�8��F!�q����P.�T��H�ھ�'���T�,��������C%�r��P�IJ`��rJ���MS�\UXm'8�Q>�&��Y�C��A���O3C,���M'/>Da���aS�S�R`B��'�D:����q��)�+qjZy!c�B�m�s��%U02��2N�2�ԩ�ݦ����X[m�p.6�����\z��K�k8����لxN�+�p�4�jfP@�c��NS����=��d�@�iE���k��p�y���o�R�E��g�< ��YF��H��իV�qM��T�z�a'5����5���͛��l�1��|�*)#���A���#<;�UF�"�6@6Y���t�5e��[m�Z�f�K��ώ/.���Ͽڹ|�^�oo���Gg��.��9}������W��x�|�ÏwO�^�������g��={����+���W_>\/��Z=,��?����.�}�N {���b�9��~�:�]���߽��?~�|x���o>��_�o<�ݜ���OO��]��[\]_|��_��W__�m�����w_���읞wW����l'��ޑ+`��_��!�<��@͖ôJzC4���V�e�h���ڼ�lȫ�B�ޡ������q�wB�"5�V��q�"����e��a��>���B!��J��r �a6P�sLA/�	Ƭ��h�k@^`�����'��!o���#
�"y����'U���%��G�6��D8Nʌ\�he�M�a�%ec�1����! Xaȥ3,VFF�����(�a���>GLH̼��`�|-YFS�*)�	4�#���a�k��as1Ԋe�Q���$[�^:�p8[Ϯf!��ڤ���y*q>�p�A�@+*��06�@5;���#�(0��F ZL��\l`��B�Z���L�.
��l��
q"d����ņ���:�������#�I��S�eW�v��8t��	�5C����p.���S�ZR��8����E�n
��*��O�\���� ���#���8b��ڶr�e�hU�����>/�v%%RiHX�l�!�5I�kL
��2B�(=D��=2�o����0�(�=j3� ����x!EM+�z��)d���G+�p�b�V��whV'2�=JB��2r�R�Np ��!��d3����ZQt���!��{� #*oH3ʖN���=`�2�� {�BĂ�1K*���1�2
�b��Z"��BR f28�#�o�Bj@����}!۴A��`^�_yI!��E���f�K�Cǰ6==��C�R@4dH�!�T�!NCH-���#h�d��?H�pe$�ɫ�^�4!�l�M�g��h�#�B|<�Ja���!��
�2{�qD�4�\��q`����Rv`IC��5gx�6pkb}��Ԓ�Ŷ���m�pJT1*R	��~ZIü4d+?�ћ?�2�Ǟ?�)�쌑���D�b��� U��м��,1�9�S���e�&��S}��H�^:5�i����h\!����|"�:��Vae�9�d�S��kB��=5�]q��}~�̊��݃�vk�z:-��^��^�8���eǇU�<�K�V�W<\�^j	��9���w�����]w*:u=����ͤ6��
�6��(.v\L>t#L?�t���秇Gb�ur|��(.(���{�r�]���*y�ȯӯ��7�:�w������ӌ �|7�5�黕���h��_�l����O�����s��N�k�N7/�����=?������ÜWo_��ϫ���z�����&�^ަؙ�p��+��oIk��˂3�:���!P��ޣ,C�7�s��Vؐ�Ysd{ju~ߦ��4���$f屽Ow��.b�?��
���fV�vIM��irᳵhz^��\��B�5���քoKN-�hc�$"�aw�Ϲ�_������������|�s����cH�z�琲xLY�$����Se$[m��e�S�@�iVS�����:����ԦɎ���N�a�(�њ�XI{�z\�4�!��l:)�)5�V<����G��!�fC&�j(��D5C���b	:Md�ZO�;X�f��#Xꦏc�UR[`!��05̡Y����kߙS�)ٜ���1�J��pd4^�1��T)��������uA��2:���b�Xs��׿����֙������Y�Y'o
t��I�� Ԕ�d�2�\CSTIc����AC��	���C�*�-�g'��cS"�E���"YC˅cS�rQ��w�p�jJL��j��Z)��b�l_�!��J�U��Y>+(}ߧ�W���	n���nw�+��3b1�V"H� ;^��W�i)׾�zrx�1|�~�����_,�����G�G�^��o���}��ŕ���]�뗋�~�{���ó�����==~~~~ws�����s?p��wx��?;==��x}sq����]o/�\�z}�9�=i_�?+���������t���My��V���if�i��l�b�_�Po#��zڈBr�5\)�'��z��V��CQ����
4��*�N��QR�|#�ʛWU��],���)��
a�_/���<[���F.8���'���<�1�oO��#ߋ�����G?�)Q�J��eH�ᡢ`Yd4sTMO��&��BZ�!�IY�D�,6S�^5'�n=�ZG�t\-�J��	��Z���Q0)Q��!��*���#"�YX
̑�,4��3��R(��&qs���a��%��p-����m�-�AG#b�W����3^0��JS�+)u2&0��zG���
�g0�ɞ4�C�2d�������X1s�)#}���g��!S�,J�!����ܔ�)��e�B�yS��S�(�j��������iF3婣�١�gDF(V �~����\�B*�R��U%��զ���]����� ��5�k��^��=��}��ޜ�|y�sv�vu{7���;<x�١ɜ�}���9<y~����No���o?:;>�qvp�GG������\���������������ݛח�;�﹈��U�鳟�_><>?{�x-���so��./.��������ݛW��7n�����EgQ�h2qs����6;C����|ͽ��l+�zrC�x�0�[��a34�?����G(�0:F�	w���ˆk�1$�3��d80BӇW3��]T��*�͋�Hv�NQ���C��/���@HF��3�Z�4�2�U;@L�6�M���)$/;o�V���ALv���0( �X!�#BRh�3dGS�آp�^3,o�^+�p�,��F�b�cW�M��e5囧	L���le7�I�ݑ��pU�`�(�2CR8���i�pCx`����X����jQ��Fcs��������+f�B���chIeA��3��]%�l-#o4��P3�U�C�!b�� �!��w��%^��H����Q͢��8���9�6�������mX3�Q�:;�����IM`6��H���q|3F���V
���Pv}��^�i"�<!�5��!#�Ͱ"���W3�Ԋʫ�\� �{���M?�UlL}۠u(jJ���U�\�\b�
�Z=�Ƌ&���t�b�(����r���N�	���+�2p�2��j��~*��&��b7�b�[�GRFd�$�
�ԤC�b3Rc� �#d��qU W&B�����8��i������p�ϋ�Z�J�Y��Qy�E��a�a+�B�����H"� �KĐQ�G.v���[x�!��x��ư:���Uh���R�-�Pn8���J��!$o�%˦�k��������1��1�E�)��}^�h坂��i�R�pU��G��G�����5:Z5�'���;��3�MP+]ϫ�b��p�1|���W����Qy���f���[I�C�в��7C���p�:�l�q2R؎-5�*�6V�`�G�\lj@�$Rd W����h85^�@={dQ���2����t�>�.��ȅ�Z7�w.h��Ψ�J��t�g���!)�1� b3 �+���� �͂�,�ed��r�bL�;�(	AHL�EA\Ó>��%H�7o�o�����r����W'w]ּt�����<黐~�ũY�ǵ8���9�����d��⺨��/�Kŗ'�8��<�|���O���覴���t:u�R��>��|��7�;{�랊�
�O`���f5��5E�+�0��ݽ���龴.��-�)���?��+�������ݥ�.mǮ�zL�������"Mk�;������Pg��������\)x�3]�U�t���M�x����8��n���w���}2/��m}�=�a!���K�h�p��]S�    IDAT��x2�������Y�ސ@��bB�D��b@0�z�[,��![��!l�o�r55xY� ��+q�&]F�#/S�+{�y}/���ؾ-�駟Z�?�񏾑�t�In��W�D\�@�å���*�)8�҉e Z}Y#��:3I�&�:4d��J�5��Y��ZRD�U)$BQe����rU*;�thl�!Y�6�ā��W��&�7eQ1���g�)t���g�}�i�5�����R`3�{����F^C��'����4�G�&��-�˂��;���GyśE.��v��!Ǥ�7�E����:��@z��Z8�b:@%�=M�Tj�@�l=�s�fH�n�/Ό=u��sie�B"UH��-$�ƱƧ��u��%^ۼ���欻XFӷ��P���4���D.s����?���r'����%�Qr��O4���š�0��1��K��!=��F���&�t������Wb���L����ɳ�g���Ƿ���<�}{��������<ۣp{vr��5n�~�v�&�����?�?�]�zu�:������7��/o�O�>����p��K�Y./7��6�/_����s�������������绷__��-}Dȃ\�
�g����U���13��g�y���1�p�l'޼�;��y�m�l��Z4:.6/&���7����T"���@-��F��i�hȕ6��1D������/WL:�)$�m�e�U )�XI6�?5<oze�!���n��e�1\���o+ʖ��^�����=6�����\D<\y�8�6��o�pЄ����Ǽ��z���2�'��n����@
�Fh�\4� �8!B�B�$e�	�2YQVI�C��	QM�N�!��2Vd+9p����zL�)���SjQ�B���z��W��e8}C��w�v�}v���R�8�rUjj�f�Ѭ��e�Q�wQӞa�3���t���&��P��}�����O~��h*�+L�/�ՆWy�ja�eA�?�m(Jk"\�Zv�S���m}����Lm� �����2��5C̑��R����VY��bëh�Q�WBKG���3�&�ʗ{+7�xt��@v����(�����j�������?����_���G����Ol����=sys�姐ӳ��w�t/������ק��tuv�8>�v����{>(s~�jy������n/.|������ɩ/^��zy{x�|�p����~�̷5.ݜ}u�����rwy�x{�g=�6���K�x���Vkb
�G����j������x��t�����!OY =/NY�[�I}nt�������*���A�J���ei84GN�0M�ڦd�^��S�Ç]��D&�����ʁ�D2J�7�Z���6=��a�6Rj�t� ^.^H=p�j��G:��!Y�z����
aT!5C�����IqD�N��ň�H|�y�/�-�7#}:D4�D�j�◱E��U.Y�m��-Be�s�)E^�DЪ��i5%�4~Y�3��BY
^F�R�g����t qFQXd��M�є�َ��6JB�/\�.M���ʨG�9��ކ�󍤭��4�!�@��,>�8Z�8)20�YI�B��8cF)ā�T'�&���4W�����c��	�O�]� �!�Kk�l����*B\��] #��4�i�}�D3�\�[��pi���H�p�=/�� �=ȘM�X^�6���058#}�!W`�z����Z�� `���5��ҡ%b��p)�K+�p�h��b�o�
G0�U�>��\��
�'�H�Z�CX�)�KH���`������hy�*&d� 0Ax��fa(C�F���0LA8Z6c&NK�UR�eG�̫5��9�K��W�F&�1����`;���j��+o�0�.j��0[x�(�(��#N�Q��Аq���Cؘz
�#7}�RNx�\�(��g�ifg�b�M_U!���+�\����F+6W��V���V���)�Ր�����ZH�E�њ�(�S�޼0G�7=r^�d1SH8�%/��R(*���I��H9���@&����\pL�+<A��>���3�2A�fᢴ�JCj,D8�t� I�aF+���CJ?���\q�@C����� ����<>�Z)��4�0!lgJ���ʫ�7��Ι�7쨵�l>���@=\S*�D(�tm����`(WC�R�ѧ�>)g������@�@\�������t>�e1�X�׮knܸ��`N7�]/]t�u�����}N&��f���^��N�)�`�/\>�T?}� �>�uL�_�ܱD�;�1:�v�@b�q�[��"�iOg�Ι�f��0��vszl5ޮ�ܳ�|?ӎ]���b�����Ogzc�1�_�<�,��k�6��^�`�_�ܙ�H�v�����w:�u�������{����{��lVK+W�w6�fv�w4���]�^�uv}o���T��~N�9}+t�]���ʒz�pt:.d2:�mL�t,�Ê�9|����zǴa��M��+�����(�nw	��(;�Ѵ�#� �8�~��ڨ����uz�j�D�@Z��@L�t�p���l�z�@d3;c�ِ���E_�t-͉>�T��fl�t����ट��>�
�'B��A���K3")�����Fk�!��TU.yeG�T#]6&�&�H�W C"}�s�r�5�R�=�k�+�@8&<~�1L�PK͹w`�UO{F�)(���X����	U^+O�U+'f�\�h����(8�)�����cX?���b��d�)�T`R�����c�BZa�h�c}x1!z-Mx���«����=�,�Y[@�ie,�u0��2&<)�(���UI�7��rQ�kJ5 ��EyT���`y��$˦������֨�IRaC�!�\���")�'mf׿��6fͶ�2J�V��e��j�և�,ھ/Ye���b�ړ[L%2a�b��K_��3�u�̻��`P����u�qS�/9v�FzX��ρ<76���x4�B>��LW��Wק;�7o/��	|�x�̻盓������c������������G�����n��{�/~����>��}�5�,\#�<�xI������拋������|����α���/��_��~�t��#��� �z������g罰y}�o�;��y_��N]�b5�y�OC�@Z@dH�v���A,#q��0��lQ��~ ��\rr�A#�n=��H�H�<\Hi�htC"p��!}3
IvxG%��}%�t\��կ~�f
�Zٽ��yO�2j\v�+�����S���R�j�h&����=�.�;�����VF�B:���06���J�	
D#WyI)�!ca�Q�U1d	�{K3�������2;)�a�Bx�/�rA�W��:�jh��S(�2$}��b����5e��B�얥��B?�o
��3�ojz�  ٚ#�F����]����pq���4e"��"��V�Ǎ��)Rs�F��K���.�Ӧ��3�����7^S�@;p��fhp4d�.q�6� B�� ��f��1O�A���eȎDI�6��!�H�ҥ#;/$~����Z}KW%4�X"Bj	"�B��eB�ا�yY�AcczsFd�xᛕ�ݛ�߷���r��{�����W�7w����������϶��g>S��b�ƇVw��9�Ծwt�|��nu��� 6�_�{��|��������>:~��m�>
/�/��7�o����W���/���������$nOO�O\!uW�ǳ��˝��������x�w������=qܤ��t�S� faǚ�Y[�fǰm���N�ķ\�h�z�*1�)ɫaB�6��a1,�����h�U�7�H��,=�(kA�Po�L9�6cfM��=mG�WUՏS�a�m�*V�S�R&aT�eR�r�o{�㔢X��0j�r�!\���D�>�FUb�D Cm�l8N�q*�1�����WC6ox ���9G?u1�pv�&0YF�)���)�M?\ϥ1�%�b��)�Ӱ9�DN��0��B"i�yŦ,E��a��y����Q+P""C�����:�p�m��2*g�2�3�ƌ�C(��EfT����g�m� $��URC��R�9b��G�Q��B�(����*��K�h���OJ�{RJ!١o�
͋ͥU!�r�1�Vp
�\!�)�NQ��"������	�k��/Đ+H.�@�!���7�b�&!I�NjE�b�Z�V
`�D.6q!�7ZRU��J�z.����
C�����+�X�0�X�ڔ��\)�!��6�Ԉ�lXI�� qx��R�5�9����F�FF.���L�:�\h2����mF�c^	�)�7��!W���U)�j�&��=
3����IY7.��Ua`��~!@�d���2u��;)�0��d.������!bS�W!NkHSl�l�) �A����� g����*�Q��ϛ�a
�l�QCj�m�����VF�����(x+�H�@ĚU�3���� ��[�᭛	r�����P���!�M� BD��QP:�!�Q��C��[Iz�SC�̫�&Ŏ&<>[�ف�\�B�B��U�^�aH�����Pv�-۰���Bs[�Y�.!*C?��zR3<�a�Xx��`T[. &Dc`�=F�!���@����9���S���҉S!���s�;����wʮy������Ͻ�r�`�@T�U�˕�j�Tl ���'�]5!%V�B�x��d�{K��4��Xv=/�"!�!.6����[�kr�*�f����t��q�`��r��:��p��:���Z�M�Ü~�r��tQ�O�8��Գ��9꺧�㞯��?{yR��,|ӯV�6���b8�)��uK"��3u$�ݭ���*u��a����uJ�o���3�{�>���ͦ��r�j�w���yX��Ow��=��4��Y����{�����w\<]/�:���*����D���_�6n��G?WKv�7o�^�^wo������?pvg9�>wڥ��;M�<�Z��1MuZ��߫��cWL��n�Q����MG��C��1�9��ݫ|��U )C��\l`%�2R����\e�3F^á3�S��=d4:��q�'��~и0��PK|�
o[�*ˎO�#�7���ǻ/u9���g���=�zO hֶ��p-�s�j��j�F,��%�l��:�fQh\��+��G�YH!���2�u�#�=�z:o�N���R�P�!�f��l'��S�3MH:�Q��B��\z�Iy�c�Ĳ�bB�wO;g����y�v�_�ͽ��f��5�\�B� �q����"������nR@FQ���1�%�>$>;W��a=�іì����8z.���a��[4
�hlL=ZQf�V���%_��[�X��^:���kFUeې������v�bkp6}
�D�AlCC��*�����k� ����}Z@;�2�ǝ�+8JP���_@�
�o̳*G�K/%P=&��f!"GӷL8Ѧ�G/���%w�����p��@ǫ�O�xP{X?0Wk/(+��7�^�n�o����dy}|����x��|q��ŭ�����������^|��:?xo�xx�㣕�
���j7��������Oַw9Z���
7�_?n�����6X�_\�������
}�h�g%�WJ{��ڧ?B�cfsL��>�4]����jML�ݰ�k�-�~p������'�=g���G�#+���T):.�Bڴ��I�7���~�I!��e��R%pMx��ƗN^x4	�2|��O>�4��k����S %c�+O���yظ�e���&;�>[�?@����K��!�H��V#2�X�!��q�����{�\.T�(���Jek撁֪
gSG����4^��׊j�22�����L��fQMj��J�"�����!ӏ��9(�z������� m�O��@�(g�VOJ�\��w)��Y�˕i�);vbe)D1��*w�|��̨�vy����N%q�e_uS�������Hަ���M�\�`�*6�;YÁ�d˨o�l-W��8�*�`&��y�x��/*r|=f!%e�c�F�38$¨v�o:�9���,h���rb��N���s����,��w0O�}��w��<N��?88�[^?\�nn^����3��|��g�>��X-��~s�\�����n�'�f�-�N�֏���Ճ�n���jws��&�W�m��?���^~����۫�W��^?m�t�]܋������O�=;:��k�p�%������뻫K�i��+��{��S�+����K��r9-��YU;�sW������P@s�{8�'���J�#�G#��:CO�e��Բ�gt��{�����kX��Q���#0�dD�4�A�J �-C�Q^xr;p(3�<~"���2R`�#���S�. �ebZ^H��-�2B:`/�@��F�kq�-�t�p��bp��+���fn�ӯE(E������p���/A����p���-Q D�T`��m:���h�2�8	����@�ehX�4��	���;B=�"+�"�h^�2 f���o4D��Y8���7~G��2�f�G3m����wP0q�UC�G���Q@.])����x��&ΨH`I��B [^�!��Vy� 3Bd�¨H�V%1�V?�sۨ*�$E��DFl�\�Jj���t2�Z��Z�0{�f�*�~[.c��"W�"�S�@�z��i���1$�l\����UI�1���0и%2dWj��U=p-MS��#٣�#�Z"�2
�h2�4����z��\������ll���	��Z��������Y�\%5,N�y# �ŁC&���(��Em)v�\�P��\y����J���ke,]�8��e����Ԋ���O��DF�C����^ [ao��Kİg�0z(1��`B�4��f*I��"g��PC�Óe�L�w��b�@�^�p�F:Y^^��&�w���x�(�r�h=<͑�p���GT�����-�F�ʘ~.U���м�Gfh	�,Z���#ԧ�OsT�-�IGcT�z��3��Hm�xB�­\yi깴�b8�(XH
���ܐQaz��7C�k�˰����,0>\1&8DF:6o��.����lL!Z=Y-GOaR�A
��ʮw��u���:�8!��W�¥p��G��i�{���U�T���s�@޶.��������IY����3056WH46�T�<8����*�X"�a�le+ ���eG�΀��ד��3|sz��+%�?{�Fi'G�I��Ӓ�O�Z\Wg^;nH=�]o���\��M{�����{+�f卶s�ӯQ>����Y�CW]��j��p��s�����N]�K߉��.��Y?X�}_���d�X*lzp{�>/�|1��vN!N#���V�;ݺݒ{���N�$��)ℯ��-ܓ�oe:r����?���7�Y_�uï=_*��ݺ�낁�
<<,��wW�{o:��掚����+���[[��c�}8 \F�s�O��犌f'�5��"Q�b"k@��W ��Q"L������	a����:h\!HA=�1��~�ђ�ׄhB�0�5.|C}v�
�jay�Ph\@Rz�F~�����o���?���w��䡍)��~"z|��!��NkŨ��q��Mm������_�#��D������&;�p5L�8�=c�w:��qiM��@�\B��#VcTq|�6!4e�Zgx��,!fīW'�����s�Δ����r���qi�39�i.I�/E}��W ��~����Dё�bRe8r2>��p��i�X��*D1�צ��6_��12S���S�b�D��z�hʹa��pR����Yv4^6���zGAU� �)s��Ԑ_�!)HQԴ�	gcF����Qcg�bWg�^y�%���� ��m��A����=��:����U�K?���F�wv�K�k�V�y*�ǳR���F�J���Z%�j�Mm{��JOo^���X/k�N站��� ����i�^Q�8�}�U %    IDATss���x��3������}�l||X��{|��}������/����������������a�8ݽ[]oV��z���z��b�z|{q}p��qu���:Z,�OwwV7w7���@�7=_���z�޵Lo}�)�i7�X���ҕ�!9g�w��=��u�h�"'��ƞ�<�z�5�:�]������9�%v,2��m�E��23��ybN���jm���MD �����5l���<����E|�
�l��H����~��_�����A=}�s� ��؞"]����?��~�{�#�U}W��=��+C��Z|ف9v�Go�zZ�7�# ��`�r,4���ԉ�d�[�R�sQ��5��!�2�)WOj�p��lO��#;.E5��6�E
CF6ܤ("k����2Zj��l� h&U�z�x�����q��� S����ȢY^�q��D\z��
��IJ�!���:L^Jَ��~�xN�T	�2T(/��#�M%�s�YQO��S����Xa��,eL��@c`j��z|5�o��^`LvC:����M_���I�UvU�&5�R��
��3<=��C�H�#����*��Uf�����f4Rp9�����-��>;>���gQ�>����o?<9te}y}y����������__�Y{c��c�k���O�������{g/����i���{����7�����^/�o׷˕�5������݇�=[u���y�?��~�w?Y<�-�����ׯn�v6w>Pc)V����>��p��ʓ�O�z�����h5pL��g���`��54Y�P�i),Tk�� ���b �-����b��C����\�75y�Ơ�C9�b��"*�QK$D�A0;��@��t�8>��a��Oj�)*�>&�X.�]�F�Z4�?qC�!�>d�\!��5���1��Q�i��h�[�8Eɋ�UUb�j���A�X:%J�>�Ȉ׶9������Y_j��J<~�1q�?�S��H
-ن�r��� �~���T��,E�CǊ�S���/��@�kH�&cԓf��Q�j�%���Y�*�W>WQ�ٚ��1��N����J�@vx�Snv���)5��r)�g�!zLͬ���&$�z1�FQzx�3�0���ӋA�aʭ$q���GH돀_�`ag�-e=o:q�W�����&����^kA���(Cm̨zRŠ�Ǒ�D�B?2���!�#�����K�˰��I��`d^F}�pJM!~��d��\�R��XC�4;�Z����D2:�ْ��°7���$��8��aؐ�(`�2�ů�\���p�4��5��W˥o���JV��X�p!� ��u�/^U3<�N��/����Ze�ʛ��WLp�hs�D�;�M����Ta��$5���!e��0x5x��c��Uj������>^KΈ��Uv���j�|3*#/Y�v NSf q��-q=2��͎x��5����s�bznI!�����c��(`̥ز�&���2*/��7`�%e7=BL��Q��Fal=CԤ�� !�&Ȩ��DXx�#����7�&��U�i�)!C�-Dy������z�
N�:#�d��rd�u�yc9���P�$~R뢿��6�;�#��J7mj���d�֔U9`
����g:��[�����^{��!�D�P��S�.�d�k8��/G/&5�L'�7�z�L���V5ޢ
4,�Z+V��1���\�����Z�.��'.�t�w��˘N���I���M��;���]��	�E�R�E�!�3x�qy��p3�K=�i��*F(�wUI	$7ı���RN�p&�!J��Dh��8E�'�i��l�x��i8��R�ln}��-C�����������W9����A�ھkZ.��S��qy���{}t|{0޳Z�q�su�9G��{�e�q�]􃃕��������˷��/�� {��;�������H�=�֣��c��W"��wG���q�<�l�?����
�]���+���sU��eeLʍTo����ʸY뾬�Le<|�x�N�ō;�����f�vߓh�0�e�����Ҽ~����j�O���_n��3wQ����/N�>|�m���ˍ)�~�/#�F6�[pCa��r}T�l!Z6/[l"z���f�
�l�!��l}+�NUu!�]Q�Œ��e^�;Qz-Zy��K�V�ؤ4dC�#�^ę��_�̅S����� ��O�?M^�˼~��/�����`g��c���X��ղx��cV,Y�֜`W��.Ͷ��T�XU��C��UE�BSp�\��T�!���J�@6�DUD��MJ����W�FSo��1����+D+DϦ�	�rI�Kφ[O:�JdW[�Y(�i�5��k���5��?���(�
h�D�,]Y�dK!#&�P�)#2��i�g�4�:lY"p�@��6�2����4%5sы�_��v�٦)
���L�E���-���Ŋ�,�z��Y�Y���/�>~�C�1䝋�������a"�s���HS�*4�m+7)��oU�^:{�\�K������2*���f��&������A��L��Z!V�b�A/q4�B*�/ʖ�c8��/<��汙�]і�">`��=r9׏W���_�^�0��Aw1�E����C<�^�V;���ON�ח�Izq�D�zp|�����js���7ח�q���?w߿z��>|���g�����������������������Ϋ�v�s	vv]���۬ﮯή|�ǫ8�6��;�9��tLA�m!v����˲D���Z�8����18�2:YLe�ֳ!�0���:\8�H�4�@�I.�C��1�Y6�05�2DԒmLn�7dW���V�9���O�qcɞ� j\N��M���d�)��I֟�\�O��o~�� B��!��[^!�dvc����VG޼�����gC����{f!eadSk�dұ�$C.�i.�ɫ�i"hH)��IŇ(hX�b�5ԛ�
��m!ͷ�4���ar���P��S���֊-J��0�Ext@�r�t��I�,�P�\��o�J$�/���t��m�~�o)��X�ʁ���������a��Q�R�L���NCIx�������dy�*�@}L��f�VU���pB��@v�Z����siՓ��0d�@���U.<�#
��Y�ȅ�ـ�bF��Y��҄�g�Y�|�fS/|ܻ޽��8�>���zk�O��9ݻ8�asw��������O��ڹ���7W�~�������q��)]ﾺ�;�����f��n���敧�lVwg���������Ϫn.v���8��_�.�n�6�������Ϟ���|������/��ƻ)�,>�쾼���ɇﻋz����l��<l�;��x��J٭�	��	Z�֧ukWas�r��U��bq0k��H���ΙN����@��m����j�
�GV�?\�D�pJ��>	D ��	�"�R�fv��^| �Q�޲ e\%͠�;3��B:�t�U'�XL.�B2 \Z/�6]�\}50&���R��P��E��m#�T����1��/b�壒��b�R#\��,��M� %R�@�Wy��8x�������2�BC-A=�BB��f�u�)�J
��B�-���7W|�F��G�;�p�-�¢��ׂ4)D@�M8�_��b�HǮ~� C@��9A6B}�����@����lE&;�"�Ψ�Y�Όh��I��~���k�G���ɶK���
a4eS���'����Yҙ����r�D�$�b�\��ËUqQ)H����~��Di!�)�5w��j�Ld�cjb�h���I0)���(��h�
���,]Y�s�:��[H�>�~�W
���
���	��()��j�s,�za3
�:� ʘH��)��=g�la;�&9��_l`�Q;C5C �(��"�����056q�h�����x4���	
Ԕmh[̹fI_/*�&5����zx1��,	.���9�"p!$��N�YϤ�p�ߐ��E����	Ξ�� RD����ר-�*�j!l��@Lj	
䂠e3�x'�A�ƥ7�mgc�5Ԛ{�
Id��\H�D�x��l��u���f��i�=8�:y��!%�7dk�	1��R�b{�[���k:B&���&��1�#�1j3o�����HGd�/�z#�p��!y)LMxHjj˘/�8��Tf����fM�!��Y|�L����e���Z~��b��sӏP$\�@4:�ܻ ��&S��60͙���+�e�$��m���'�S��NA|���I��>�Ȑ�+0�rٟ;ᷪ�:p�*M����qʚ�fь�N�U��2j��x!���Ԑ!qإ�s�*B��V�z�zF��Ś䊃���eX�����+�7��:���R��������.7+/�����7��硬a뾧�����D��q��ݵ�W~3�������W�|����S��|�s{�����g����������o�w]�����v}��Y��tC�cl�<��ƍNŽ�?P�Y~js�ȏi�;�I�b9�%7!��ZL��il�?��������ы��^^��_u5�b���]���g{f�-�/��\
V��F�3�5���۫�n��?*l�k���6�%�d���Ҷ���Z��g�q��I�l�C�vW\f��(C�ƶ����K��K�َ.ͭ�DD�bN!Y�rM��f��W0�(|~s��g �(�ʥ��,���qڇ�A��Z�BZ�J�7}_Z��O�|�E`���]?t,;��my����,R��lM�y��XEc�Te60\oj�!&����f�i�qh:�ȮQ/WjBZ%�Yi� ����`��G�炐-V�ټ�	�Ѐ���R���@�,q����R1+ch������}��&�Bp���K\Y���&";�������(i�1d�窏���Z2�Y�*_�Fy3"S�/W
�C�QCHuZw�}�(D�,)fä��I�孤2Ƈ� d4��0&����r^��.$�RKWv|�VR��R���2�[Uz����	+E�Თ:N�ldGÎ�l���\<�͞��{��Pt�����4*D�j"j�ZӠ%�����B��'���0�b����M��6#��*�X}��Y����ʶ3d>^�<�����/9�8�뫻��ݟ��O��ǇWϿ����|���/�����3�;��k?�>|������ɮG��<z��=gN������{�;��^~���G�~z�K7�>�ھ��y3��ystwu}w�5�K�]�j{9�Ni�v?+��G�3�2w����s�j��g̵bh������mm�#���Z���e(�H!����H���@�R�d����CRf�^���,);r�،�y5C�q���q�\ߎT1��t|�ҩ���{�N�vh��К8]����H]p�\E���Ȏ%�z��@�Tl� d�^���A��HS�蠆�&Z�R��w(ɛ��%�f\/im�p+������2��Dy�ND4C=)��C�N[�:�F��@�8A4^!�N�_����J�^�)�`N.S��C!&Rv!u���A�Df�������I��%����@�r*�w��G
�p�#U.��������A�x�e�|jF(�������!5=$2C��2Wd��ټ��Bk� 3Z�-p�L��0[_�B�Z�\���h�μl��
f��G�-0YR4����.boN�4H����`�C��,������ࣴ�7/7g�~��K���������ӏ<�������N�=�裟��|{}u�����F;�[���l=4�v�7*�{���<�}tt����˛��괷�ٿ������vW~d�d��6��Nv��$���{�y}������ۗ<|���Ϯ���������o�/'����?�r������g�5p|�u�/ƅl��\aM:���-#�ܭ�Yc6�%ʎ���UE�����b"C�rQ��h0d����WR����aj�?l��"����P�^x:�#aԪ�-����U�`Q�҄W-���6�#ܐK���c���@=A���bg`"��jheg�5
՟B�m��9���
�SKj�34T<BE[Ҕ�j�8@}�\���{���2�p_��	Id�!�x�k�C4;�:�l.}4�hI����a8(fl��pDxcΌ�Cn9�	V|de\�#�a�Gn�%cE���7CH�a3�6�0"�m��s�l��^.�]��D� ��� 8z��T0&ٌ*�m�I\� I\B!�Db[�*�/o�E�����8Ǟ�'>[S�>#ڬ�1��f��224`"�%�&�����]�N���ן��>�y��"#��?������p"KЛ��P���Pԏ�Y*o�ڬVU4:-2���y�%*��N}x}Cd�� EUF��8��šl��2[yp�b�D����H��#TpL����4m2�>Ğ/\_�P_�aL.��&P�'eHa��!PAK��B8B�_�c�s�|�J,f�C�d��[+8�F�,*�3y�Z%�Xv�M��M��2$f��<F�@�VT�Ԭ!̶��_CL4
�U`H5�b3� D+�!0�Ѭy�Ӭ�9��݃��Z`{�L�ԏ�5!��9A`!�c�\I�F�L���b�P`"s��� X�J���gH�KG��T|����L�X�R 2$W�³Ñ'�>�n��I"��0��}��f�2�bk��8�����&�Z���F
X�gT Y�@��ː���a�X�>�2�y���2BF�%K \K\�3Ɇ	��	fD�gh��	���23.�K6�5�NХ ׈��f"�:��H!�U��4�K85�5˅���G ˖k會f�%ݔ�рD.�� ��괁�Iqɥ7^�K�ҁ��	�(KM*�W��Gh(����qaM�D��#_K%���?��v��񻖣<�$ٺm)�1��εٗ�����gº��z��uI?�9���`�ķv�"����#{��Un���v��&]��?�vs�>t�r�{_ļ=8�_�T�:�{��N.���?O=r���e�zW������b�/o��?:B�t�ֽO�u|��՞�t�~�����飇�z���6~�l}�>�����7�w.2��z��ݵ�����pH�QO_D]��Ȳ/��+֛����.�,T��ʳ�9{l�e��i۱�D���P[�cC�0�6[�
������[j������O?���N{N�_��҉�и5LQ�I1�ū-�7�4yU�VD��@��rH��OZs���;�4�l����w+��'SB�q";��¾�mMxKa?��h�	�E�c}�����_����T��T5�
ٙ�ࢢ����Ȏb�֊u�vSa���8�J4�GU@�i�ɪ��
c�l��#��S"��b+�`��	�hd�ZS���~�k5��3�[��C��I�!�"�$��k�U� \�Gm�[%B lds��o��59DJ]�;�������c c2��Ue[�;n�?c�B���Ω�s%nh/���G"E4=�!�&���)�1Z���FIeG�H:��ZQZ4N�z:����Gm���W�Od;a)���J M5�ʢyh|i�%ʆ�񕍿gg�r�C�	fH`�6�jҷ�w`�q�TS���4'��go���g)�^hJV�����W���`��o,Ğ�>�s�y�o��������������N�g2�����4.o������{N�o���8x=�|��ç���}ԋǏl������w�_}��ȏ�=~w����k��������=�?�؜{��j{s�뚾5�ڰx�|�F�ZioO6�	����2�q���[� �a"����ؘ����F+��P�sY�7��%��� [�-�,�Ն�[:�d#O���ٌ������ة��svE�-6$Ӱ�9S`䤊jÌ�l{��bݝ�կ~g7S�]Q��'�&V�����#�kW
�DT�Qko_B�+oJ�8���I����� s��z:z�f�� {K ��S �U%%��[��&>��j&.�P�6������k�:�#�-<4    IDAT	�ԋ�#0� ��pT2����Mo�ЪA��MG��!��;/#�@ؚ#�k�R��Ԝ�*5�̢$�z�[�~0�v7�����^H"�'J��Y_K��D?��O�}ꦦZ��]�b���PMFS���ZxLF���\��U�fjA��P3d�]<�1˥�p��Ȭ�:�&���j�U�%[���£UyT3N.�Z����h��+`zg.�u�Ps0b
�lR�������������47�ۧ'�~�����/<K�'{N��O���޻{(�������w���v����4��|s�w��������m��=��]���ꫳ�>s���έ��<y���V��ݳ��G��99:��ϳ��۫���ѓ���O��M/m>�svv��+������i���~� v�5�f��������i�k�� �!�5�"C�5R8�yF1x�HP����'���v4�1�)c�"jz����� !��9�R��G�d8eC��s���kȥ� +���@=h��d+߰��
�lM�Vf�A,�!��*�d��R�ܛ?��I@�h�j���SFx�;C��\�6t�G��'�����׋�C��k
��ū�q�7���2�O29)X%�ec6G�@�(��Z�V��ԁ�S(���Ϫ��#�!N�vݶ�a���B!�WX�j�e�M��.m�DK!�zL��R�d����=�
��@��dEEK���r�[gQ�l�"�(*����kB�͂/K�Q��e���cH�b���5��aIg.!�-��z��v�y��
�f,A.��ұ�&Φ��`v�jk�z��&����	,$�a"��Q<A4�J�s�!����Ѐ8�2����C3��lhZ��y�U�R!xqJ7{<~I�T��j�����3���(k�g�UI
���s%!d��5��k��I5�~�(W$B�����a�[�l��"� �5��*>��q1�8u-T^=o4v
�м֫o���P3�*~�o
�Na���l.̒�@f�t���
�	�8�1����s�hͷ,3]�t��Wrh �¯vd}�6C�3	���Q�20qx���f26�V/`�SG�����~�3�\��Kd���k)|Է�E�R��a�a�^���f�ђ����8�0�8���ǯȅ5h𶝾�L����e�J���E(]���3�^/&[k�
�%5�Iq�[jṦC��O�����!#��KZmD�ɴ?#�V �bMM�`ء90����2D`k�H���+��$C
��!)�Ћ;e�h�43L����RRi����e˛W_azx�歐�b6���>��$��ee��Y�a�z�k�����U%�ST��(}|F`j��4:��Rx�7��.级g.�E��s]o.]��cav���˻���]�kWw7nj��
�dG�G{��޽�^�A����^���Be�_y�.���\�zs�y��W�������n}��<�V���R��ݺG�7}�dg�%�oo��5,�\��;2�N���@w�d;Pseݍ#BѾ^J��f��O�S�ۮ~L��s����6��q��֥��KK��/��©�n�>��8ݺ��_?gQ[����d܂}�!��&ΰi���孥��1Ԅ�]�m�Q����K���0�,�p��d\��U�RL/�'��������SAI%�-�Q�2��Mjގ;���ó��!���S�%#He۰I��M�䔷��d%��ŭ���/.y�eG_Ep���r�'W�D��5:l�a�(�;2p���r\Ѻ�R�y�y��ؔ��!�+�0;��~�p(�UB\���0�*Ml�!ڼ2��Ml.�p6�F�J	l[��T�t�(F3�JaԴ��U?�N)d�\�/�X|v�z�m+��;H���ykH��S�f���>�>(�\�R�z���R��(��E�!L�a��x�8J�H��fRIA؋��3�45�YK�:- C��J�O��,�JI��*����d����``j�dB�jC���MO��gT��Y��JN�q�6[SϮ�\ԀCᆥ3[��>OAx�@�ĥxwL}+�TW�����8�>��T��KA��1JiVj�`�U0[kD���*2�J�zF�W�&����}Qnd�t#�@�u��2����<n�8<L�	��/��}v�����''��GW~��臻���+�����=<����qs��/N��<��������/�|���V�gO>��o<}|�;l^޶/}���;O.n�6��W�<�vw�����������8 �㱺sԯH��������J�.s�V`���9��l`|�8�OZ!���V����p��8m��i�k8�I�M�NƋɫ�z(���"0څ��K�ך�B ����˦�,;Z��������H�F�;UA�s�?;�x[Cd��}���-.w��;B$�̫��;��PR�+M�\"�c��g)[�^��p�(5����b5�4˥�<�X�ΰ,MPO.K�M*>MM�z`; ��y���7�&��XHj�,\UU\C��
g@��(^6��(}���U��u�	��Bn��I'>ے6��T�C�X4�3�
�1�-�fJg�m�t��ݯiR��/�����6�j(�^��9�y!MMaPc eiQ�t���~��fh�ZKQ%@���� �1��\�D/c. �,Av[j��9p%"]��0�g�X��:rʑ+���0�^ ��e��� �}mM�̦������Ǉ'��ك���ލ�����߾y����ͥO��^�~�9{����������G�>M��>�qC��v�.䱻+n��<��������lw����<J�!��۝�˳�W�7_������������ٳGG'���<���7.�?�ykp�S�������g������:�{�C~��������'~VIk��7�`C��)k�Zkne��X�s�=�2Fny�)c
g�E���lGP�¥n�#3����`j\��@����������\@��# C��닥����9|��D�я,�j��j��l.RycU?	\V�n�̆O�U|�)|�YƜcRy�� SFc�(^����15y�
K
���&���ī�0}���PC֚`�樗������N0�B}���?8�D�O�wt�3��!Ԑ+�:�2x���ND=HGk"	�K��nH
�kB�sQ��9��G��̋F_?��!�>~UA�d�:��Wфӄ����$ʸ_0�>��?�rUd
zQf�E��_��^�B��~��I
�`H�2��\�f/0<C �VҼ�J3A��TҐ1SL�4��ȭF�G#���a+�P��M��Z�\撷)�+2o�ؼ�B�;Z/��'�OdF%5�1Hi
^;��0�sXTR�5.=f
� #~v5���M���3���E�͟�������H�����@`}����c�yE��a�	i1+C �YpaF�}�(}|�j6ę .oSNp�0 � �W����QcW�Dl�&�K/D�|�g��T�\��0��b����)�4��&*�� �ƴ���3'��]ZE��/���e���U�,�X�p�V�>�M��G}��Y'�&o�\_3o)�D�����R�g��f���.i�l�d&8E�h��fQq��P*0D?	se"Lc"ٳ�pCm��0�K���p|�R���&D��!��N������/��!��df�p�6J�"�f���J��CZɩɨa��E#¶5�\�j��h!8�G� D?��-C��pv�F0l��4o=���)�B$m���a7S��,b_��~��7���!�u�&)�D�*!@z�tZ�l��[.W6od"-;Cޒb6�B�
�r��S��EšS8pvu�!�Mfdh&��wR��#��x٥�N�e���o6�����MKoO=e���[�����d�MD�T=��z��XX�X�';���r��x�8�㻌�ٮV�w�nd��̣�ݕ��AX߭.�P�۽=v�ַ07��W?�-�_��������֊�﷝;�x0�rWR]nx�x��} ��J^����8��8�F��j�',���v\��)�Ks5�ϒyp���@=����������������4W��\�ξ/��݇>�;{�]ߺH�V���}��֮}f��=p;��q��ή�4�jm-5�m�m)6���&PTۑb�i�����U,�B��X�����ۥ�i*�կ~�k?l�OA?5y5��Y� ¨'(�>���XF�ΐ��Z���M�1���oq"{�P�dEY�q���O>�eM_Kp������!(��,�lH��#g؛G�aEB\���]RE*N�D�DЫ0��=.4��Ech�&C#%\����h�sAӗn���	ds6kQ@}|��Cǩ�d�2)"e!���
ck@�M�BK�uT��v���s)p(�t�9���}gu|�tx+Im��lÒ�!1i2��B�@��@��O?��g�D	��8��P�/
��b���!/�&�uз!��Zo���t3�@��zdCL=Cm	�Ȣ }۱�������,�Q.���k;�d��m
4�Ԗ���)O�/�Kl!����Ȕmt�e��!H4C� ������/]�wOG�_|�9~���{��o�����������-7�>�*��,+�T(��iEG��p-�$����I�4=��=���s?K[�{㇚�F�w�{��w�N?��������w��]�^o�o����݃�^^>>��󁝻��|���θ���9ؼ����O6W�~�vu��S��>�[g���Ã���G{O��;?�����������w/���!���ѳ��_�ݾ�򹤻���ˋ�����?(�O-�(�_n�j�oKs6�51�l+m,ʲ7sEA���Z�d��B� �f/���(Q;Y!��h�饈�%���h�y���q�X�W|�� ՠ�j����tR�׀\�����p���F�ݺ3��V�E1�v}K!6����o�8\��Wf}�G��u⫖�BU�E�u��������t���� ��T &���&�����7MH��1*[�R@V�����pD�9.6BF�p�l���@C�@%E`h�#HVC6d�e'�i�L�g�:��4Ѹ��B�B [�Yՙ���JdX�V�P��(B�����
�Y�����ld���hZ�C�N��kΛ���o<�����[��NT�@�!���E����H�Q8�1]	�c�V�8��qbj��B� c�˗�� ��%RoCH
�[����F�gC�2��F
ٰ����N��5╗&�>�N(�A��Ln��L�Ó�������/�/���Y�^�|�|�3��tﭶ_|�����ѳ�����o>���������~�c�U�/mz�xu��`��ؿ�v��O������{t����?{���}^���Γ�ӟ���������߼�ዿ��\y'���~�����W������>�󹏿: ���=r�ӓ�����2q��������2Zö���Z=x+����ٙ��m�|�d�`�������ph
gP&���\@�a������+)xQ��3Ď���N�B�PД��?�o�Դ9d�X���F�
K��F�z�ə���{��,h3��!�jh�Ӑ+�}c2#�MD���� ��Z�O[ZQ�3��U�,��gkx�+H &��0�f�+*)��(�8߾� �2���O7��Sk:�h�������6eF��8lH:��Ӂ�V�aT��DM'8B���ۧ��!�eך;���[���a��m�l ��\M��(��T
��dC�1[(_ck�!hl������0%e�U�x��R1��!e}���\���Ya����p?B��l���,
�#āLפ�Bޚ���O��x"V ��XDOY�ۊ�5^"v�&�+���J?B6G
 ��!��e�fL���`(���-��}�h5�m� ����2��9�YXF�)
ӰX��`LBI�-q�&PHvd��j
�㔷�W@��t�#���U�Ym��n��q�C̽����r��C��>ͩL���K�aeOy5LH��+R�P�t�Չ�TF+���t ��9)��V�z-�KǦ ��YL|`������El��g˫�9�����J��N��S���!�-�(8;A�6A!h�z���Qa\���54 #B!�=}=NI���d�� lMH��C�f�ɦ�U҈[��e������bE���;��^^���eW!o�a���hy+#���8����Q�hȀ��V
��̒p�z�fȶ�������j(>����Kmag=t����IѦ��[�z��#�G�KcO�8%"��Ǫ7��j��PSa�h�)���y�V#!z-�\7!�S�+F����KgWF65�a�L!b���ʛ�_�������<��"�#/�V�������+�I�
Ԁ�� ¥Q(�ǐ�����r���7�ƀ�9�K�Z��nX�l�)0�Jl�R0���U*Z�mT�g�����˒�4��[�7+_�3��2z��{�;�Һ�+���ͮ�Q��˩���V�7�^������|�����v���o����c����T�R�N��w����j�טּ����򬾝��Z���^��,�>����Ea_�\�%�!9�5��^��]M��2��?��V-��z6��y�M��uu���w[�Է޷�f仛�@����7�7{;Ǉ�Eߞ><����+�7;�Az}q5�#*�o�.G��ȶXV�ͽ���\��a��dLeyS�?�=��(
����mVC-��|���fq�N>S�<C{`wؐ�3�>�Ta�U�}56�&J#�7����yi�_HF�C�B�\*���Z�0~)L��A��
1�?��Ͼ�������Hs��C�)w�2�&���2>�z*@
���V�} �V���V���t���fJ��!�[,&e.R��88��b�)��T����Ί�	�H�(=��(�5���M%-���h�!��q �"���pU����f!�;��ez��\�����i�	�"|�
O��*��X�ZB��3J���Դ/�f%ҵ���q�r��L-�~��1q���pJA�۠�u�d��%B��#�ۿM��*B!Gdm*��Ip�&����65�I�b'w���Y��bHl:�!��l׀��(\�ʨ ���4��%%I]����t1��}7bL�ԧ�~j���o���m��L�{S=u�m]�(B#g/�b�դR�t�D3���N��wy��%�y�gh���#��!������ײ{3.�����;���t��^�|��{w��|�bw����ًoO�g�{�������._\_������������j;~k��������t{���/Ϯ�_����=}���ΕO�>:x���?�n����ǟ^^���
�s�{�w�*~�勿����û;~*�K�ۚ���a����K/�&��ʵY�\+c�@�^�VD�B ������k�B�-
�M�1	B��M��g��K�X�q��k�ƕ3���� 7S^4 �m_4�dm�O�f)�0K���y��;8�릗_��裏���?93: �{�@7�1;l؝C�l#�Y���8���[�HIE�K�<ۡkh"��d�)=&ʥ�iK�qZm�l�˥��(�j��i�nڵ�6_�c�-r�ȧFӌZ�z�&V/V/���)� ����Bp��'��V��\8Y4��8�`kh4��8l~C�t)��Z�6��ռ�Ya�^��rY���㮉�'���N�$y���@zQ�ڨ��˨�`��o��5��O�Sw��`8�զ��z���V����A�g���t��ٌ�������!��B�Ňt>I�!l+o
b�����2l�P�}F/ o�@HC��R�ij\��/u�@��j�M���U5�:���8vo�N��rёz����3��+�����G������9>x�>:X���<��������T���~�����OM�����bu{��؈{7���������������j�3/�y��<7��?|��oe���o�����\}�ݫcw:/_^}��7��轇��n^_~�{���������/������n��ݬW�ʰ_��,��1Y+ �P    IDATj=-~\��I5Ģa�ucD�[���m�e}����3�����F�7D�Θ����㐔QH&!�6��U;�*�j1�|�v	��{��kB�!��5��1�~��[��,zo��Y�t��Y�GHJ
������5�!��95�l���p�����ZØ��k
B�%K.C|�����\�L8��*�o{lEʕx�Qas��$�p��9��."�)%���C'U�����6)4xs�g`�K�ܤ*/����h�9	�k���6iB 8Zkȥ��6���q���OgJ	d�,��%yui�ʫ/)�w6jh��a� ٰJ�L�pxj3{QB�J�Y��������L'�tB(SЫAk�y)B� �Ph3�:+z��2�����˅�J&���y5���Q\h�NW�4%%;iC�m͢*#�NC����U9�n̥���0
]64>G_U�
cDH��o��"0��s������.Ӝ��Hgr�%�o�WUR}�!"P��,8��t*�W�-PxY�m�I(V����75�E�GT��9G6B=n^��r��)#[�6���f�����f�� �o=)"����b�y�����E������( ��A���ؘ@
�P�~NM^|���J7c'i:٘�Z�x����b:W?[S����*��)���V6;��F߰X��ᢣ7Ԫ!���ā���UWˋ��>�zp��%E���T��R5�i�l8e!z�Draj�826L���:G��s�/J:x�4U�5��[\`x�U�ǁ�2��,\�a}����ق�
3H1��+ _Fj1����7,{��)N��ʢ�$�×FWҼVI6�ܗl�y,����Ґ�
���p�\�IL��x+�P��j���2M�C$�7PR}"m��%��G��Ԕ��g󥉦�K'c�m� ���F@�.����+�E�Ťo(j@�{����ӄ���U&�ƫ�?uJ�T���
��[9W��4����K->M��T46����*�f�+-���-wo<s�WM|��n������/������G˝��e����]{ڐ'�^�_�������û}?��J�7�����k�oubl����K�7=��1��{����\?�v�e�s���QKO���)�ֳ�|�t�Z�΍oUڏ<U����g8=�v��t����|Ut�~�����]�u����ǧOx}�EΓw�W�C_3=�]����������������������׾��}+�U����l�w-�ˋ��2�r+~,�h���E!Ă��Q�J�����1��k�ȶ�
O���kz
��c���sA4�8���Dͪ��/��+ꅄ ���z.�
ȋ������a8!k#�-y2��܅�Ҝj�	�%�5t�O�{f��_|��~�K�.��gL��Bd֯�2Z���!&�u�ttC�e
Gs'��F����t��f%�6����4h���oa�fQR}jbU%�a^RRb���ec�!õЪ5q�h�B����$B��!�a�pr���p:�`��-+�BL���z;AC�@h��߆�l���Q�M_
�����#Gj8�Pg���Y'9�)R
j՟l�B&�&;o�c�A`h\��504�/;��F�Bpس�pW9o���+]kX��Ʊ��=_�O~�_˱������u�n#�5v����fT%���}�n�V�R���٬� ��(PH�QN
(Q��!�>5� ����������阋^��qW��:�h�E7<���aY���B�r P��1UP��m	$�f��ǉ{��@ηRlI��>�W��]�����[�y����eI3�z��47Wׯ_|{{������ٓ����>�����ӓ���G�}�Y	< �������������{�����y��l����o�W��~*�S)����λO$]���qw���nή�_�|x|t�����������w�y���º�<�ye�#��cG��lML�ěr�dqZ@=>h�2��f\@��V5/So�-#��("������va �q0�����?��H?i1��H��v��9�4�seѦ`Ƭ'oC��4��rT8 x-�}���R����}q�/E;b�%�ՓAMz+#�N�`p$������)����A�E�씁EI*�&g6С%�a���������Eͳ6�V�!��*C�����T
�ȷ��	.�7gpQ�� �6�-�(���ژq��e�o�z�b!1sQвI�1#�S0�ع�v�@QZk�U�M%�:�Ugw�E�-VI���2����{�6e���w�m���*O�N���`kj�rGӃg��_ڸU.D���2_�l4���I��畷Q�5�&0M:�mD$���hʹ(
�$��Ф6ԇ���˖��M!2���	ۅ�x�ı�I�{7�)4ǲs�k�X�Jp�e45^d����{5�?���&�y΃��wm~��r����\_|��4������������Ͽ��<���xd��aK9��L�����UL�����c�z~����vowW�_~��w��~p�>������W\y|��շ�����~x�g�����;ׯ��W_m^}���/?�⛋͕Ϣnw��㓤���2����Z�0�V�ni�۲�Ma8s#��z|+�z&"���a�ϡ�S+�A.��&����8A|����B��,Q�J"��XmeH�4�\�re���� �Qc㔷2F��P���5��
�E��\v���\�ҵ�����C6�LZx�d�S?J�0B���X^QDj�G^�&�@��ɲ��L"�9��!l}j��t	)Q^.�|�)�a�B���U�+#�f11q4�����C�ͅf��A�K�ͥa��ѥ���5,vzq!�-�Tf�&��\��zK��ގå���E�U�Ϊ2�V�0\��/ѣ�������ֳiʢg�w�4L�(56���ˮ	Rf��p�xDӗ�09p��]Q1�0 �������z�) s��t!S��)������%��VO^Cx3��Q�2��񋢙���H�;�Xm)�5���'�4L�t����MGß�gW!���5�|�^v�r�p�,��y1q�)5���� ��3��. r���nȎ_��z�������ń��@����~ʖ�8WYؘ���V�q�J�"+?�}}�aY��"�]�#+J��=MI�)��`���p�V�'Tg"z��(��6�z�W���4|�e1�BC�@��9噋!�I���G�D4�T��G��h�`��iX��@QŎ9�[��g�8�N�P_6)���΀kpeW-���RL}��D�\�	��2�,Q����f��,��$v�fa��׀Vvæ\�\���ᅰ5���jXR�fX���v�e�*o�4c
g�-�^�o7f@��J0���3e���TC��P=�lr�r���'�̘s1��/��ʅLA��Q}��;���^q�s���h/-�D�ܷs����-�>ي��H65o@����R�$��84�#����hX �}U%ŖΨq��>��հ��Iq��!���	V�Y0(L�AY����qd!��*QR��;�3��Sybk�\��Z^R�l�D"���b2y�|�ciݖ�+-���r�T�մ��,??�"����B��\���д���;��ؑeL`X+�9W��w���9!���g`�E{���m�X�����޾�!�#���x�79�L�]Q�mߣ��+5�޺H����&��| <@ÿ�#�#�ۍכ�迻!�B�x�����w����?:==v��u\����j�Z���Mn{;>�=�[o��/v�[����";u�6�n���\_�\�o�wZ=�h��>��e��c�UL�W"�p������
���������a�;�D�X@ ���撋�̞!�\��k�Rhcü=��eo�$��>��PO�1��ۣ�Wvd��p�E�0C�V��b!l�55�^�JZ�tf�����7���z�-�E�8�T�a��'��6� �̅��CвC���v�k2�B�m���>}�mߖ�A���&���9G6o���̷�4DVL���Z(��m}6e.�ܐ���å����/fC��p��3­�9�-�M��j��'���ʲ]�r~&�������ժ�A��ݲC�ʨ�)֐���Ɔ3�Z��9��rv�EU$P�/�X�ֶ�i��"(��$=�X�^.L��&Z�h�p΂�l������n��֢�������Ծ &���Y�z�1SӤ����V���	�f������Ԑ)�S=B��V�A��yU|� ȐE�1T�u�9����7#�2:ݚOܤ��V--{�x�4�欩��iX�s�ie�
Gc���4�M��mJd��ݣ½6�K��x�V4(�cE�s��@&.��z�틿߼������o�?����''�<������\
�}�����[^w���>z�g���=_�9�x���/�޽ypr���c�t3zqt쫠㹠����_|r�9����-ғ�}h�sBWce���G%�ON�����j!��r�9�L��hsFV�˲��b٭*q!���p�@vd}8�E(Q��y�q ���2s1�����l��!\����3�3].|M�������pG:���M"ǀ�X"C�i�E�:���O>��o�rZ|	�!|C�b�Z�hF��<�V���Y���$oG
)�]���ͩA��/�G;�X�)�>>[k��� ���m
�TR�	M�\���m��a�2v�j����&�p��r�1�N�� �Ĺ��ԒB :gY��m\��Fq�D������H�jd��:�-�Mc;�Ha:��.mk:@QI����5[ж�����MMC���
G�k@vj�s��ц`3�U�"hl5,zW���[FC!�M�0D��f,PN�
UIIգ��5��V��,��EN����5��>����U��.��B 㗈˰	̨GЈ��@n�!dk��϶y�W��O<r�̯g<z������~�������g:�?���}��W_��[�+�~�h�k���{�+��99<8�'��T�{����z��������Ǿ�z���o���u.oΎ�O���/>�胇��<�������w>�����������ŗ�~��ŋ~��̋�������G�|t�%[`|���Ol��S�49���EzHKdz�`۱m&F����n�E��Z|3셻e�EA �
`s��4�ES}�t�8zQ13�B�kp �\!l}�i3 �t����ӜFm���_F8p&�F��55 ��%5=�-wLjj2f�֪S`ƜiR8m)C�t�b��:�h�z��Dp�g&��T�4Q���@�\��Y�@�qڑ���E�T��y�땔w�h�J����224���2D����B�r��ҧ#{�%��i h��zd�t�sH�6��B��B��f(jJ��9�[^��椤FЦf4Öe8B�˧�����1�C
����ƾ�>^�p}+����+9N�*�P?�����ψ�~��Gn
їz�!��GH�RϨ�KHY��rL���aQ�� ��i��� )^���AK�϶�J���a�4�l���:�El���3]4%UCx �V�	�|aG.�PkˆH�H65v�|n�D���5C�b���J�nܰy�Ȣ�Mǐ����_��1�q"+/�U��\��+�K�J<p� �(K�&��#&��p�!��7,�!Q�2k��8���4�FŇS&���\��Iqip|�#"`Y�l���Zy�Շ�����VC&Պ��E����b�CC�F|CMMT����&��5�fZ1�B�bj�Bac�Y+��5�\���)׷;h�� �5,r��I�!Ԥ�����3)CS���7�O��QV���^T:1��T�(:�B�������Ŋ� 5v��D�g$��H���P�Y 
�[��	�g��t�Z����Df�������y��T��b�����ͅK�h� �&U%b�ZCޔ��S�K���
D�_@�8��+�4C((����� ��@��w�.�xώf���0�6D������jB�n0AH�&�ڙ�+���&ҩ��q��bd!�H�4�S*M�C}��4��d�+o�%�H,
�P��%���J���պ-�c.6ڈ?
�����y����\o]���I���׮/*��=s)�-K?���Ju��軔�s;�;WX�Xܧ&��HLm���U��r���G�?+�ݖ����&|���,Kak9��E������ՊWeԗ7��y~�V4[��{+��y�W�Ƭ�lFn�p��yl�v����]����N�r��qe\�];[o�Ǐ���Ν����1�˷U�X�R{8���+��,;�8X���揍1�eOX���;���-H�i�jm8����!{�޺�@{���B��aC'�V��ζ�)	�nY��2�s!k	2&��>3cr���W'2�Ky�e��;�0��Lg�fj��6�JD".�6>���g�Κ$9�,χGx�H� �5@��Ev�Դ��矇y�y��z(aq�BH �X�#���T��G�P�z��^U3��,���N�qw��Q������u��o�q��J�X���;���u�+��MæL����} ����g@�J�]=���uI��b����͂!���) C0M�aX��d1e�ҋ-dzK'VR��ɋ�IQ���h�B 8l��is����Ԕ����n+r�F�ת'�XF�H��Ojzc�>��5Df�C�����'Is��O*�(ţ�Z奀ițK�fշbhB�Ŷ�4a#���kK7����]���o~�_��c,ݲi�	J�����:5�bگ�'^����)�!ܐ��)+�]d�{��@�Z��r�mj𹁄�J��P�^��2�A�zԯQs����ʷ��>��1n�fO���g�~����}팳�NXf��4&�֪G���udkJT�m�G�0��B�����W"<C�k��b�xoߎ���h��F맟ɝ��߫�j�_	m=���ų�����w���y��_�>z��$OiX������z���������m�/����.��ǟ_<~wt�:�3x�У�/�קo}��������;�?�ޜ?{�]o=��+���n���y,��,����Z�xO]�������2�1�6�\@�lq����ޚ�zE2�0mFCQSb(
�fȀk��̛Z=W䆓 /�	�qAڔ�H_#�����,A�������a�$�d�
Ȩ*�U(����6zk��0vH�׻�Ү�A R �y5�#؇=��K�����嘻c�P�C�Q��$m9\��6�&�{Q�^$C.vQ4լ�V�y��'΅̆+����]�������	�5�'�B�
@P5C
�f��K�ʁ�A������I��2�5T����oz!�����Պ��d�#�N)2ؖŋ���^�_�b�;�i
�٫�S���Q�����p>)���LA_v6#��]/�aK��%u��f,�B���D��'� ����S��Ȕ�ɥ%�ņ/�(Ȱ�v +���[%��������
|{�b�u�٦z�/��YXF��Bz���g�H�P�RyM�����{��pd�@���S�WGi~���0K��������˫�_�����du~���W��7G��:�;v�~}zx~�������G������˛�����*�-W�ocG��{Ǘ�^�_�<��n|�zy����v�CO��׿x���o��������>8>�?�x}���������������Փ��k;.�g�G�{��2���4+i��F�<VҶ04�v��lXHK4W2��@v^L6�!�y���h��Al�S DIz�:z�q"��C2�1gU�z��5iV�Px��i3�#gWr��56�+���B��6ԗ����sA���Ȧ)p�e1�Er�%{��8�ʈ@�fI�+��4�&U��MR���B�\�����=ހ(�%��$@���@�%��q���\����:��1�r5\X�F���JA��z^Q\�Ӏ�d,q?\m�\��
7,�w��+W�RaI��RaQ����2fͦ�)D �9������Z.�]R���,�&_8ܞ�(�-�VC�,����2B�Ț(yklqq�    IDAT�\�Î����'8���ҙ^�@�lF:�����*�hz�e4^��'�oj3#d�J!��a����q�es�Yg"�y�Vm�ElLA�QUq�E�=p�O�w�1�Z�5,�ް�rͨ�U=�VU\s�55�/MK��V���Ef�8����JA�Q"�hވ#�?3�0S���fX��1mD^���j���xkl8�	�?P�P�)�~:� a�8Ԫ?Pߑ(Pc���]]�a'�7)�9�?���
b���$�k�2���dI*eLxU���!;r}��|�'f.#�f>��£����D�D�(h���-ض��\M���b�5�u�j�xI�F���Ϟ�,/5p����z��Xs�%��nl�`�6�)��3��X��]x��7�R �ְ�DK�=�A�ܝ���(6���!~�fR=bґw	7w=Wn#�58rƒp,u:���K�͋/�Pm���L|�
���3v���D���gL�a�*�a�^
����]�\s��ݦ�\�j3�0[Og6�y�Md"h��k"��s����[�o�����1٤"O>#�}���,�K����;��">�Y5��t�>�Ɓ�,���@F�l_�����If+ MRb'Ӑ텱h�@C��ӶJBFX����fXy���6�5���$�4n��ތ{7}ޱx��:������N�����B��rT��6�eJ�������9RO�����]1Wݣ�}�v)p\�tr�S�$;=����ĳb#{�'Ǉ���Ooݦ���<�G=[v{��JG���_ [��_�.d\�K�̤�ٳ��p^Ng-��vs���͚���7;o�Bj�w�{Gk�����ʄ/�����~e�����_<����2���_>$��߼Y6�<�]=w�,/�0���������4Ø����0��ڎ>�Dd�pjԐ-V������R������`�oo/�-�����!1�\�iϼ!��$C6�^K!��b&(������tvӄ��NR9�gv�h���p�R0�O)F��0L� �wyyi:�Kկ_d�[v*&P �CO�U��`.����%�K��5!��rR
�����Ԧ�o:�ʖ.�j�(�#�D.W�1ӁW����"!K
�ÛByq���^�@Q.{�� �������%��pf픻3��֭��
���U
�L4ov�݌3uj1�I��͘��t�2A��� l�z6٪��@,E���p̑˼��a�1R�)�P����OV^��}��<��|.��E�iCy������;m^"8/�Ԛ��� 3BE�.�i�{!vl7�!�$�hz�M)NgfQ2:�f�7�v<Qh\�3;�5���[����\ Ms�4��u1��R�b��`�^z^�&���9���Y�=�ݥKjv��/.Y6ވ���M�]�Q�#p���ni�ypp����=;=rAss{u�]=|�������۽�W��������z��w�_]�����c����|����
�g�=���e���{�ף����?9|�}O�߿�� x�P�����x��w//] �w�q7�x#t/�Y^Lo�5�k�͕1/Fh��C�2�#Ѭ�c�(Dxg,[�p�-,�S"�'2m�h�tp������W����(cj6Y���C��D2����R�4�bH����N���8��vT^K��KS������7�Feo�?�Ya!vQU�5I!����:P�:�9Zh~���@#��F�� �L:h�NRhz=�Z�� ��8��P,��0}�xW ͚DRk�����ovB0�P@���&�GGjp6L�A�)��ڤ/;�������!����?��?J�jZj䝂�:{���fy�{au9Ӗ���7L��D�-���hj��foqþ���g���(�Y����Q�Xٹ�%�
�"�f^L"��#e=�3���B��#�T�ح��H�4:����(�@ӷl��u@0�2���OƦ��;XV�"��?����)�� � 6���R�]��"T-p�z��*iȺQ�Pz���~�J�כ;�ru���G�ח/��zy���������/._<�8{�؟�����zN�z�����T��Q3����٫gs�Q8���non�0��Ʒ����O��={��w�.����˛���=98y�����\*}����5����C�}s3}�W+�_�H@�o[0�����MY=�܊�CLܖ5\�Pƫ�ՃXp�<lZ�r+o�Pb3���5\�F�^�y\�
c���餆#h������w3�%�Q��E
��5�t�W�" ��S \_����ƅ���8�����hf�L9���Q�e�V^�f�i��1���X� ����ȹ	���ռ��t�C�6S4�V���~��J����	�(>� [�WoGTv:��0�^%�B2J�UK6���K����LQp4.x ~H��Y�Ag�"0�ɯ΢��֒���p��"v>""N��@�%P���Kd(��i��²i��a�*)�]o�N�\yM�%d$��&����/�8c���b5��i�A���ҧ���pS3������e7�^�X"}(o=��Ry��'��[���A��%�J�q�f ��A�6�,�,4!�1��'�Z��Ȯ�@�v���˫�o�W�AHE��%v�E3�).�:G�7s���e?/�ɖN^e�<)���@����QJ���.){.�L
��љ5���=K��H�$���U�š��������$D�,o+ � �NF�Z.���/\_`��7�e0� k%��$���������j����AЗ!ؖ"�@�R�^Rx�)̨4�AW�٧)��J�{�!��2��U�Y���	��l���x�M2��F�Q�y'n(�� �h�0Kͨ$8�ު���8I$q�X+$A!�ē�WICe��@Ƥ3�l�d�%J><�2�d���a�{3-����B&� ��S�%o����,�t��%���K�&�>�n_:.�b�4��5
z�fm(���@-&�k�����[�^'y�X��c���flޑ��,F�eʕ��NC=fY��q�Z����g@*�So%-M�q�Z���_s|�E���I������$�R�������䅓��z�� [���NA �e�Iא�l޹�E��L�2(�X�)���[%�!D�sȘeĴ`��A��c�|�6Zn�t����%�?�u>��&f<�a����{��j9��jWq����8��w	pܐ�+�2��͸��P�j�����cQ��o6�כ;��5���$tl�Qز]�d�eqI��N���f�-��#��u��*z�߲U���|Iw���嫋WW��[��bㄳi��X�4g����}�l�9�`zt���������+�7������z���0�}fy�.�
C��8n��?z8��7���e�~���V�{Z���*d�8\2r����Np�2���"��h����kuj�8b��fO>9��풁Z��z�DB&����(�6���LT����v��9F̝���O�5�8�2R@ӸP\b���M��/ۖR�(�C�+	PTxQ�%-�D�R�&�m�Ԅ� 1���H��E�)����*)�thl�&�kY��̀�h
%�=�V��R^�Ʒ!^UE�_%���Bx3"��Ժ&^v�&sM�E׺�B�\K#f� \�KR��W!>W� ϕ7�pH`��Ӭ�^Fᥰ�{��&h�#n�]u���)A�Og��	��VFLnhC[�_���~����s�i�-E��pBrѡ_�s^��\h��
�k�Q ��g?s��t���?���'��MAx��T.����^��1��q*�@T!���Ү|�i��,��
��O~��%�����0��
lvG���*9 [*�j�շ�l`���i�)�7�����Ḑ�=�B�;�0�hn�$����ݟ��B��ۓó���g������cw�����f��g���[�g�ަW�U^^�z��_�<<~�ݟ�z�[��#���x��@����9-}�;ݘy�=S��~�s��������^z���W/.7�wǧ{~���1���C����?���sz��k�lt�f��~.�!�R�w�����m��K`;:;��f�m��R@��f8�X��7��p��y�EA��Z
�4RE�� �K�Ԅh!�i��!vS0�\.6�1�Ǚ
�vRq�܋��6�M6�	�z�>k.{渥.�&�#}��]�	q��^�ͭ&[߁Sal���
�@����_�R.-W���X�5!�(4_Rb�S35L-��hlR��2��ʅ\T��#k�dL6���T3��H D� jR끘���4��2~�LĆ��WC�d_�*� D� 0��0��c=�|yIU�j1}!���(̊)[��>�^*g�%_���{:v����"��D��B%D.��P:�PH5��8�@�z��7Z��L�����p�8E���R��#��!E�qM[lI�KĈV��[�cG������X��|�hjB���(s�W$��E֧:R�1�ƨHW�(0���ي�el�U����.��)83\/���~s����]����Ml{�껛w~��C?��b|:<�J������v���?z���b{����m_Į_]z�::<�^cJ'~v�p���/^=r���O����؂����n�t���~��w���k^�<���o���ѻ�m.|���������d����s���f|�l��Q���D���C ��L�M?�޲[g�)PK�f�ق��XM:d�z6�����EX��T+p��!�EH\/VO�F�w�Eq#LcV)�z�G6�%���X(cL}��K�����X��)�B��!c+-�0Yd��Y
>��2���f���Ԋ�7,���<�4�VZs�� ���-)5Q��B��Ȁ�O����`�a@�ְ(iOF�)D���f��N��-Rq�&\lv�����Ւe�-0&p6��Y2��������Q���	A����"��� 
,)�a� �F80C"�V"8�­#f��1�∝Qp�XOMv-�n�yE���,�
�*dk�����N_�f��-K�f# �Gq��5�kV	2\�ɀ1��kp=�\�h���[�93�*�(��	x�QR�n�WI���t��30��p̊�T�" �A�8\*��E�8;eH�@Rȳ��Բ�Z=C��eg��
a�&���w���#v�i�U��К4͉5^
�rgTH5X��z!��B}tj�U�=�M�+V
ޢ�)��z�z�{.����7���!85sRФ�#��
D�Q8�!��d�q"}C�z�pF-� �7#�J�J"Sk�8�MS�ף��Dch��5]D�-eLCR��ƀ�a�7[��
(��Z|�"�����@�1�4�l��Ym�\�A��H���U���Q��DA���8mWsߝ`Q,x�c�,$�
d��b���y_�IV��\�� 7�dAS������c8k���U
#fj� ���2����h��a�y�@�
��G���Md���#.�@�V=�gTCh��h�1ԥ�,
��H!j��5^MI�ᭃ��ԙNU�g������1�C�D�r�{���Y�f�#�jR �)��WQ�o�zQ������i�I5qje���+��__���@��:ͲT[Rz4�3���(v��J%��#�����Ƌ���ʆ�S�i(�
+�@�+�C��Ѭn(q�I�Z��;�O�����<�K����(�j�Ie�ev!���>Y�o�<��ˉ���1ϰ��6���.�K�\��}ٝ��]���f�����ս/�N��n�:";~�_��A�fgַ���B��s�+?}dWqEtt�����i����;:�����=�{y�Lm�+���Csm�#'��Tz��K����V=ޙ��C��ݸdI�E��s���m���ּǵJl��wY���h�_����o��M��_�E���&3w� )���V���0Ј;!R��}��'�E��lm����;�ޱ��,H:�s"h��m���MP�	I����C�t\;g���/~�������,�Ԧa�Kh�0�td)���q�W	����)�K�
.$e�(^M%��Jm;�؅�#	L�U�Z�c�iV�"��Ň�P_=��0k�!�VIM��	4ljDr�W��VR��C���.�,�5�*!����w���[�ag���J�4�S�p�)#���13,c�mX�Ը�Ȥ؁�enay�h��0)C�DU�i�=�N^�A�J�5��(�]
.Q�
8�s���[��b�Aڍ]�s�����t���fI�����f�D��JOG�D�J���>��c4�p��y'�{V��M��
��k��Q!;��2GMK!�bǠ��Ի�O>1_����?9�?���5���*c�*ݦA]V1
�S��0G�J̪�`��S��L^�j@߫���LcA[�2�����[�xD�v����~��~���'��I�<��d���]\��F�>\y�����/^n�O��������~o3��6���߲�[����v��^���^��_>�z��H�/_����n��ۋ�wwj:���'���D�OWX>6��+���sqA��/s|}���K��F���&жR�!­X�mO�5a���m���C0�A����~ [a�����/5 Bj��z���C��!CKS/$5 ��eW/�y'_8N��х ӱt�����g����w5�_��_<ڑ��ƮN�kh����*/�#Ы�,]����h���3���� Rm2L�ш(��*͐ ZjD\�1d�x鑱�.�yA�R���R@��K���e@*�@�\U  1��@d{>�������2�1��ҳ�:�*�\C��Z/��s�N��rT�
��SA,M.��R��������rf���Qm���Z�4mQ.�y���袵+�n+�Ex��B:�bEU�@�&�����L-q��=	ӛ���fPNʐ8;�t\q�sMٳ��!�sedO��TT=C�}��E�}�K����C	�B%�7L��O�����%�Ӱ� ͥp���0B�i"��i����:�h�%��#Q߻������ް���=:}0~P��ĳe��w����F�}q{�����o�l�f���}��#���Ə|��?�|wu}��-f7�[ò����g����|z����xu�9\������GG����P�������?���ϯ����V珞ޝ��������3�7�9nW~\s|���C���{�2�q8��o{��&bYRs����,�ٱ�:4������������4ʆ�=Gh4Q˒��\c 3��
�ߦ�D(]���~�"�lR�o��煈���s��l�K)i�Ѹ4Ìl�f��O����83��,v�	����-�kwH�D\1�b��$UI�VO޹P4C0��EuW�Ն4Yj�Wa͎^:��D"��@C����6��v9��5�8,�FS��V�zxE��༐vTx��3,0.��R)��IR+�=	ei��E���\S��?\xQi� S��4s�Y�]5R���S6��C8���%����uug�y�� �-oC��+U%�^".\l6#�Lݰ�/D=�lC�D"�\�Jo؆�	��[����>pN*M=���,���h���P�+P��2��!
�ɫo
Bx�lFQe�`^��-dr୤>)=5́�ƤC"�Ɔh� !lL���4���/
�5��An�h��z.�,Xx��q(��Q#���/�>�|q=[#��]
���1�j4K��k�&62��75��0�����LnX+��!W�
���+���f��zQ4!�+0���RD�S��hU15���S��~IyWj�aR��z�V�!����R�KW�\���%��l��?�d��Po8��U���,�l�r1v&����sV� �f}�� MV�JؚW!C�j˅�5��m�zm��{� >�w	��E��*>s�7o��b�S9Z+0+�~C��3�۾��-�
�IW�)o�8�RbBJ��)J�/Z;W:�r��OP\�D�j�6�I�YU����C���@��Y�Fߐ�d'y��xuN~"�%�7f�"���U��    IDAT�|���p!��l�-�yx�n�X���W*gr�ފߗ1Z��4K�Ӭ^..m։B��jcWI�lM���,��w7ټM���m�2:`ي��w��J!�!��1p4F��̥6`k�p�����W���Y��Hw�9K9n�tS�wR������˛�B��4��>gX�?�s�Ӯ���8�ꚥ?���#�k7?���q��ӵ?8��W3Z�/�t��w��}�	��9�������P��o�������v:�'�8B�/��6�1ǭ��6��ۚcA���F�ݞ�>�w�[_�U}�ʨ�p{����_��������k�o׫�[t���8dV�7'�c��]�t7�]`36�h$��m��5��y�1�����ٶ�؇��B�t�L�-kJ��O�!���"CF�߹C��q"�2��*/o^
��E����w]�@j� Ռ?���-N��?Y}�	6#g9���0�7:��em�m^�\:렯G������e!�L����.��)��!�@�.��U+6eUe��%�k��%n{EH�(E�j}���(Le�B
�O!A.!DT�f ؝�Ѭ?D��^o�]*65�4g��4|��ф��q-��줢u.�����+
��z
U�>oMT�9T�������G &C�D�HU60B�)"���x�����p^��q��}��5�]kb��I��Es��G��p�(C�M8]lm����HQ6q�qv	��.��m5����%�x��(�D�mP��R&%��Ɏ�F�H��%����m:�����������/����۞��֎n�D�븢+�]Yq�2��(ѐ=c�bo�\���8f��~�rٳ�Z<�޲�]���ٽ��iW�=�Go�����_����������������i�����%�ǥ_������9rc������#��m^��@ڃ��#7x~��7o�><����\�|��g��n�<��{�qK�f{t|t��{�O��~��'O�N8Y}p:�@�{�+��Z�`|i�ڊf��rY����8ȁlۢa�X!��1�������3�Q
���%�Dhs�k��V^��(W�$pr*��F!)�!��%7d���)h%*�(�����N� �;!D�2W
;�����'��}��綝�'�B�A����c�d� �^�r���`s�����H!�K��(��� &M��Z�`�Z1��lM�}��*ɼ�j��e�Q
�f�z�d��R0 C5���V$�p��LM��"W9�����hh"t�h�o{&nj5S�0�4���8�B`!����Q
^q��nk�J�_���e����rQ�6�����p��S������� I�?����K��:!m>!2�xq
dS�K$/��<5�l-)�l.B
g45����5x�����2��G��v�Dx3��j)���G����U=D(�K����3�������*qYX^���_�u�#�	�,�M:����v����p����&rxp����p}|~|�g�7�'�2r|�����_����_��'�o���������]�]]\#��N�-˾�<���i7��]�:\m/�<��7��7���ɡ˧�?�����������WϾ�÷���g��t������������o_={�w��}�jﶯd��,S��\�r����cXO�����]o),Z[�e�C4F��ty���_}���z��Q�	����,&p�������ѸBx��Y�4���eTd��Ϋo(�͊_=[�\zL
B��lF r��ٕ�å5d  �ڮ+�\#fi��2�a��]=�e��]�IM>#e��)m��奌)����2√�h5 ��8-,���d!���ƕ,�p���gG*�J�^���iVC
�
����U����G�5��ZL6ClLKĮ*4Ӕ"5\H�9켃�ih4�l�VT/��8�2�\�<�)�bT�!��z�4x���F��ҋ�PvC�L���pC-r|C�/M�\���P�, ;q4�V6АT�k1l�B"�Fd:�#�X�j�=�c&Ҳ��F��f���/#^I�������%B6���5	�8��v�p	aWvLR����Tk�e����%��(�3*�Jԉ#�g�T �a����q�20#�C_"�@�&
b��	ѲIi#~���A
PϮ�]�
�!�46rRR��z���%eL�YaLde�q&-�jH<ej8���%t�HA�[��٥��3W�Y*Pj�p�%
��x�)cFH��#��[��r٥Cƴz6��o�E��b�^ �V:���"��T�^����ܑqr�#M:���^��\3���rQ�t�yk�L�t�Ε8�1�"T�� MF�I?$�fȠ� ��r��R�	������d���OJ c�5��X��^K?eQ�Z|E�7��oX
���Df�K��'G�a�4:6:�j k�*�3��L��;�8�h&���q�%J<pڍ���f"-<��-u8�a�D8Z��
!q�
m�j7$��ѥq��Ń6�p��f�Ne�˛ fޔ!���|~h�
��e�	�1|�ė]x
B� �B��d�91��4ejh�-�X�r,�K�ՏI�ڒvЦ�ِ�Y^6�j��H�y��k@��t}��j}���j�
$��Z��4;�գ��ӳ���R�p㦓;?���2����pos��������n���/_�O<�����#W��6�<ţa7�q��k����S��:o릖Q�<��\�ݻkҷu��k�O7..��N���vh��N;<� Vح��C�A�/�ݭy��9����\�P����-�W:c���e�-�����/������Jr:w\2��Ӽ�����ԩ�gc�_����w�@����r�����9�qj�Vp�>c%[�V��ȹ�m���<��3��1�t&'&������I;�@��
�K�҄h�ymqj�X���3&�NŗH�f�\�GK�465|H��
�� a링 �M�a6�ɄTL=��2Bؖ��Ġ��j�]���A��Ւm�g�-�3`��,�MJ��J���ּ�9��hY�cW���)����4P#��W�X\��V)ʼ\�!JH��D����Z�*���A`ӁC�� =5.-q�����z/�գx�t2>�Jb#��	o5�R��@�ALMR|g5�8nr~�v�*qM��B�Q��P�h�^�⁋sx5v5�lXH"%�j�y!��40ټeD�
&�&V^��p�BLM+�D\�j�M��u�3�_12R�jm����)6��dkHR�z��l���()U¥Q({+����Tw�z�� +�`���4�EFp�@x�Z�2"tӢ9:4�`�����?���W�5Q��x���i��=$T�M�<E67i�CK�1�V��6�kȥa«L��wqg�G��G�u<*�o^����I��T���k7A��o.n�W'�~x�~���w�/^m^�?s���ήC�*�-8������x��[�N>8Y�{�}�����~��;�vj'X_�a�ԑws�����W���������'��=��Ӈ��o�ݯ_^?��\�2���?��Z쵿<�|�|����� Y��zw�4\f66�a�6&��Vɒ�NޱU����˖��62���ѐ��B$2Dck�4 ZdF3f8Nd:@�iP�����f]P���E���zM\_yhl��T6��vEF�8	2���~k��4��H� M�����*?4ޢ��d/���xq Ss=����Pj�t�Q���[�l^�	A�\����q�齐1�Wg ?@��dC��� �ˆ��uj�!�D����Ta���\�R (D��� ��^[q+Jo������24/^�z�����M.�������7+c��-��*A͊�y���D2,��`���|�a�D4Q�z�&�7����%�D`�h�)$7̮ǉк�Es2�8��g��>f�7�
?�bRC6�������,r����$BS$�+�� 6�\@���B�XY���05)lDF��OeK�,�	�90+;M�\�K��@�'�V������t��oF��������+�L��kϯ���~��?������'�~}�<c��^�.tw��������x������`�������o��6���S��du��?^?z��w޺����%�;�Ѿ����ܽ�����=��w�??����w�~{w�������ѾM�~h�o%V̡�C�����I��"�]!f��:�Z���M�/A�^��8�y1�C�e�X�?�z�Jg���<	��@R6M�)�3��8��p����l��B�D���bF��\�� d�E��$6��ώ6���)�b�@6��6�K�~ ���-`s��m��JJ
����I�N�QaȆP1�e��C6PC�e/����2/�0M�0٤fR�@}v���Dv�ht�r5 �4�XQ�\z��,	3}��g`��/�c�L3R,0��Q�H��E��"�,�\����ƥQk[�hN�xL������n�@�M�С��$�
�ʢ/0�rULv"�!-qØ�� ��+�����3ʅ��!0͖�����)V_�b.�ɢ��I�+)Zަ�Eհ�hC�پ�ch8��P�(x�U�/�D8k"��	�(HT�*)�+�k7����h�E#4TX���$�ɻ�˰p^4=/�&�&u����4Y�آpJd��mbXaB46������քT�����r!��ri�x!�TI��aI��l%� h\-HH�֬��kA8ՙ>Y�@5��a�E�'Ux�B�B:��z�曬@H��炈�'��a�^a\�e��5�i3x�
0_j��Ca7�V�>�#�@1��aE���"0:���\F}:8U>�B���X��ذ)�15�F_�wgs꒔`�bչ8_oe�*�+;�:�[�4_=AmWd�di^��0�^I��RaTm�N��,|"tqfa�֛���%����(5�]o���W�4!DS��n1%�L�!��\a�*L�����B�4J
l^[ۆ��1��X�S�F+�\j^���k�*]"1e���:S��9B���r� �8_��/�^�=�kO�b굖eNA�Oߚ7�kE�I���h�!�c������-�a�j�5�k���^���U��U���.{��9���pL�����>�"55x�*�5/;���1�;>?0����	�B�:@j�Z=�B�����^y($R?EW �;����ӥD_=y]t]���W[���ڢ�1VH~��؏}y,�s���ܿ>=�x%=��u{wg�<Z���<ܮ�=�b{wG��٩{E<��c��ϯ��]��Ĕ�gR'���}`�9��Ӗ��^�v���qw�g$y���ݛ��������=��n�I�l�*{�qz�g'i�cl��c7sz��������KVG�B	���� ���{i�Q��ˣ+��=�\��ܯ]�u�ŵ��r����OO
t�����ϗ2;�9��7�
�l���ca[g�f#f���8��va赶8qk5Ex� N��������a����g���esW�h���ah8��o��JRp��G/
�Mj�����d��7& �Xv�@�����"$�W�\zgS�t��^��,;�8�IYXC^;
e�8�HYU��-K�f.
�ܠ�+Ӊ,!lR�,6�MË�x^��z��8z�d���ש�&��\L�,�B4�C���H���ҧܤ�cGF����D̗,})����[=��d4�E�#W �\Ų��	*Lk��^�y�#�E*��E�=�]�_?AL5��[�t��Z\�ņ �Z��pU'C��	ZKaF�fW� �ۼ,oQ�bd��M�eA,Qۗ�Y1켆�YƼe��T���cB��ڲ�7;
U�Zoj�8 ��\�pFו�f��� ה*��`�h�n��d���(���5�O>��%wk�� )�����}͟�������`���"U$-��Ui�
2�9%6C��i [x
ddݓ���#�������m{}1���u�k�x��hۻ�g��z������9ݬ���_}|����O�yb���U����c{x�[o��~���������۫�����������G�>:��gO�_�'��������;::vn}�:��|���}}�Y��;8:s)t��xC�]�b�m��9�e�uKGo5�JZr�hq�f1�Vn��ml6N�6��tLb��q|:��n����g��9�|.����c�S+5|���G���P�x�=a�U�#xY�B¹𵊷t"�g=cx����c½�~���y�� CGԸ¿^�=��Ý�7,QY��W$^;�>�U]6��[)�\�OC�4!����ER��e8�}�R!�\1\pS�ٜ,к���\Kߋ�)��"���*���@�a�!���+�����(@O_O�Jz��	���֓����N/�@4�F:+앫z,�{d]�n��V��d�Q��1	z��I���_���)\�DT���p�]�����Ry4�Ʉ������rajht q�����b��I����Z����X.5��.��?Mߚ���򩎠���f��
d��R��#�om���Wj:يQg�����:�ctT���>�Z`���°�w��?߻>8]]^o�T�ŋ�G{oy<�_p�wxw{����]<�~{w������7O���G+o��^�{E��w���%t��<:8�R~%d����ŋ�~�nΕw_�l4�������w?zxr��|���/����_{6���sz<������s?�����w�������_\m.�FǞX)[p�6�9�i�sC�Lٳ����՛����H���.m�BD�����4E	�$�eIm�)�� l��Im���\�A�f}F�
\T_��g#$2���Éh�\!��'��^��O�3k����!M<N�q�z.�|M`��/�]��V`�Pz"6\F8`�z��&�=2�=��4F۽���p�`O+v	z�y�Ȁr5�M�f�"/�Wx;2B�g�4�b��!8z����d�Zތ8lQ�9}����R#���@:Z�R�E��a炴&�d�E�ъΥ�%>p�G�.L�Z����5g@�3k��@���p�&Pj� pC6#W���;&��ShA!��$"p�04B����N(v�W-CS_��-M�2���;w`!!��Rak�p�eW�ny1ŢUU�q��DJg�,�L7�i���������p}�d$;CD��kX^%1�����(pw�`"����F�ײ񛋐�O\=��	BD����)�//q��!y�×��kHA�^��p�ͥ�.�Aք�h��JĞ#0.��؋�E���1��" �n�1g����t��7G�[�h��E*�4��it���2��J*
h��x`�%k�2ԦZ[JT���2Єhd)@�@rM��'�A'�E���.��rʥ.�B;�6�?SW��5�������]�,��f�q4x��1	J]��bV9�:�3�!C�ի�����S��5x�02�
��$��TO�5SY�R�B�|�XĆ�Ȓ��4��P����`.��A����������V
��@E2jS��g�A0Է���Ն���
`sէ����ԛ{���'�7~.:��J�#Ch�yM3�0�adW��Z�BfFPKSl.dv8CH%U62�6s-�?!�Y�)��I뫫�����d1��-��c�1��d��Bak�T�JJM��'Y8�!�K�;��Բ1ɪ�,f�n1�Z)��&댊��!��`t�J
��#��bI1�z6��z���3�C\Mh����8�۸�oe+쟺�c��'��n77�<^{�����Cqݝ�A�N��Nzzϑ���x�����'�S;�f�3�>�;��o��x���='�}c����˛[�+���5M�����Z���ޒWV��e){�������q�{ԭ�`��c�9����g>��>8�Z\uY�^c�Y���\Y]�_\^����;|�w�B��HW~�ƭ�n!:>�u��᳿w5~p�Y���[kom��בl�WS�M�����e��'�Ҙhsc����)P�o7�W8i����K�mj8!����:W��ԉ5Q�T�U���6�k��w�y��%    IDAT\*,P?���!~��Z��	B�s�2�Sxd.!M�yT'����p�5�z����/�zZ��I9F�I�0�d)��k��
8���*djlG+q|G%_m��Dc���#�6bk�u��գ%I�%��Ԡс�/&</��H%V��k E��ۚ�#hj��ʅ�G����h8��V6o}�=�҉�Hm�Y�
G闌z
%����rEo8�@^��ZQ
l"�CtiEUsx����а���7���l��k�hj�Z
E�eos�v�z�YeCF��NYo��z.��!7��K����+/AC"������\�:^�<tjݵ|�T��6SBҬ!����Ԉ��M3��qj?!ȫG�{�g\���o��ŷ�8�ɮ���u�?���qj�&)X�:WۡBT�l.��zM�p��-�7t�T� ����v���"#����6ށ�ݹ���r�*����g��?��w��o�?����������������W냷�/�^�ݼ���ך�]v�_�x�;;޿�y���/n�w��;4�փ��6� ���ڃ���th{w�ٻ9�·>}��{>nx(���`{�r��	惕���<�A{.hz[u܏�+��;����e�N�%6)�gh0�,�>�j�������%D?Vf�m9=DTe�)S� )|��57D�B��S..N�� V'�]�>0DoIo;VR�
g3���J��a^�a�,��9��t �t�4�����՟~�������\'�W���0��֑�+5�(�ؼl���4�d� ��o��VȔ��^e�X���pB�B��:elǘoQ^5RpI�F�C�r����Dj�q��R�F��MeQ@R��e�� A�S6"-ed�Yx���F?M�D��#h�h�a����[�C�z���=_�U��(�)�+��^�d��Q�9:p\%���~��'�xY�Hv�8���W�����4��@�75�Å28�߼��@0lA�lQHʉ�$&Wx4C!I�G�mA�����7x7-�߹X�bGB+�65kҲKצL�8D_�@Î�V.j@:V����@��(SUl�3�";��.kE�!#A3f��[al&����,��?�G���+�w����N�}���~�����������>����ի��������<:��?}v�d{�Ҿp�e<��_dn�9ϝ�=/{��������ٹ=�װ���7�ӓ��g�?��O��}?{r��xz�������o^�x��������n�q���[;`n��y����b�˙��j��2M�֡-���f�V�e��'*�k��M��p�+yq �=���²!���Dfh*�	a����&<W���|C|�B��n�f!C�j�K�z�Z:�)b��P��z`}��%���OaN3��"d�@�}Y_��L"\Z�e��Sc#�E��r��V����mk�����ϕ&^U��ό\B�-p2E��"o`�^`H����R�3�XL�tx��BR�p�1�B�"+A�;�C ~�
���34|j\��l`������ !p���ꓪ�b��2 Z�1h���M�V�-�b70}d���\��Cn�b��1C�g1���2��FnX�V؝Ev��hZ)�&��`m�Z��S3kdSÇ�ى7�fWސl=�#��h�2�1��ߧ��Jm����p:�Q�Y'#���0/�dR�����^�>�$[���Q-{z�A��iIqE�:8U��«ǰ6�yC�q�3!)�ة��da��!�9l��.��>fYؚ�p���5/xH:�Z N�-������Os${Ӕ�|��͘��!�Z�����rH!�U)$�>/)�L��f��P"������oy���|�5��>o�(�w�Z�*��w|ͪ��Ja�����r�ߐ�) D.���l-2W��2/C�D(c�h�������<Y��7͒B
�V`.8�R�L��@�]�ʃ���iX�3|��URᶂ!oL���[v�.���/��e�Q�cj�V�U�(6B4�Z�@����+��ke��$U��@��0d
��W�Q���Z5p%Ґs�A/:�â&9��tL
1�*��8i��n1%JAH��i S���$�
h��W��\d�F���
�֦R/
���a.�a�ɖ�������p�`��@�n[+KSk�^O0!IAH��n�v�h��
ח� �;ߧ&����x	$"����OR٥�pN�v�>o����|3PF��Z�?��``�������JW�6rצK�ˌ.�}��~qe�f����7�v�=���9����3�\�;>:\��7N��ݹy���D�׾�{�Ӛ���E���y��no����J��1�4�\���n�r��1/��_�Y>nYz3�0~��)bnƷ���u���?���\��L\�sw�}u����������m��0o�z���v{������]1�go�^:A��sj�U��sYQ�s���j�S�3�R������ݶЫa���V՚���\�mO�\@d�!l;	��k;�u��Y�nE	A�������,q��pT��ؤ�5Rs�b���I�0Wj��5��eAK|�L��B#N��n�p��%I�N�[O��jp��[Ҕ�yS��P�S�EN��ӑt�"DpT:�%0}8M��l:\�@D3����I�Q��&0F�1Zӡ��jk�p4���1��5�j�r���Ðg��ƔN�KA�0�re��1�K
}��]c[[���l�٦Ӱ�r	�N�p
��H=c6�Y�LJ��֍��,˴�R^}R��z-<���)Cd�\w0/[_��&(٢;�B��!�GM,�B�mш�+�^����X�wA��a[H����(CdQ��m?B��&��0{�K��|�_#"��Jj(jԴT��+�,1)sI��aT���f��~�;?B��_���!e�q�P甕E���k^.��R���_�����1��4}r���&��������@�Ἳ�X�=t��D�|�窻{�_��\?t�����u��S���R�K4Ϯ=���3���\��w��/�8�w��;���/�0��7oߟ|��~uz������������?���b���ɥg�<������������oܭ��e㰹[��̎)#���[��]{8{�mi6I��嵻h!X6!��� w��j�d��S�RCR������2V@@"�B�P � ���R[h)&sl�7Q����
�����^{$��4�gFDF^�΋$6��Zb�f�ݻ@��w�������E�b��Ӄ����(��H�R,VVV�3�w�_uMqh����\ܣ�=�#{��	P�ukQ�+P�DU��\%��S���R���*�Kׄ4v:N��_��=�O>��ǒ��s�Н&����<���u�I���5r+������!݇s�|��,�ҹ-��xJ%��*d& \h̓�,-�s֬�ab�eH�?����Sn���A�Da�b����,5 �'�)��u�T��Ϋ%�1k!Y�l^�2
`QI/G��[\^�f3��N>����
��Z��`���-�y�U�!��Ƈ~覦si\*�$]<��hERvH:03�$���a�	x:�s<\B���Z���@6�A�y*\D" �*׭Nmu]F_c�ඖ�?����n�E �f�H�N:��4]ɬ����T8""��`ǋLFxQ�v���Ѻߩ�� WX��k�O.P���T��b��{7���z��Ë���������_������G'G�w�������;��������W��Ɯz��#��/��=���3�W�&�-�͞������	~�c��e3���~���W/_�n����+j�N��������z�x�:/W�>��֏�)�����"2:c_�}�M��a�ct�(�� =�&�L��h�̉	o��	 Wӫ�rjHB�@�`(o�*C_��Z�J�l�ݐ2��o�q0�I\��2.�7 �	I�(��V9��C�["�nád�� �օd��R��}V<����EX[%��hu�BJl,�'#N0�m5�.���pp�%,LE�`�vT��t Qt�L��kr�H��� 4Յ���k!tѲH4�p�)J��7~F2s	O!�Xw�
���nF<�b�t+�f�%�;!�4c���`�#��
�B!� �+�U�Թ��s5�aĂ�T0#rF��:�mH ]-/��,Q���
��f?ᢀ��u;�d���U+���
�b� ����\�]aK��)�����oo�ӂ����*Bt��B�&$;;�f��ȢEa��Q۴0
)��>�<���hbf��������E�j�r�\�\����>�x����\[��գ�h�Vl��f��d!ꑂR�.h��˒�N�����-���D�E��s%? �eG�kjY���5y
��ȵ�3��0"�O���ݨ)omH0BW %/ =^zlfFw��l3���u����R�t���z���Q�5��c (%6�DV0��6n�~暴26uʨ�����Q[�y��&�9��I�R4�c7N��B�*X�.l򳐐��*�.)����'f2��钩���sN�B?�O�.A�"`F#-)���m���`X��<J� 	��n0��m�a��<�x��D\a x�8��9�0�Bp���W�V�H��d�7���3�,���UyF�l)�0x��[�`3iF��?1^_y��Ԇ�.�9������]�9@F�p6�R0�2Wm� d�2K��-dpb�H���X��\�����j,14����ڄ�W������x%{<!���+Z:<;:�D�]7���2Rt!�)E�h��@�����f6d���b�G�B��L+��`���G��!�x�����/=��f�ş��wW~J�u����/�[�#ח�>y7~���W{��h�g4_\�����ȉ�������W�oU�I��N�W�n�x����+���W��ã��������Oȸ.�.��L�w�RƜ�{y<친W���]F��s�����ۗ^��ϊ����B;�V����W~bf�+�w�W^�ts���v���zsxw�_;Ϫ��r�w�ħ{�~D�_�^ջR��<;�o}lE䣂%E���C0�m]]vC��A����
)
�t��g�e�f��|��I��$�R%�fU7r�Z].��L��Xu�!c���q�Pіn&�M��+E
�0�Ė��]q�]0s¨0�Rmǋ(��}��hj���ueެBv�~�xsI��$"���]�Z������jX��w�*��� ``��"i�&PI.�0*�����R%���]^���<b2��U]�D)�»ħ% ' p�ed'0��B��.��T*@
��]Ǧ�-��	�"|�IQgUYdWI�K-�KҫM��b����ţ-\�:�wv��"a���ƞ>�9���~��`�$���D*.��v捖O�63̡��*k4�\��(0��`�
G�-���dã�f��΂�W
��ky�R1:G������P���}&��f$0�0�',\�͉Jl�V��ZݨԿ� "}%�x��qQ�����q.�2J)�dt`�	ʢ�9Z�8��[�}�e�0A�W��\�xu��������M���ý��ç�~�w����o�j}���/���������������Ǟ�9�;�}^�:�߾�Q�w���ܿ?���K_1r�x���'�<5�y�����틣��O�x���5��A�:��G���Q/W?��%����x����C[�����	�,ơ�4,o�jمM��l�(Fa@�#�0�~ ���ui�u�YN-��0cS,���S�Sj;���q.�
�?�m:�Y6;h\�(���H��2Q$�R)�6���+�K�
c(��RK�Xꐺ�K;�ݜDK��	ǡ���96<�֧ݶ7��-#�u������@u�Ƒ�)��Y�m$������Y�Z�P+�,��5K�L]��P:^'&��L�O*�-�&���W�y��:)�]��W[��"�f#E�2J�%b�NIمT|^-ao�y��ʶ�M�J���ʿL&1`�jc�k�k�7���d�}�c�)��)M
���'3k$�2�)2ri� YLc�XHx0Ɛ���S�Bx�]W�D�+;X�t�S�H�e,Vx��Z���L2�EM�]Z��V$��D٫Z�T-#	`����
�*�ZDm����敂�Nt1��ǢF �p���bt��!dL�",��N���/�(��\98:>9>�xu�������G��K�}��������ߟ~����wO����4�?��3��ʭQ?�i {������C��q�Y�����v�&�}r`Cl���~���<;�}�������_^��<�\~������r�h��3��~���'�>�\߮�o}�gYAD2��Y��6��)I�i~X���<�mv�<����ziͤ�%Z^��+�@+�pac��06KF�l奓\8���Z��0�T^ѝ,��EtR�`.dtlt�C��*�:�������b��NA��J�wcg�,��>���e��� �"�D�������^�0�W�kE�,@Y tC�1�.�X��$�^��Y�D��-����5�t�]a�3GQ��\�����Z��H!`��!6��8�ԣ�3���@��7�Vꉡ�uf/Qx��F�K��������Ko�gl!�����P���bK1^^:;�Ldx���)�$�%h��ڔR	��pJX�	(ф�N}��4\ʎG��FF����%�H��%/;|�0��P����(.��e�@��΂�,�tZF��e�@[�B�7@5k�y��MKb`�!*-c�\,1�.���SW[��ꡓ���ӍW�^����DKU�2�����@��Ѳ�j��ݝ�8S�~P��rѫ���T{ƺ�H!�I�q�s�"u�>�Y�+����9��R��0ȧ�	@��M�\�ꇤ��٣G�;{\`�}��Vw�̨\����ҹں�
���V�(]-��(<Z-�"�)J&s��L�\A� �BВ��[y�,ڲ���W�(.T�)�<,	<�V�8u�~�@ oH��Q|$���GW%�TO�H��zv�hy�̶��Ə2=p�`\`���_�*�Ȟ�HA��iOa��D!��W<~�H
D�����E1���i���������$TXH���ެ�9	�U8����.YҎ���H�Y��SKW|��ș}�����eg!	�t^�vl��e\�,c<y��=��2���'0{����P��\F*�0���]�o(�Mr��*�O4]�Fm' ���X=b)��1���lzwg�W+��
C ]�����ļ��*H�h��V���wEL��IDb��@��yd//L��,>:�3��A�}w��˻Y� 縺��؞��������}��ͫ���i���7�=���鹺w��`����~��od���V�<�N�����k�7w}����t�c;y�r�@��&�K��x�f�8����Z�պj����̽k_e�k��0x��vL�������'J]b;�rܱ�ݬ����.�^���)2b��f�����8�o�./���������Z}W��v}���[d�w9\�S�i�(cd_.�W�l�L^�Q̲c;#��g��t)�1~Q�v�F�C�	|�K�E\]�q@F������MK��hI
#�	�Y@a�]x:alNf,#o�n��t�\0�D�,m $0�5�lht�TtD�rYi�K
S+�8KG�UF]��L/ih��
�
�����US�0`�v	�Y*�p*�KA��	��R��AH��Ө]5m�FÈY���9)6^v<��F�K!o�KB��΋J@�\�
 �B����FJ0 FT�XR^^̢��]�79�0� ��_�" ����XPq%\,�B2b ޅ���e����L/��=��gv���O�x y��(֢��>��:'9;|�"$�x �����d�Yv�l�uE 1�6��qa�<���`�0!��({^jS|�7���sA� (�I��wĹQ�Ƈp��Iï�J�6��T���d*��� E���v�+��o�[�����u�QM]đ/    IDAT	{#�U����D�R�DI�T��. K5�93��9���_��N,ˉ�Q�����|`��帾=�F�1;d{t��~��O�G{�<���ٿ�CW�G���'���������у'ۣ���� ����yyyu~?������������� �d5�������|xy����>��/����&<}��x����٥���>�\�ohw\���sѿ���BF�f^B�bB�!�IfԶ��/t��ѓ tъ�Z<k�u��al� 粲j�ٞ��"V���v%����2RT;w�. K.����Q,` ���ۗ�,Z�)uDU	c�PЖ�>s�/V�Xx��)��a�W�� yl��}t4�����w����S��
b���>��0;m�`/{�44�����9�~�<#(�;v6$p��
7..0�)��3R�)!��� �SG�a�?��sl-�\a���k�Z��V�Ü�/|u%�*��KD����(Na�XR���`PSM&�`��ƢB5(U*�h�p��bEMyx�r�3�y��:߹g��RzF���e��ǧ��K�*	fB�"���6(��`3
�E� ��/#<�.�'=����S��W��t��2j�Gef�O���)/<��E�m��P�Z����94�v�	��UvgZҹ�f�R=Rӕ���± 53JA��0���Ba,p̃���ʋ��/Ǘ3�g{^��]���O�������_�������}��}�[���yӸ��\;M{�����V�k�`z���q�����v��<���ݿ�w?���g�w��/^�\��ރ�/���j�������������������o^]����Kj6\�;5"���i��6?��q����� 4'\�8px����r;��m�ӛI�@�C"��Z,�ɬJ�DBX朳�:�-�������qaK����Y�`�!(36%���DFQ3#��E	S"F%�D;�L�L�]r`��a ��a�(�چ3��]FFB����6%~�JV&oY�J��a��2��h	W��a��,~Fx��)�9yYDu��-�˩ *-*�ZR����0�
)��L��a�V���EKf=,�t<�WUK�WLC��%�n)��Z�2j�O%�C! �Z!�0G*u5������q.oxx'�ac	�6{�ҹt!;�u�;c�"�^ /c5Wo2����BZz��KO��K!0���E�K��[La���*	S�0��%�Xۘk�^D��YJ7�RL6��쌍QQ0K�g��p��ovoQ�6j����IA�1O#$BF� (��r�(	2��K7��(�B�Y;1�s\�j��,�&�$�e�+@�Z$�6�≟K	��$a�[��,����Zv����C��Neꕤ;�>�Ӆ#��I��e�:��L�P�g�264^�����"��Ȝ�Bl�h�i����te�<zR  ;/c`<G4�)�� �,Sa/V�`Z ������Rf�
���)#	`N�k!)ڐa���¥%`)s��8.*y-�I���xg��60UG$�`\0�*)��. '��� ȋ���к��V.���#,�<����2��/Q:�X�0���U�`S�`�
#�[<��Bgh�`!gHl�Y!|��`�Z��Y*W[���@/Qz��;cg���
h�	�m���5��a���5���޷{F�Q�Ś( JF
a	Y쌂!�Z0��b�B���g�,�0)����&��5FE�^�b�4��������cHDaH�4�*�C�-u��kII�D�vj�Pp�3��U�n'UJ��K/�V��KũXa�U=Zy!떋N�7�G�N����%�̦��E<�t^
�y�1�~zr��c�rl �.�W���.����������^f���k���<TG$o��xux��ޣ����{�q̉뽞|ܻ�����9Xo=#j������捩�2���R�8f�|�Y�;�j&ͭ[�+�W������`���o-V'�@���,�3~ul}�����;_.����ե獌�J�_\]z���ß�n�"]����4�1��1��un��F�H�s�F�2Kk���ո(����-6�p"�p�NVZ�Z��*r�����1�owW�20�<�Z]Ƽsh�ja*o�[/6��3;@��sE	P���k\\���&�+�B)x(tN�.62*�4*����@[3	�-Q�[tD��E�* �x(��Sp�R*�V�E�Wx�jqj٫y�nܣQ<N�Z"�� ˮ�P뒬I`$��V�	��h7�D�z(Z��!��Ϣ�U�� �d����0���7<��f����BT���N\�t9��sxb��&iM������7%#�n�E.�^�Xa�a�%)�&,]I�7�9�V��Ph�YDQ�FE���?�~m!F�F7���2�3j.�*�2cڶ�C����`2��D�n?��c�8t�ʰ1ړR�J��A,�,���M.W�_�������T^��,��Q��ڶ�\byu�������"��O����|���}���*��? �����}����/%�!@��/�p�ƅ�tt�ci?���V+R�*�R��CY�?o2�sǻh=��|���q������j����l~����|y���M��ç.�n��7��>�����/�������C�I�/_�<x��fost�p}�x��p}|�ws~q��͋�����wr}�������7�9��>=���w�<��7W����w_���N����}��g_��s��������z�M�>ޝ�[C6F$�-�	�b�Hz�bmL��fU`+-�>f�Ǩ�VK�ؾ�`����q�د\0 U�ARv�*�2J�nQ�HJ:@`]��N��v]Y�a�),8C�Q1��i��й���(u] ��ԥ0]�dr9>��#G���A��j�}��X2�mn�/E`��(
�H�~-�p������ n����Â�1���E6R�r�b�_����; ����¨��)Zy��(�� ~g"��P[��q�%5K-@�V9K���RW�S�v����3�gLy�͋����(@���R��D��������O�k#�F2j0v<b�2ۓ*BlĴ�J�e�EWK�&��e!0t��e�-V�NSP�r� H0ze�7�R,���њ^�8��Q�]7g���[����������XІ�a/��mu�	 o`I�M��}����R����"T��O
;mGǄ���D=�!����'�u��3����������7�����������wg��9�]_�p�H�\㏜+_%=�l��3��^���2����������$[ߏo\�6���~���Ʌ�f~t�:x2^�����o����ۯ������{q~~�:��:��V�w�[��~�2c5r���Y&�htf��|v�d�@�MZ$��u1W�8�B :	l�X��L�r��1���� ��.�z�pX���H)u�tF���N�R %L�
�kϫUCQR���Ƭ+V��t���شL<6���p�*$c����c^K���l�TR����	L�˫M0�WHy��u�z��!��+c!ZH^��t)`�hEf�EN$@�6KlbE��1���,IἉ^�$��+������X]TF:&��2��bS��®LAW1�"E�ʘx� ���/K ��¨啂���+]ސ��:ET0K��2fgi�q2�����$,\������`���)���3�
�=f��5��D�̌�=�cU����1um��0���T�( <�E��R��!Ŗ�nε�S
�G"�n����g�lF�(� 3@̿t�3KFl�+�(ݨ� s-��o#�X;�L�K�8�H��yq�I�*i��uV8 ]�XYD�r�&u)3��Fzs�tF�#2�Fs�0�bN�s�����v�fR�S:�hY(�(T#~��EB/*��XXR��ޘ�81��gTSZ���VOE��˫M)L�\��uFeP"�Z�Ζ��H�)g�,� %jh�����xa���GW]w�͈J�P�� ��%@T�g`Yj�`��"d�I"7�0`��o���w��$#�$�(`t-�����«�@���-j�t	<o����*{�fR0��0:K݅l�ӥWa��IUTH!$�6����gf���n<j��Bj� �%F������]�R�`
L���FU�+��C��&\6p� fwf��MKzl ���~�5�H����R����]F�,��0�6-s5ٛ� b+X��S�X���!�%��F	�"���Vp����(�_4�u�w����.f`]
���̈��T�� $����ʨ۸�� =�LT.-�VR�IJ'x %M�$H5��@�p�È�ђ�����v �𵼲4�����$L�J X��#�?�鮏��a��-�z���窻��;�\���=����?�y�O^�;1\��ma���b{G�u��?:�x��߼�u��G�?ǽ��#�[��=yi?��w��aN;����p�4�!ǝGO��r������1�w�	sG�x���#��>�\���&�e��|���׷�#3���\��s!��O�]�o��ý��ۮ#����\L�[���K�9�-�E�o��N2��e��	��gȹ@c,�,7l��A��b�3
�g�W���f�(�5�MA���g%�����QK����aX"Oi�ϐ��M�;s��)��E*2a�L��sΪps��K�Z�1����J�i�B���ZW#�9���q$R�2��T��e��YjT�+�Ƌ��ђU�(�ʬ�b�8l���Q�y���R`�` ��wO.�.��^e����=I�E�\H�����&#��(QU �(#P%��xH�Z0x��Tv���%b,+��K�V��@�t}ҍ+Wq��Q=B$��.*�����U7E��f#`rr�jS���\:��Ӟ26vH�2�5.z��%H��+�/Dk�0�t-���]w�}X��Ll0���ږ�3�$2��V���q�pu@as_�t��5v���+�9+���Z$�ƅGI����0,s+�j�R �mIm���1�tȨ�2�T�V��Ƒ��v;^n��Y>FR}��V(9�M!*h0��	�X���*��;ǡ�����龱��[�����g��!�W�^�]?x��;ݽ��W|>����_��w�/�^\|����l�}������`�ݞ�ݮ��������~{�p{s��?}q��Ź��Gw��^�z߭\>�,����kf���֏��x����k����_\�<�꫻���۫� �r"������4#5	4��t
1��)�	L��dO؁M���^�zn	[W�X^S�߮����h˺Km�E������Tn�
g���
V�D�ұ���t�X2����%Xy�(���+a����2�2�%�\E�ڥ���b6����ц��^�wDa��}�4�=��4�`��f+��|�d�6���r
����Ԭ@�@�N��P�d���ǂ���!26QB�.���H!E�+rΧ\,�eV<��>���� �e�ʂ���cg��H����Io�6p{�94@�2�%M����~�<r��Ҡj#Ǐ3Z)��tj3�3?��C�؅4�Zlbg�_w�g���+c�EҦ�E�Q�
@Ut�p �q.�7�O� 	{��wc�U0
�R��@�,�nɢ0x�zU9��l��a�o]f`.;S���J�9���g��\��S=%����n��y������&��ԕ�*(��D,Di!ubה��'�g��ϯ|�r���зP���s��yY�������!�o�Wwߜ^�sĚ�RͭW1����K]��ho���3����'��ã�7�ߝl?<9�-ί�y��t�������������gg�ׇ�ϱ�����M�������+7MW�+Okz��RV�'ǩO��7<�u��A�F��7: ���.:o�Zk��KiNZx����A�.��;jP5��I+�I��b�1� ��啈�6��]�+�X�O 	�(-�6}q��S�-�1�,ņ�-�QƲgԖ�+�ٝJ.Q�y�Q&�.Lx���K�6d�Y(�e��	��b�c�΁й���0��� s6ĦO�.�DmF�������9�)U2	YD����f�B��+*^�,�H( O0�4f�+i�FQhKWUtvFB��kR�� �(�^�T�<���}��ed5�c�:���J S ��,B���Ie��`'�k�0��\�����$T/L�\t.ʜ��2Vv�i�Uy�6����SD1��n���6�͑�T� 
��N�SɅ�0FR�MHx^��bu��)6��P.EI�1�P��<a��ju�*��p�0����ʢyc�Ze%	�Ւ�@l��OZ�8gI�a�[�\`,%��%\*�JG �Dqѵtސ$K0.�j��26
.���%p$-$*�ƨ�y���(�t��U�K�-��q�6	)#�`�(�����:�=�MZ�Q�7
����M�Yj�3r1�"t����]�1'^-��u��_h�Ɂ,$#L`<�ke,\[�����9��,�n!=%6mY�S
O���;�P�Œ9�f 3/{��@�Uټ3;�tm��ל;�`�B愳��U��(F�-�-;��9d�dѪ�,�%�(^)�ju��VdJU�a�3Kj���+��"KW�4���H$�`�,`����K�»��uk�.ݙ�X!���B�WI��Zvm1�gԆ��Da"�X�i�Y&m��v�	ƅmN�n�D!� Q��npQ�H���j����hy�����Vo5��;�+;�V�!�e�W^�t��-���`],{�jӒ³C��I������������� ����Y�Y���(Ӯk]����(!��L��S8�,R�8cQt
p�X22���90o薈�p�!�R�?-�
��Z���@�%�&d.x]�1��+��oL��D+�&�Wԍe�����խ1�l����{㝱޶w읯�S�_�^:{�]m�E]�.�J��H��|��`{�ॴw�VW7w7�7���������Ç'�=O{��O��VW q����uޏ�\je-�_<�����-���5n�o�Pjo��&��A�����L�^�t3���B���� ݠ��=P͘��v���˫q�����@�;��m7n=���W6�����˫�ո��O�7I�c�YA{L\�U;	���^�0M�(��G	�bi�I�'�1������U������xd�nt�*ɘ}��t���+O�@,�K�����̨<1���e	�K��ajY�'#A�XT�Z�i��,�O!�.:�8�]wp�IRl"l�Ys`�0؁F�X�*U.e�*�(vQ��eq�S`W�=3S"�*	�200j]�bg)�X$.GW$W�G��D �1JMa��.��j�1���RS�(M56^:iDl`�`%������u1ha3벃�L^UE��7�n.��-V�,iǙV8T�$%r�H��H��)0�ZY�u+U� '���S�gl�bh��
�<Fj�x \d#�M��Ts�g)�)��l��.;�����E�Y-]��:">��sp�P)�pT ,-���	rE2�Z<��V��G��+�.�.:�t*'�� ��eg��P�b�y�{���\������?��?�A�������H��կ~UVJǛL*��rs1:���+�p-�8�ck�,�C��x���\�w\�>��W~�s��
*�_��/�s��_���6���Coz�����w���O���Ϟ<z���ٓ����K��~w��x�|�zxps��϶�{w7�_���������{��������'����O�{��}��]�{!���z{�S���l��ܗ:�k�+�c�xW��]G����)����"M��lv��D���`4c��ah�qY]��۝��u#�Z���E���Ngnh��CN���#����7*�B�(ZB�(4
v
�\0t��`ڼ챱`9 %1"^-ݐE�V���ײ��Y䍟���4��*���M��;�ɤ��t��������qFp��
�W����O0�b���A�t^�pns*���t���G���t�)�.���Ki��r�����[R�)s�"�V���DI�3<�M{
<W��r�    IDATى@"hB�*_l�����F��L��\rArE^j��x����S�Hx%�ުA1��>��*#"� �v2ӹ���8�vKKJ��֭�\Ut�S����- ��t�����X`�����.�\�ӭ��`��͹�pB���qZk����^0�MN���`�R�����"��
ŊBe!�t�,\��g�0Z}5LL����K,ѕ[��2t��Ԋ�������;?����}��W_��z}q�������w����积��WO=���#���:{���7_��~}s�w�o}��wǼ��`ou{�Y���۫��H��|��W����[��~�_����b�������������]����n�}����W�������븯����������˚c��������4g�<��3�i�H����S���@��΢�L�6l�1�@���j	�氩"�<0yY�� ����QC^�[5���*ȥ���&\m�G[^�*L�Y��/Gn]v�8���u�6
z!r	?����d���@�K�R"�á`��U��`эS�6 *���͑����U< B�d�ѧ�n�j�`EЖ���TE`|s˻[</# 0*ޅr�F.:��6}�.%�I�Zlo���,L�-U�@�Ue/P�,��ظ
�%��\lYP�J��W7c��V��3g#��Y�����DM��T@����8? 檪-��T�.��t�� ����T�%���A�3�s #�*
�b�?������%j;C���@f7���t2�6��1=��B�5{eג�� ,Rk�HR��)G,<�.F:ƙ4�.�] ]�i��R����U���1�*A^.��$��>iu�]�t-;`��#�6s�����DNPAƦK��h��NK�5
z�J�X�ҲD���;���"���`LW��0��RDa���8G#��KĂ�TF��m���R%\QMe������hC*��Ȯ+�(�����2Q���d��+AE�ɘRƐ�*$��Xz�\��E��o亐0�*DU,K:XIY�L�3jax��⡰kq������Z<����3�x�ՠ�<"#� ^���!Fz�"�-��������.E�2��0d��i�*
�J�F���bc����J������n?� �"�XQUŨK�!HB��L,W�(��,p�OK4v��6��#
f-��Tºeg�;iwC2
+#p�� �OZy�lF1�:EU��*#!f�K ��Jl��(إ�m ��v7��3����f��`LI�)0E���pZ`o�������KT��~���~!Nڤ���nT#-����d.���v#*�E�^-VU�h��,x�V;W��^k uQ�9	<�����E�DR���]	�^�y�Ф��
�R���`P���Ŭ`h6^�7~X��o��7~tţ��g_{�Q^���<�y㞠?^���ޡ���x���h{��j�����L1{�c��}��;���?���+�%�ۼu����n�¯[�+��.=Fb;�W������b�(iD���)^z�N���Ͼ���q�~���YΞ^�7�� }������/�ܟ]� bZ��x�V����#��썽+o�=���~�s}����i<^��?�9;����Us�t�xL�S�J�Ie4	�=C�2�&�X,
 K�C�셷4s����qe�f ъE@T27�@;C��|4��	�E�-{v�������C�R�+��׍P#pH-�	���u���e��(����:y'�>\{d��P`��� I1s�4����:��wa�qV�ؑ�U�.�K��8�c��C�p�dGK��R
e���X�9�Fg/�t*�D�\x�0�.�9J����X�S���B��Rjى\,�,��kbxa�c�J2Q�=�E1:	�2^ųX�N�1s�V��<-��(���2Vv�j���k���(�@�re��� F��r��e��b��TkK��!d!xsψm��o�$Һ�a$b��z���û�Zb�*�5T�����rQ���e�.�j�,0/�DZy]#���F]�h��+�@��2�c�Eкt�"���f���v������2�~���HԹq�߱�,�7A��6�4m,��F�&.S�7�X`�a0� �Q��a�o!�ݬǿ�|�0G�o���9�v�i|Ih<��#ղ��yy{������w�ׯ�l���Gr��ә�w�G��X������}/��x�`{�N�k�^��Ώ~yws�������Ϟ_���蝧koK??�f}�����ɓw�;�'�C�x����?D���{�'8:���j����ۭc�ƹ�E�Y�����ɔ1��в�I�2���;�|��&�f�u)�W�B���0�:Z�����bû���d��.�,�d�B
��p��I2�m	ސ�Ɣ�0K��`��\t5�PUZ:W���,t"K!e���(��gT �0�%b䝉��N���W��o~���G��plk��&=��2��	� �B�������g�ѥPf.�nM{�ZB��F�ر�N�MX
0l���X��\M��DEn��R�B9�MF
i�x�1Vc�s��|�*Ov�m�0�7o���x�b�,��%sh���ui�|MÙ��@��f
*R�
%��K��"���"0;ou�3J*��y��G;�C�SF�
a�B������3VmQtB'"ݨ[D`�ͶJ��.k��2	����\�\���L�#yM�t�m�,M�*8��d� ��e�R@���#/@/�@�S��@T*' ��Y�ZH��2���s)�ސ�^��Z����������_��W�|�}������盽��_�ruq�ۯ>���?|�ݫ�<�����ޝo��M�K�������o������K��Z��ޮN��n�N��W�z��_���������/��|o�Z�������������o���|����l_�{�f����K1u�ݨ�M�y�``�4E\M�QK��T�B��g?3	VPH�&?KYB������A-f�\,���xlɐ�
�6ET���$œ��E��0\���S��%��Y"l��`S(!c<���!��ŀszY��rU{]-@�b�K�Ѝ0�J$j�fI��y��H
�T��*o-��ʛe�.��Sa�P�L1�eDE!��Dr�	�iA3��ȵ����2�]�a���]��k�˫eglt�НMB窆�3V��4�6�*	\[yt
WlZ]2	+ @Ij��b�e74�.[�&F�R�V�n�D�O�'`�K'�K����c������N���2�ɒK
.�%2[F 2����1bI���9
`.�T���4L
*��qn�j�b��>��\qґ�1!P��@]����NH�;��a�VF�Yb��@�ؓQB7{M;��t"��V�L-@����Y
$��T���N�5)U�G��(Zz��Tu���Nn�N�`�	N��ѥϤ\t�QD�`��*���!3fY�,��>:��TC`-NT0�����yk��&�2�7pI�!�`u�ިY�0P`�
�B��媌\r�қ��EW�'�=L�ML.��S��0��ə�El��y�s)R�j����;S ̱P0p��8���؁wy��RaZ�f0 !,�tm�W �+��t
W� 񳳰7�SB�YHv���t��)�,�y�¥�X
�3Wg���ȫ%����pJ���7����dG�T9 �N-�.�8��5W��I'bE��Y��A��[W�������N��y�y1�F��S�f�� ��^yt�Y����MI�Z�>1YJ�>?F�`�m��ċ��z;�0�%�S�����(	 �e���ԍLo�,!j�)�n.)J���Q�E�a��]����0j�H-����,o?�������;g$N;Z<0�Hy�'CF]0��!��,�4E,�8g	�xb�V�,��܇Ny��2b`��]���0�p	z� ��P!EE�"6m�
0��饮�Fx<`���
l�}���&��$�k�4�7�TZ���x����7�}b���~�K���k�݌?Po�^�{|su��F[�m�����Ft9s�c<j9po{��C�g�7��t赛�nl�=7�ҥd��5��tw?���g�0�}��F�e�#������W&|uu1�V���sAA�^�7����xP���MP���s	��޺��&��v�_�u�x}i���/n�my���,�Sj���`�0�a�'��I�%��o����F�v,��W������ &�B<�uʒC3&Q[HwԺ,��Ĺ��Y�Q)/X�t �\��	#�@��@r��.�7 :B�D���va֩C��*��~��"�h7��(���DRT]��+`�#�,.j�c��DN>�
Ѷ��*�x:�\I�T��옕G�*<��*����F�7����x]�E������=$���.�IJ�0�V�Q���X`�F���Ȓ��"!o���H%!��2L��]�JFIqF��.�hJm'�s`Fx��!Tᐁ�LrF!Z���m�x�LZs��^��!��E{�&�b����IB���o�u���i����d�E���t����4Bҥ�9�Ū��+�K��P �@�Ka��0 �����_���3[�9R��50��E�
�%Y��q;F
��)�'�|�&���?����0��^�
 �ѡ��h�Wh�:�7�sU`��,�(So�u�e�Ɛ���_����qʳ��o������y����Χi̍�����ݻ�?����[n�y~�ӿzt�=�wW�6b��|�|����������W�/N�{��嫣����w�~��������ჃG�L�̅��{������6���^B�@��GO]ӿ�fuy}~q�K9+�I�Q�14���I0�a}�͞��5�H;fn^vs�č��c-���2��RD(�M8A�����I!VӲ�8s���O�f�c����8���H��Z�j �k��^��@z��B�"E�1�=A�Л�ff��U�X]<j�D[��"r�HC�vY�b	湫u!ye�-g���ۿ���J�F�j]?)� i!X�.��,v`Yfx����!��"BrU���
k��4��)K��J�^�v�s�D�V�c�fc\*z���b���&�9�J@1!n�2*�EjcS��^Q1Fȕ]�$���HXt�^I�y�f3
�2�߿]�c7v�rI-VKJ!�-�D :;ef��K1�x�F2��M�a$��EN�e��2jy�c���)�R`H����_����$��?&�4
d��Kl]�� �B����y6?��h*�.)*IK�L- 0*��f��RX#�m� �o{[>��p�R�MXI������I��T�\�F�d��e��W������OV�>xx����7�_�>z�9���?�ޮl��/_�]��{�s�O�՝�c�4�����_g�=_��;�V͞��U�Ց'�WG��:���;y��Oq^ە^O����Ƀ�����gc�:`ǫhO�~��_��/^~o�EL������SL�-�x��4��!Z����f� y)>�1t��+-�Y����X�\RБ�#�w���L�ya�c�{�œ�E".��)թ�v#�eL�>��W;��0嚱B�TT��0Ѳ��d�.:��g,V8LsX=��t'9cY�؉SVu6����Z��&�>'3i��R!q��K+)���,%�y���͆.W�)���̲L!�J��.�p��fAyF��(]Q����D�24�,��f%BJZx�˫-c䍱Yj���pm��(c)�9]�]X�Q[�*ѭ��F3<��*=�� �kwh��/��B�C`Tv%�)���.�C!ڢ(#�rLaPy,!g7���o�!g�ʵ���BR�@zEE74.!�9��jZ& '�VpÉ�tc�0�8���C�F(�-���,�(E�`Kа3OB
�O�5�.�>��C~s΂��]a�0ѭJ'+
�����E��7�����E�(:c��b���-@��`�G�΋�H.%��Lg�,@l\�*$�	,W`F"�(zl0��K�5�,�b�Ǔ�.�R�9<�,S��<vx-�̾[d�����.�.�"�Nѭ��Y�
�SJ����.�.��Q��v�f��(��u\��P%u��]�XF��js���ըi�Q�"0o{��3�X��G^�\�\."K��x"����bؤ��yM,�5ǕR1\ �v�銢皁��xK	��۴D��� IŤ�-�t���*��3�XQtƦR-=��^���l	�'�l��o�R"�}R�f����:�k#�ˈ���Y@��1:e@@"�!�����F�DR�KD��֐����J����^���>��xz)v-Q���-�������h!��89��Nl�~�m�fg�J� cC�`l�$0������bd�K�XJT��,��Q�V��j�Ȉ$��T�"CFB�4�&�EH���!�6����6BJ)��pUIx:m��Ǻs�1M�%�8��.��X��;@|�ʱ���]��n��%|�ގ��Sq��Q
�⃻�X����1�q�g���uq��o��W�ť7�G:.��ݗ�Mbo�/��6� 鸷���:^?�̌��˩�H��������Q�F�^$W6��ח^�g!���nE�N���~���_|�­��{�.��������Q�p{}w�w���kO�z��v�����ܪ�(Rm�҄7�S��N�sf[�2Ʊ"x��|��Q6O{���z�yYJD�Lv�T�skU$X�v����v���y)�n逫Y�k�ٴ\�f���
!��nT���.�K)���ZS��:�&� ���G��4�b;`;�+�Z��&�K[�2�u�@���{ H]����%����:E��"�²�%*�N�~�.^QY0��Jj݄W"�\�B���bx�c#\����X� m�F��(C3K� ����Յ�P��TVͭ,�Ju~`��,����2i�˸+�ÄT�*a�!��<��d�L�Xw���(!0/��������52Q�F:�yY�.��.�lL^�o�����,�����o���m#{�Ye� 
R��bS�r���c�GV��Ş��u��O+ȋ�)��\j@Eq�q��Hi[�b�F��uH���A���F:�\Cfw�s�n�[_�@
�\��Q�;L0jE���H�%*�6q�`��rU�|�)�=�������s�`�4���~9^�.�oX�^�m��/����{_=��GnV��ۭW�ܼ�x�������������?����9��Ә�C��[=���A߹؜ln�8���w~I�/���<8��w�����{~v�9��}�js�����������t���>�7�Y6�kB�W��]��ͤյ6���䢂5��,Mi�&��1QΆZvTyM)���RN8Ų`Ck))Z+�*�a c�1�A=�	�a0u⑅Dg��E�+)<��QKG�]7a�1�@�	�M�`K78	�Q�)�t$t5�<�;'e�03<d-`w!������`�� ��G}���;�L���z���[�fL��D���¸x[D��+[Em�U�+/�Xt�I���O�I�|�/P;9u&��V�-�!LQ9*.T>T�)�Hg�HUMJ!j�w
�����P �ִ�HGofȢK�(�K��0 �~/^��^_�|yo�]��Q5��<
#Q�E5"{v
Q$�q1��ĝF����@j�Y�t3�!�0�0RH����0F2-0tl�[�b�;Qa�O �z�y[���T�5ҵ���,~T,��\::aJTHx^].�uU�6�K���R��0�����A,VP
�L�1�\�6eRI��Ĭ�ױ��U?���g_~������ܿھ^�ɫ�O_z�����o`����Ӄ�����/�~qz���~t����G9V��f�n������ Ǻ�t��}_8���{W�#�>�?<�z���/���7������=}����C�y���������|����z���*���*o	ݬf7���\0b�,e&��M�i��S ���I�.~` B�6�0Yt���Q    IDAT��W�����_jW�L�$S�/�d�>6 ?~�?���@��v�Ɇ�>::�iQ�Ⱥ����\�]�<�I"sĈ1�Z��r��L\?|�B�,
���a������pD���s jM�Mh��[:8ešÑ�M�5���_H"�g��,�L95ӱ��	fW����	��p
�
�ᕫ"�B�KlEB�9���( K��P��;.�������[K@"�@�5�m	�R�@���BFP�#e@
%B8��qj	�B" �5j`��E��ZBE���h���3m��`���ckc�x�|AJ�F>'���!4{�5q)h�A��@�rZWʉk�ө�1-�l�o�ɖ ��ى3������)�~>�BZ/?��a˪.�f�o���' S�aj����8	�����ݦhK��zՒ�t.G@H��E�]M���G��[�>��#X�5�"Z	�p|��pv������R���&��s9)wJ���C$��y���O�/�Ni�|��Cx����I��Q�����QY�ʥS�=G 2|dS|:�����@��9���V�	B:�h`�P��@�o��vՄ�4f|������٘�BR� Q�Vs0���Q�|�,�y����)MY8�|L��gc�M�5��ҥ��[d�p�2M�VW�_b
pN��Ë�8R��1S�Ni�BM��\V6�Д`M��s����S�í�_4�,���r�N�Ur�jB��ӡ�P:��>N�*�����vR�"�S"�ijj��.�m�ꁈ�Y7�����V� $1����,�P��v��R��� &;��E-���c�FSNj��i����Vd��*�z��F �����s��-�h*ـ�q,���u� ���5%8R,�t���2�@05�2Ĩ+��, Ǵ�"���]��B��J� $ȆK�1�(��#�� 4�Ax�|�II1�a�GڷJx	�\����%v�ɢmb+�2G�mզ�v۞}#k�5*��p�k:}"�/�Zt��Y��;4���v�Ff%
�1�h@�L��E!�����h*�-R9�BQ�ҩm�?��r�֢�w���O�X���ھ�N����ݴ���u�������p��=+yv�n�����M,����O�=u����l���ۊ�.������o{yX���K��EI��\�k����(����{�K�տ��kjS�+����J�}r��j}��}k��6��[������?����߭��k3O�]������l�]|��O�}�𵯽�=��|w�43�U�v����7p�����gk�2�>��觀�vG[mc9���m��;�:/�s�c�0�p�MK�ㅶ���/�NYl�5N�^�F��+%8D�"qajR�31g�1��;Q����X`��)[���S�nw�ү=�Y�U�]E0�%(t88��Z2дn�'}�&)�"��B�@���i�wz����D����H-�py'�Z�8.@�������e f����-M{��:��O��\A�Bq���
1�JfuX���	�ҩ.��hY!M��ԬT�;WBޛ@sI�Á�0b��ZZB� 9��_
�Ҝ���F2���m���ꢱ�0d�I�l��v��9�#b7�-��� w���X5r�Wb���q�iV���.�S	��\�ae�#��'�pV��;ʎN!Vn�h��Xc�q��D�H-��z8۝!�e������*|6�Cr���t���=�N��֚!
�
�rLը�Y��u�#�`Ԗv��[��v���η�{v��똺*�k^O!k�֓�Vn�ӕG��=~q~wq|u}rv����U;%�}��[\ssr��f}�s������̓�����C�|;�۷�4O�۟���S�����q��}&����˯�_����5�o�ޭ?Q:;<xrvx���o_�����8=�D�O|�����FÆXu��)j8v��� �m�c��!8c3�ѡB���N�s�]X'��pYl� �ܮ����Nm�:E� N��A� aE[�f����X D�>�-ʴD>�����J��EY�u��3G.�H|�(T�#9�I�Z��݊��Ц����́(]���_xty3�c�3���uD��y��%��m8&٪�B4[���ԶiG�����#UcU��J"� )���r��� p@�I���c�)��AߒS�p�cE�F�I���-GWR��H���䇫"wDZ+�Ef��.�9u��o_�gK�C �O�3υ�#BAh�T��|L~����h��"���F8M�t�b� �i)�hD��v��2�R��<*
�yd���pR0����8�9���A�>M�PK��BIq��l�)͖&+�sRc��&Qϫ�V���hNNm8�ʢ�|�'Azsd�����1Y��V��gm���(��Ի�����߼����|
�'����W���w���z�X/��}�����ɣ���|s}syr���Z��1�z��!��k��i����*�Kq����\��n�����G�����'g_�_��Ϳ���޿�.������_��o_������_��׿�կt���6��[k��"�B�-ٔ���=~�R���7�7v�W1x�c!�ĪTh�Q���uP���8v��i�eE;��#��)�>qj���~�D2�1�)#BV:&�(��s��[Q>��.��d��<��+$�C�r�#E�︋B���XYR��[i]��v��%�혨�ٵ-�~j��	�dS:k�N1T7m��:��1D%�j�@JǑU��hpc�\��L"l�kc���]ͱ�+D�&!� !�8�b��|�h)B�p
�gk&k7�E|KZO�t�����V�6��bJӴ��˒^
&|�[����Z�z�X3�XSYʡ�T�CAh��w�����c�b��$�&��B8�E�Y
*�rG��j_V]�4m���Bf���.Š�OVQUT���ZJ��Q�H'���*$��dqp"���B�p�h��B��۽��
�(9~;&e�I5m����D0�d�h�B,A*�c*���VByw:/�#Ko9����P�r�^i�J �y)�����X�r%rL�4��r1�UISuSY�9υ�m�,�@j[iC�n����?�t����T+8=W�T.�MS�Ȝ��=H�:}��'�P�^6��b���DÇS�с����UH�3�3Mz���۔�@�h��|�iUR Z�r��8�9B-��5�\� W�MJ����Y��e���ڛ=��*��k@b�Y�ȑ�c9C@6�������9�Lw;Q��~�DLU�/�o7���4���7(@�'R��*�8Z�!�(_M�U/Q?\{+��������ΏcZ�3��v^�BR*T?��!���$� J�4�q�������B�٢�B;o�RrRKY�f��26�eh���
����u-�,U
I�2 �N��p��rˇ��4��f��F�rr��t�o!�hm��n��/j�99��?K�������ix�ԡ�\w8�c�VK"��F������kU!dR�" ��55�=}x��Bj�#�Dj@Q������2�/�e�nE�@�ƊF r�"nD㬟;X��\���ެ����L�n��ۄ���G����_z���_=;?=8�;��{r��'���+���_����~o}��gJ��x�S>�#|�����V�Kb�Z�v=,���C�ۋn��i�'5(j��j}����5�9ҽ�S/������G��g�Oϟ�H��7��Ob��>ۿ���s����?y"��K�n�8>�Ÿ~r�ڽ�>�J�o���N=]�Y��<>I��n_��c 9@ƿ��:NM�^�i�l�]?���s"��W,24�h�Q7O�`�KTǹ�%�Ԥ�. f�C��Fm�kc�~<[��C�(>� �9�J!���7���?�r��Z:�ZMM��#H�=j�E0���X;M�f�6J:�i�hmQ>ۿo�IP"�!
uWD9�aGH�ˈ����K�|���b�YjX>�>����N0������ڰj��m�����)�ڴ�:��
V?��q��Ȭ�G�@�|��䶥,$e�i&&����1����|
v���͆��Ro���Ԋ��*�=d�O!�r'��jbO�]mu�|~4j)����+�3��	p|VbgK�$�lȝD�������@o��ڕR���)�:-�td)��ꆐ��ɣnE�N�pj� 9��o��`�2�5�o@X`!'��w�bJ��0��>��z[��_�Azor��b0G�B�%u"��^����4��A.;N����BD�é?�-R�����Rv}5���9�}���ݳ�Z���_�xc���GGO~�%��۫��'�^���Y�ﾸ��;8��>:str���y�==����o^ݽ�>9}�������՗�����w���'�|������go�n������ޞ5_��������_޼�9=����E'�C���ɽ}3��ն�v�c�r���F�����a�vƁ1EvxDM�!���Aqt9d�.���`��*��)C��ARe��ށ�_Q�S95�{�:�R�*�P�EP�5
qZ��\S��pR+y�MSȶj8q6�Mf=��*��D�3eL`�o:=p��v,}jM�,�Z�De�����C�o'���y�͕�O�f��8^��ENĴuI�I�T�E�hD �y����I�S5�h�L_�h���������>��ZN]9H��'�Ί*�涃,�&��i��Ԟ@Kt糘����p����&W��9ߙ���we���S�w4e�ɶ�u��K������5L�F��E�'Uۦ8�IR�YH
�B1[`�p�c�(��j����%���LB����\�r�T��#��;� ���
��|��\=Ȣ��I�_-m�S���BDe����í�>���soZS�&ToN )h �U��%+a+�����x�?>x���ߛ~����l{����Xz�t��dד���;��^����W��7��p\�h�Z�o��?����ڸ?�[�Z��9������̿L���������7߽:�|��������q������\�?����z&�E�6�]�9Vd-�n���q ����J7�,�#n�L�����=j|�\��)�r$k���I]Y�Y�D/�����y"���s�5��:��8d&j��+�`��Qh�1���C���:����Q^GH�Y�> �WQ��0����"b�CA4��ݽp�rR��$�43���ml��"��94��r�A���b��� [u��I���R75NS�����9�m��/���Q���e̔k�nS��C���һY8E9�r��~! g��G#��I��.M�ԄaU)Z.�(��_,rӲ���9���	I*QnIG�A����}�z��*�$BP.\��ϧ''q����&�V�tSC����pSt�5�T�%�0���nC��l��*�p�e���|V?D\��3��,��,;)4C�����9�hqj��"���heU�He�lu�F�OJx)BE�p��|��UM��O��|�����Rpؤ�`�d��ҏ	��n���xp�D�j b��!�R���b�T�p��ȑ�-
�̆�;R8u1j#5�(��V��ϙ��6����t+�tќ� #N%+eM4|@�o*:��n���6�ϑ�����i��r �8M�jUW(d��H����3�
QK��t���h=T1rG
�B��fB�LNm��	۞p:�p($�VBaґM�F��
a���g��9x+j�BM�ڄV��:�U�/�>Q#������`;ꭕ򥄔E"J��4�N}��7�؈�W�|d8)~��%=�fEk�?G���������B����Z��e-SV|~uٞ/�FI�F)I�o|��rY���̖��֔����* �����ԧhU�$NS�9eU!�#��)8;L_�����9m�B�d��ؖ�V�io�S���M����x�i,��x�#�e�)"r��OV:'B]�G���+)7p�2r��m����@�}�d���%;;�<:Bp��)U">��aq*v�"4�%��R"�BlS���6d�G�x,(�e��s�M���&����[/�qM�Ή�������a��������㇋�����w������蛷w>�rqv�������=������w��\�eߘ��//�����w�u}������H�d��s}�߮�殷:�b�{ہЏ��OMz�ћ�������>oJ����{�����'GO��]����mI�yw����#a�C_����K��Ţ�4�����k�>��8�}�����!Q������b�՞G�����%�hu��.�h ��aq8�p�)�( ��E�t;�8��Jq414��Gn�9��4��E�rq�8���	�6rX!����B�:��l�үh
��(ݲ�pl�u'܍w�c���]�ҘV-L��)� �R��ʲ��A������Pa)�,��SN�]5dS�hm�'.\�Rc�!�mͧ,ŴVqDeiX����U��:�1�=���B�p�_׽Y������<��
щ�C���q�iR��y�h�T�zn[��
K�[Y�1LG����E��D%"~�t�^���'���Ϫ��~R*��/�ZkQh���5E�d��@>���ו������Lg�&~��1�g�R�ܹ��"S�U�	 Rn͔G��GS�B,^Ϣ����P�-�2�\��������b��d�u��{\;O����ݴ(�3D�������N}�?��?��G�O+9�Ҫ�o`��i;���-@%L�hW�R$B֓Çg'�f)4�}O���qh�<����or��Ϟo��w��⣽��gO}������'>Rz����������~�3�������uG���~���������ׯ����W/}�/~������ׯ��y~�~t��U���ԁ��~����o/�<�nN����ώ��ܴ?�ٞh�ӌEm�Y��%Xc;��	,N4҃�\Q;�u�c����'5;A�Q����VK9j8��"UK� ����wY�t˻Z�q�.(,q!���B-p[�z�!h(���Ae�6�M�!� ��2�r9�`����h�q�n���2pL(cVb�V"��"��fj6��O?�Q�6�'��~Z��9v� �Q��|�a:����cV���4�����뵇���j���)��	��J���dղ@��#H�Nbj �-�NCEʵWB
�#W&k��	�*���p����zԡsթ�,�^���w���l�֤WQK��e����V-V9>5�
��Sh�X�m)p����Q�U�4�qୗ8!�h{�B%�$�,$p��@�Hq6�㓢i�f�CU �CY�::p�@(p �Ps������<��nȊ_z�,k	4�@F��IU�,M�<:8B,�Cp�q�6J|"��9�j��Q]"�c9�C��/|[ͷ߾�Gho޼s�V�6�_���ͻ7��&�-������ők��"���7�W^�y!�e��� ���H�������>x�#�'GOϼ�y�w{�p�p�	a��7����z�_߮/��hГ��M���X��*,�cV�v��e�×eg���t����7c�@;vޮ"���/�=��Z��D)d���Ҏ�#����_am�� �1�����#����pH�[,�z`1k`��K�P^��C�t�A$҇C�l������h��7J�e��B�4��l�k�cr�y�������$��\6GK��)jJ'�2��IM�5Ukȵ�&ȉ�6���N	��!�j�F� ��Ł� �Ds��|ъ��B����<�Cp�R�r�Ѷj�̩.�{Y��f�M+A$2�����lY�D)�rԵ�FJ�\�d��蘊Fc���-:�Q�\)�ZI�Y�fDS�G4�9��$�&�0>�_��˻K
h�n���B9�h��Eփ�R�a�pJ�yYp+�C��5 1�h5���y �!(�rB��h9l�[�ڐ�s�_9":'K�T�&�@�#Vkt$�hҋ�98��Br�%U�8:��u�+�#��/7D�7J�[:�PYI��� �ƚ���y��$��8J����V��P~�0�y    IDAT[��U���H�ZBKsB��HŔ^���R6%��Gt�pjl�rӗ"��)���Bp��pS
�a��" �eB�2�H�2���B�K�e�s��F4��^�%�[lK�Ɨ�)�&H�*��9[�k?E�#�X�U��gww�H�m`�B�Ek&�z`�lp��`R+�)�Mvp�@!Y+*++�BL)4���ã����S��Kdk;�r!�Z�Z!��G��A<?�8���8!1�R����q�I�E��Y/�-qD8�˝��y�$;"E!8�)�A��=�L�l{�����Ĥ��NJ���5D�-�� d�T4����8���#�&�)K{|���&�$[zە_u�[L~��JѤX�dE�f�^]�'��9�%��$��B0�[��3���� ox�c�َ q#.G��p�m�G|Q/�&����խ����RQC.�r8h�!G3�ϕ6�1�(�z��(�b���#� �����k��_D4S e��J�f>�(����:���`=��ߑ�%�-Ew>��E������������m�� ����U�7��)ʋ��>�����'0���;�>?r��~��g�o_�yy�[�z<����zx��t}s������n�\�?���J��'��'���Ӿ�X��A�p����k����Q���g,-������}MO����>�z���[����]���]��S��^��_{��Zzqgt�x�:��\z���n���D�g9��؜[�_�m�������sLXG�u��uz,��-a�Q_m!���G%"�!�v_ˡā�B���3Й�;�D�DV��.Z���,
��c*��A�b�ő���S�]P�
�W�E&R�4YES�7��@�^����}��ǈ����9m��c�TQ���Q	�f�"�c�C�eSjh�u�A��#	��I�� �K,]��B�z��(V!���|�JQ��!�2M�AtZ�.�6�+�H���"WΔ����16)on�&K�$���	�2���Zƶu)K�1��AJkD�6=��ƙ�����f*рi��gS6�,p����Ŵ��>Ǫ��t�*��m�NQoиq��vhQ
J ��(��Qr+A��7ő��D|ӚM���d��'%�ө�a�щS(�ĐޡaMqXm�E��b��z�k!���8\�!ZQ�iҩ%D��[cۊ���.dL��%�z��D�����?�s����>,I����J
��h|�@:R�Bm:�_jTݠ ڒ���r��^��V��������������7�}��v�r��}Ϯ_|������o�x��M����/�^���4���u� ����/�<��{�gnn�]_^<����S_6xsw�y����ۃ��T~P���g����S�ݕ���ߑ~��x��_]^��O�Dp�?��C=w�ڊ���X���dtj:*|�	!W�E���!�)|R8.4dY�#�ƦA#l��"��*��9�dZ��?��?PEE���q�s:��S��\�:��:h�KD��hMKLn���Y [���pJ��ݵ��8��Aǔ�aQ��BhYjU���R�rF*�6�c�!�NR�e�X�`�ɟ���|���~&�#��qDl�ZF;�����*�s*gc�-j�-ʨy��5`	�fM�zn���<�S�[m�97L�r���E&��J1�6T�O��X)�-�/TѲ���z�;']�����]�Z��uK�2K�'K-H3Y�18u�Ɣ�	����G3�"��B��R@h�L��I��!Y�j�X�%ҙiQ��Kw�tw-��@s)���^�9E%u�Eu."w�x�w'A]	��f��cXK�Bt��d�*��t�r�wtz�tm8�&���г�Y-Q��HG�C\V+�Dk���	�滄脆B����?H���w�/}?�����뛓�c/�}�����_�\��N�h�ʧ�o}?����?��θ{o���a=:<n~����ų�������م�Q=�z���9��9��޼z�:���[Ǣj��r�����Gf-��ꃂ�������l�2<�?��3�>���A&�>A�F�OL����IJz{���C-���K��d���$n�˪Q!6e`m�@��*9pr"���� JP�&�����Z!��FY��щ� dC�b��cLU�AÇ�h*��P��l�i�	J��,R-�_m{@�%b�IL�����Y)���������fP3���<�$���S.�>�dk^�Om�#���a"��!,�4�"���hF�&Ԙm1����~�p����m®�PmT��7%b�>�a͟*h�K�#�%�ρ�H����g'�f�-��j�$����%�uˆ�Z�W���b�A��+�F-<¬�H)�!l����T-Rq D�j��I��lY�Yc�6���P�,�r)$5���T3�::A�F���@�]M��!�6��x��Q�Cі<��e���Q�d�]C������#�r�8��h�PQ�����4�_�H-��������{��YC�����2|�f=�9lL8����pG0�������Pʤ���)Pnd�Y��D��9�Bi�M']t-��J8��8R���_n�$J��ڛ��5���B�D����h���Z�4���>�DSE`48eH倜����j��O�*����B�!U��?�C���Ǚ\����Nd��#>�\�� W�p
u��>`��ӱ������ζuq�@�2&���\�ZӤ)&�m�@�)����S��ï�I�(
���oQ�B'�P�i����b�JI���' ��7Տij��� �e�s�1S� G:�Ѐ���WI�4L��G�VMk>�M���4&�*YQ�嶮��'�t>�Ҧ��>p[ƴ��FH65ѲD[&D��h��Q�_H�Q��g��ΐ�N���%��?������!;���?��_��9��d�� ��sv�]�I��7�q��w�V����9�JפZ�R�0՝q�.r��Y��s
��E1kZo�QŖF��&��v>И�u��+}r�R��O��x㑯�����C�g�F}�ħ/��0�Kűw8��O�O�r���������w����>oΟ<���g�������}����=<�#/������ō���]I���Sw�����O�K�8���o��QOm|s�%���]Ƶ�u'���=���nܼ{}{~�����X�}��m+�������97�W�g�e���ߟ�=�\{���}��~i����~���N�O�ȑ�l�X�Y�}�צ���8:J�!�jG�1d9����8t�Bp�8"����� �
�4HG�Z�� [?�84=�^�ӯ�X�r�����c9d�sE��V-!5;O�I�T��
�����SB��I��|"��=��nE`���a񓥏������Ui�M�J{����RM�Fp����Z����L���ZQݧʼ���Y�*v��f�n�iIT'���/��~�)���Bu�V9��!}{b��ɴv%0��������jN���J���ӥ�ވ������R��n����3�q���;dj���iU�����6EM�U�C��,�P
cU��Q������Z�>~�b,�6+rJ�vǺ����O�}T[�Dk/�O�P�����A�W������60��-�r����2DG��O~����𾒻�p���ڐ�\�@�*ү7!YԈst�����N<����#ħ&�n�ٟ��G���U��w�y�~���o�
s$ ��F�xG���i+A�竴���b[I������9��c�B���g���w������܃��7��7_<��K_Z�����|��g������_��>���/�������G�O�8��~������6W�/��z=�^?�������o�3֡g)�<�b����w�{Wܾ]_{B9��<���z�or��p�Ѷ�EYQ;�jOZ���XWko3%
!�ݕ��\ȨA:�1�0�v����BW�#ׁ���޺T�V;�.�\�tr�U�2�*��#�Wh
�ǁ�#@L�5dMb�p�|Y����L�G��g���'<&K3��b��EsQ?\���a�yx���������G�N��(�?sL=!y��W2L�ځ��B��I�K�#��!��G���@�!8��>'B�Ѥ�b�
!c
����e!�gÑ'� \�=g�b)+�v�B���s�$�#�pr���k�g/��kUQN-�uJ�Ɓ+�JA���G�CGRX#Y�e%�7F��,�|�?Tɉ�&���f�*����+�n��Z�t�.˶�D�Hw|YC�o**�pDh: hR��@C-dV���z�R�(��*�2D?1;Y�ڮ.�ge�b=���ܰd)F�2���"_Q�U�3m�E����
���r�ŋ���������w��߾{��2~�|z�g0V��|;��'���nx%���%�9�Q�^=xt�
ZG������d�����ɓ���o��^����]Mr��������������ޥ�኱j}8���o�u�7�r�h��Lq��� ��/f��U���o߀����=��*�=�5C碎)u%hA�Q
�S'�4�L�q� �#����hqL�����2L|֔�"����Ro[R�M;��KW�BȥC�F���0�f+�R�.j��]Ŷ�o��A�J>�*��@]9d�dO{E�lE/n����z.T@��g�@!�!�3�U���R�3�[��@�g
	��"\�Q�f�D8�)�@���X�c��+�#��j�8N
�Ȯ�P%
E+�2��Uo���pN}�	2������P?SK�_bδT��
���������Fm�n+L���@�Mg,P�BEь�;j���ޔc��� !R��;{���Nb��NŪ�R�d!,�����!�6�S�:�	��#�Q%��ɦ�$"��+4�6"�Ʈ^���h��J��`n�Gk�8,k���8��B���'�&�P:B"�?���j�Ȣ�pZk��)�(���jm�5PTJ��xj����L~|��9��Հ��w8���;�\Q�����b�L�156������+��&(ں �`M�x��HA���V�5eX��(�,��8�� ��s��`�
Օ�F�/��T=d%����琝��T�)��l�����:,T�|��B���1��Ya*�Ȯ��"���$U��Q�(#?q|����rD+�3R#��������1Q���N	!>����1����Z4�3�r�#f;ɟK�4E���ũ7v�ǉ0�bT��K��Z���6؊��	q�N�����7 U��&2_���� &�(��l=�݊�}˩bQ~8��C��C�
��S���{(�CJ��o7 -3f%f!)��� �6�iʣ6
���a�C��Iс�'\��E4������E�W�5�>~S4�N���� )�|>V�y��U�()�M�q��u�&�!��Y:��~���x9�PȔ�L��h�~�lO@��R)��C�#9�h�j��V��]�>(����-��S��'�+\}�7��N�W�y�z�p�1�������������ώN������ٝ��D^��������o����ѻ�//�<�yػ|���z��o���^_�Q1��H�9p �ѵ�#��Q_���Z�N���Y�{b���Z/��~�}�wzh9�6כ8Vz���w_~�s)��z6��@m������ͺǇ~�;��o}�:�;��}������O�>�������ݛ�_�{{�8�����ͭ��G��p f�9
͙l7m����t&Ha!�1>2f��,jD�n��p=���>�i]�����gW��d��n�Y!��A氣i-|� �*��4YB���i�R�0�ö���*ǏL���R�_�����v�H���2p��a��)�LaY.ݟ	�閻���|���J5W���+�W���!H���Iqp��)��r���Ƥ;��V�p�UH9�@�Uȴ���-P"AKSuH�@Z�\!#��|u]H91%B�y����Zu���q�)���uB$�_Q
��� d��m*
�^��Nx�����R |���� gSsp-��	q6��o!4EI�3� b�b�m`��s�8�J8�s��R���罉n��AQG��3�� qTѿ#�������O9��|�6��J̶��,��*�mj:�BޥҭǑ�K��Om��ўsƛ����>�XH��H �H�
Q����"jX�ɡ�i耍�i+��,~%�0��:H�2[���g푯	��7�7�?���۫�w'�o^�_~�0/>����7O.�OΎ�������ϣ9����'��o_ݿ>����ϟ?ܾ}�Ż�{_�ݽ[��������������N?~z�ď`��͗T<��y_��}]���Z���~���
�&h�f���JY ���%WI���e�����6�C���)(��#�E6�}v�Mi:!H)�́;�Y��w�M1=x�� ��rT4LUA�c$4К���H�nY�BYSR8F�ɲԖ�6
�hchrL{ȁ�&�s��N�q�����luV�P��:��bd�ӨN{%ʗ���x@�؟�����7�熿��w�	D�׉����Jk��)YL:�|�.7NQSջ�Q�pXQ.�Y��O�ń�r�c���8�T��1�Zh8.���U���|�8	=�\%�E�݀�E�@v�Z;���j)���:�S:�6�פ6Lq(L�{�($2_������)��IEww��C��B��[��)�#nTw��IJ
A#�8�v��A��h��g��2���G��
Hk4�LMij�pX�����1�Ⰹ;��UGJ
}{E�A����c�����#�爪k �!�b�mxp�z<z�|����{K�/j�M[/��cy�+�����J���S��C?!���^��P����ݾ�v>��~)���U�����1���?�����w��j-f{[��؄Mg�v{R��%lZ!S�����ۣ�5h�KZ/Y[�7��S��ؖ�x
�3}�@�d%Z�����[T]M��=��ô8Ǻ8�MG���8��0N4��V%}�V��'���|x��SK���8�K(�(djS`��*RD�r�S�SŲ*�A���0��q�~H�L[�8����9B��Cfl��G(!_'!hR��Hm�.�=|4�5fq �>����"]��R>�C���B�ud�b�.�0%�,"	"l���?L��Y,��>T:��N�R�Fչ�q�pH-�:&���[�M����)�ZYCT
[?c�Z������Ķ�,��܀��EH��i��Y�1�*e�32�B-vd���2r��`YL��r��B��FR|8L��#c�%�ٖ��R?Nk�[:�D)GH�5BdIG�cڿ�ҩh�4ݶSQYI�3�R&T�D�֎���"Pʩ�8�!�*S���1�pj ��s�!�Y�';x4�1G�!�4�YN�Ttצ��P3���+
�Ҳ��z0��:�C�!Bh1��
=S�� ���
��$��lYEMEٖ�_�>����j�E3 ,M`�EY:Bq�LS�'n���#��$��B!�r�eY8����qR@�� p�B�!��9�rG�P;\bj|�I�t�q��(�V���7�u��"�+�4Y~�t͐�A�*�6��%�H�I�?Ӳ��j
�.�1��n.���r{�K�*@>�r�vh��]�4���t3A6� ����qD�+Y�G�Om�\��V�%HD{��p��c6b�;�R� �qd	i�:� 
��:�D[�$�3�ت��"bR!|�Y\:$�r��	o�U7�[���D6>}Y�\�6�z���Hꁳ;���NJ��B�������_��_�C�[5����-و<�U(�BE�^�Tҋ �F[W�+��a�ߣ !��1U��g��:^=w�@0{HV7�D����3x�a"�gk�M���l�%p"s�zt��Yd]������~��ܺ>r��l��������g�OJ:w}fD��ى/	�Ꮮ=����{��{��7�/�<z����͍��{{��
�������E����x}�����m�;~8���K���_h�����ڢ_H�*~��~�S?�^�w޺K��7~�l�ە@    IDAT��d�y,�su{~�p�#����>�郤�B=��]��y�pyxt����{7W{~�S����r$4�o�]�/�3�:��E`��4O�~�����&�6�c��@dq,���8�Qί\LxN�<����� +�V�a����/=��v�� �H6��YQH�������!ŏ�N%��G3p"[H|�i��B0[)��0��d�@+b�5�m}�kj�T���&�!�ɽ����@wk�[�7��u���%�9:Y�)�+��)��w����o8u޿O"�G��.Q��$�@��)�}S��+M��(Yz�Ԁ�^�B6
G.};V��֒�+�c��ڻ�_V�� ai�!�	a��S]H=����õm��z������!YlT�(���S���,���>!���l���!�|; G�c!'��w���g�V!)rS�"��B��� m;��| �D%��~�
w�Ue��a�E�J1�dv�޽z6��O�����9y�#׌;:S:Dt��41�����F$M�YM�9��\�Ӭ�B�Y:
��׿u��i�8�ۿ�[�z P��d��9��z��h|x��(+�V�BQ�Й�0����#�ǋ�$�H&���3$����<��'Oo�}��W�����w/���/~�������W�O�<��߿���7�^��O����ݛ�/�?������9{�?>z������_<��^�Ã뽓��燧�u��ݷ���o�$���\�~{p�����><}��'�Ħ�o�X�Yl�jj��>��p|�i8��-�uT�.�D���־�ӤC.
'�(	�($˃�Y�����������4���_���x7�`V���C-=P���"�z᭱��]C���NˡSt�9h�1x�r�[d�@_�pN�鳺3ŇW4KM4�(�%eķ%�<��z�utl>��w��������4pȼ�d�/d��8���E���{�S] �\d:���hBF�׺J��-�4-_nۂ��ˆ�#�
i/&�ڝ�9��+G����Z?���J'e��ԏ��j��������ѴA���J!� ��dM�N)����m���������+��	�'�m��a�*0�dC�
�O!�`)���96��񞢷��]�c��X�P��7�HBN]�tv��X�!��Q���£u�q�4	�,�'!� ���GJ�3Y3�T�,┳���C
h45�*����M�]'�mƠ�����{�{ֿ�L}�ރ��{rl>#�Zߞ1<%i����/sz��k�����o�;�Ϟ<S�A����	T�_��W~��E.�W���+Vm7�+�8��@S�� ��:���RkB$��8X܆�>�J��V-#jϑ���Y�,A
l�4ӑ�qiE5Y?Ȣ��"G
Dh�L5`
D($%&|�U(&9�*��/�Om�����!��lx�W1������E��U�_2N�p�f�p�����g>�����&M�8����>�!,�P��@��)��\Y���)e�O60dS��ܲ�J焉�Ȑ�Q����� �=�D'h*bDKޙ�1"?��(��\>��X~`�D�d!�l����~`S���B��6X! �N
ũn���R����-D��Ά�.) ��$�Zb:9
��������G�)#�2�������E9B���Ѧ��D�A���N��$���5����#p�r��C:�x6ܔr�,"d��?|x��O3���`�brz��;�?GTK���@ִ��!3�f
,�c�7�f�k�� ��@�j�R����s!xR�%9���RTdEWO�)�BS�F�|��t�ұB�e�J�h��>��TX'e�B�!(=�����\.��IP"N�csd�'��H�B򧨬�V�B�i�YW"iFfǩ��kF"������K����bpF����n4?Z�*"��:�D5 ��7��{�!�R3H�Q��Ϳ��->�e<�KI��,d",��Q���ᘖ���h�*��s8N��D�P��8:�T���k����$����Vі6ʭ%>�!�)(��e�06���H��j�	�b�x��Q.���;�B����t74�+���uȦ9%"�F��a[�56}m�!咚=�\���&�I���@ȴ���#��X�pj��³����`:c�į.�)G"�%�/�8-�M?+_o�����g/����
9�F$˩-UwB��5S��P͔غ�C�45r�*�S#�t͛�[WaU��i`Z���)�ߨg�R ӿҦ�ض�(�(����c����d�@ʉ�.vtHᴜ��7�R��6�<�Ꮋ�>7�gu������Oy���g^O\�}�{�������������_������+��"�W��л�v����|}����}�O�&̾۬��ەZ��%�������.�R�+��;o���0L�a��E�gΞ��bٵ	뛗-�۟����]x��䛫�<7�J���Ͼ ċ��S/���O�?:{r�����{?#z�w<O￻z�Mͻ�c��.o|�՟A���M1M���*[�}x�ac�m���~vnm��smۇ���t\qVJ�x�����N�8+�8�;n�y��YK@)d;��¢���4�PE�D��6������1�`*W]H:l�8,�u���BN��ގ;H���r���'D��6�A3�`L��=(SYY8kԌ�����Y.���+4��(��q_��V�pH��844�Hq����P���(J�%���q�t�B��ϗ"�	i�r��v7O��hB�]B��2HIW15S�(�&��Ee�-Y�t���>�L�B��/8�aV]�Vv=���D�[��+��T��G�9[�2Fy�J���l��!�<�Ȳ�UǱ�N�N�d�H�k��p�;���ȇ���I��$�L7BY��ߟ�{ ��)��:ђӯ��ᎈ��~e�w�z�AB\u�.}�B��b��V�z�O���1|S������`�5�#����;������&)Y�����V{E�oHC�'�!��O�U@�pZ��Sg8�MS��%��{���R��s��۽=�N����0��<rwt|㍑ó㗯�?.�_<?����������n߿��g@Wg�Ϟ���O~���o��77{w�7>�櫫󏞟��}��������ý~w�����W߾�?z}�����]_�W�����S����]<;�9��3_��|�櫗��^h{��
��ځ9AE�%����I�c�}ة��H�j �N��P.��Dj9�"��ͧ$�qElc�XbU�_|��n�{�M�+�c�N����Ђ�"pt�C?�t�P������)�7��v�����	�#H7r�h�m�RW9�6�:K�I��(���[Z�ݔ�s9��Nl��OČq���=��l�Ǥ_�c���ɚ�`�Ԟ�!Eu⮏��S�c8��mQ
�1X"��ڱd7��KV�SE��I������&��vvy���CY����
���S��|⪴�[p!�����Kʉ<�*�fD3�äpD#��1��|
�
a㐊fZW���H�.����(T]�A��7��tҀ\�����g�Qn!�$��a`u[��N�,D-������|"u�J��p����4c:���BN�����:�+�b�%�FKPTT�Z`r�C(ۄ�����o����ꛯ�F����͞WJ��։�s~�[u\F�}ɌE{>8<Z�S�kw�����ۇCy�S��t������^�������:�_�}�ɧ��������~��]'8��׭�k��\�t�Bv�2=dH�'���OS�&�f[�#@�Y|S�� ����>D��( YHw�a{�@�ݖ�t��6��&� -@ҿ ��ퟹ�J�I�+�,SC.}�೦����LR4PzӤJ���C?���/d9|LV4qxuᤄ�V��p�h�t��K�,�(�����Z�h�8�B����z�U�U �[Q�J-餐iR����!6�,*�-Z]��AV!NYB8���o	4K���U!�i)��SV"3��RT7D�>m$;L}�`B83�`-s�mKE9��O��O�o�Mm��T��F�,����B���[�i�K�u۔����\}vŐK��a��h�ā�51 ���	�o,��S�_�-��+Tg�H���b�Z���P�#� �#�N8h@46��t��|���ìE��5ZoR�r�B�GVr�DS�f*�!��1䲥�t;p��F|<?���i�(Q�6}����R3B� '�4��
�F4��ZȜ֒T��[B�!K�l�-d*=S��|�XjJ���� 'U9~G�~vk������%Z,DE��,Y��|��h����"-BSQ�lu%j���,�Ȯ&�T�\I�V3�9����@��Q��S6�E����Кf�9=v(�)ݴ5V��8��X��>5�G�H;�o7d���
M2��C���RW,ڴW��%ֳܑZU�YpSNm�Ɯ�qRNdEB	��l��ɟ!nH��r���r١�g�Fեt���r�J��_n�l!Hx%�6C:r"�U)4�#5|G��9�>_�Әi�,R4��� p�"�Zd�aV�~�#�Jh��aq���?��mK��8�x������@ q��`���7~_�-�~�}��;oc3�-dBH}������
��Lb~��1�Z�ٹVe&�B���v��RHv����B��V'*����W��d��G����A�^K���#$R�Ղ,�M2���8�q8�Gu�D����MPY��	��F�N�"Dܔ�)]�.�LK�9M�h�1��PS��
_WSＤh��y`��Ĥ��H*'e��|":�| ?�/���g��	ʩ�(*�1�l�D ���u}Fѯx]ߞ��9����+��\�S�'�w�o�:�i�~q��a_]�|��Ɨ�������ˋ+�g�QI���.ʮ?!v�)����/|��p�#7O1�g-m�Wy��\����(_${�st��xoW~nf}���{���������G�~����w��u�&��L�M��t�cxvt���K_�tp}I�%o_#H������?�y��Dז��鳤(V�>F��H[�g�����(�pi��t�OGg���A{�@'�*�+W�D�� Ο�SY�	%n4��\F߈�)ה3~dS��e��?|#ed�t�r����12d��q�m'���7Ⱥñ�A��`�$�n��4��
d8��-l��t�q��pS�gLʌ�;�;�8E��]�� ��/N�)�V��r8����׭�=QE5SKZ͡� ���S����2�"З����VǱWF�L�U��,��г�	2`�&KB͈#QE4��.CY�t�^�.��(�,��4C��G�Gh�f�zM�'��7�"5���b�D�EA{m�Չ��U �!wJ��@�i{>���@Q~U�)N[�_�,��і�t��A� �.:y춳EoZ����"�MAd몖����e��q�3~�u> ե#_o	
1!'���g�p�R=��@����G}��_����Ѷ������э��'w����g���T��A�$Ř�𶒏�ld�|�z�0[Pb�v�T�IG�n�US�m�7�W���k��z][����|�����ɓo�۫��������W_~�������������x��/��λ�_>}r����ϻ��������ყ_������/�;>��|��z��ɫۛ��s?}}{�Ú��ο�G�>���Ol��=ԧ��ŚZ��u�oC���/���m�{N�b�'R�9�X�i�Lq�K�(�1�8��Q�i�tlt��;u�%��.� �c
��|L�8fu�TWι��ЊZoRJ[���IA� �S����C65d�j	��P�&�U��O��3�Y�q�s,_.<����O�4���̙iN����� i��F��_�a'*�pzdB�0�����e��>���D'��Rr��h�#�ZB��x����(�C�	i	��8�H4ҁ(����Z23�O- �
&P�6��+�4\c!@��W���ap�G]~���`�c�I
���+�'e$Ea�tĉ�HQ�(p�ԭ+����f*jd�`S�4�ۣUE�ҁV����j���Q�"��s{U�<���TݑBch�g8�z�A02 �2~c��+4���L���H���t��8���Bh%(8a�)����������*gt�J�D����NA�������Z��cOo�����ޙ�8G������pz�tv���Gz��e�x.��w��$�B紋L��[�F�$�׋���uL��[�>��mxۥ���c�=��H�����Ѫm��2ʥ)�H͈	�e��
���/���?�q�:YQ[��L"�2B���q~�̏b$%d$�^�E	�E �g�ZH�F��PR�d)�F��F�����%XK��V�1k2�����@E�?�_QQGhZ��)45�i]�Gi��V�  ��UȘ�0��M��|�)! s�G��VGԴC�P�F}�12U�r,�Q��eV"_�*�-m�Z�����'.d�wj��# =j�s>K�E�'�xY||x���)�$R`@�hFYǢ�"Ƙ�1��(�> ko�����*�f�u��GƱ��*
��Q6����Jԃc,Q��J�#T�D�@�{F�gqfD�%Y����7��Un)��R�M?Kh38��K�ޯqNcf���K��=����6�zh@dN�<��Ț���A�mH=��'�HS�}��sDe��� F�>;����<`n2���i�t���k�}r:b��(�i�����%S�`��&���`8Zj���Ĝ���R�����|�5�V�r%���G(���t�8p��G���Q��-k���C0��3�,Wc*����S�"�E�H��@m�'&n�4MY�,�+�8���@Z&���g�%�%OD.H�r�ĔcD` [Z���߈z2luX[�J�d�j�LVxH��;�C-�-���3Q~����N!H�m/�%O�BӜR"�dS���CR�D ��2�F_���Fk�R;m��7En�R�����8�Z��i8�L��X�@A��J��8��#T�8�1�2�!L"Ajv�C�Sn�Doh1�7}����5�V�Bā�[�x"�8F~j��jQc��d�i�'w�+��D�ț���A�Ԁ�,̪DHG�R��Լ�0�h���9PW�TT4�(j�l���>�Q!���u�_z�i�"��B�U�Tߛq�#�\�� $^KF)MqX�i	�L=Ec2S��q�Jlԏ\�M[�[����%��USj���/��swo�8��X�?�un�+�2���9W�WN��<�)�#�ǧ'N�+<|�[�g���?%��ݭ[�~�R��I�����F�|�w)9��K��N�3���bl'?>)���ָ޴�Ͱu��mG�3㓔>�O˸�q|t�O��:ۥ5�zxv~�p݉tP���ry�MJ?vv|�;Ǘ�_��3�~uӿ莟_�\��y���X�=WE?�iq�/����)Ⱦ]۩�i�T��\���ヵ雥���Y;�w+�t�_��ڷ���g��K�����rI1g�i��F朔�ɬ%��Oy���O�B�c~��e��P~�i=$�4EѴ�a���)
-Q	�u)����@WK0Ee�x=X�X)q���P�<��!6".�(�
X�V�D(��v�k2�8��Q�eO>Z�\�%�,��[Wnq2L=�Hq\��#�*�1wt�ڊ LWՒ��N3�)_h��R�O9��5��浡
2��V�[i/:�i
��� :=t���q�M"��5�V��uH�Q�-&Q��joS>YQ䍵�a/Ř��#7߈s�!�;|��-�ӱ:����z��8@�_�h))�)Q)d���g8���tL� 3�k��R���tz���Y
g9|��T+����~�/��'�|�κ����)���C�I�p�p���QȔ���O!�G�{܉b�:�uҷ�g<�����],�omZ!�����6��D�8:k��`���!�������)�*� >'���9;Y�����g\G~q��h��������ܕ�    IDAT���/On��=�9���ӏ/���w����݃O7G/����ʫ�?�y��W�����_��?/�����?~v�����>|�+�Yzvt���ݩd���?:zq����;?��ҙx�聻Uv�S�Vu�p2��0��C�6����8�=>�g���m�	�e7:�)��[-��n������q�)�`����ĭ+��r����UxGߧz1�Z]��ɜ���a�=	*j���w�Օ�@#���b�Q�Y
N��4���Rá�XQFJ��1##l�+=�}�R"4}�/D�Z��Tb'9e8����SN{SF�0
v�C�,#r�� ���s&ed���I�Cҳ��Ǭ�)���U���K�M�ᘐ6��)J*>�+z�R<�$��ӥ�SV�V�H��)T���\YSN��j)0qSf*4mC��Y
�D��#�r�#�8�B������oK1eA渧���tʢ!��_-�����ф�,$�f�h9@�iTٿ �t!��~0���>eN�i��HS9)B	J�!�2&C��!Ϫ� I�crHՏ3b���S��%����i��rݩu"�xV3�L��*R����� ����#:���+P���h-���o�Cλ�S��wH�ٿ:,ן����ӓ�o��}�7y��D��������_��_Z�Z�"I��ϙ��w��R�?,b��V�R���HP��=�[��#$׸���-}�����%��ѳ��mr8H���Pb4)@k\��m����)�!�6���|c�V�i[8�/˔N�\��B�%!��� ���G^���'�|j�.�{��	^�lR���H�k,YQ�N��7_T��%�d�֪��&�rBL�1���D���`QD��̩
�д�40A��0vZr�L��[!%�ZQ�M�4�LZS~����6�Z?4F'Da�r����,��$[
 ���Ԧm��,飉l
�$����QRj��R�?���Ң�)��j�h� �c�	�hL��b�^H�-�'%Y@Qdc�p�\h���&�I��DVj�D 2
��[>!��� M⛒26ժ����ۺ1��紺8F�P��i!��Oǁ;^ӧ�=��'�1jJ!~R=�DeiF�FuY̖� �BB!�Ie%5����/w���1����u>$ȏP�ҕ���Y!���+dD`��"?�����}��+u1����A�z�@N
1��hu!N�N�Y�8�|L�8Y��"~O��P�/Q
�ZJ���"9JT�g!"�ϚƔ�S�4e��ؔd8F���ir0���D��~4�|��r�2�`NnE�w�ݣ�2'2��ڊ��Ac���G��ۄ�8����
�A
�ޙXi�i������'�)$�C�7`|)��a6jM[r|:@�,>���L��)��Xbd���{�D�3�z�ie�@� |Y-��Jd���J ��0���C��SVʍQ�G���ж�Z�8B��1��?��Ѫ�0�|c�$�+}@��2SuE�qL�p8E5�Nv��)W3B�p�dEkr����?SՍȜ^͕h�$�.�ApJ�Y��P�\RUJ!q#��B�ʯ7��w|�C�,���g�:���7Ds�K�y�rq*A�o4Mm�ޟ �b�^�FH�)�xˆY!L]5�a�B���L��#o���6����r:�M�(�)�5��ˋW��ֆ[���`�_��^�v�s�ԛ�����j����}&��f�t/ӗ����s��'��;�V�wg���6	�?��ꓛG}��ŭ����3��<�u&����П�y�I̶b5�{?�vg{�D<M����=�pG�O]n?7�>X�+����ū��'@�I�2����Z�U��p|v�;9�����N��̍��x����Ot��y�+sUwwSu�uA�����o!u�q��mx�j�c���%E�Z\���k�4;j����+�s/s��e�b'��7u�� >��@L�6ů�4)�j��
���k M��Ti��B�J��
1R�tS��n���bQ@3m�=( �3L��)��7�u�Э����R�bN�`?U��!��j��	���]�~�iJ��2�5Od��-�,�Vd�T�4������,RH���H�4����q��&J$�t��R��VE���1�+Uj	��8���Efǘ�ݰ�
�U92Yײ�V�!�́0j�CM��e�K�r�P�Qm�ܔ&'�8��Ac�q�Y������?urT��W���j�ѷ�ȝQ��dQV:D"����f��ˀ��V�T�(D6����]L
35������a��u�L�r��8��}��A��Q� �����fP��;�d!p|
�D8����@Л]Bp2װ���2��@������?����JL����0�^	�V�� ����42�v��Ꜯck��	f@�B��Q�MK��ë�%[��n�3ҾR�׮{����9?�>�==���j�շ�v���7��͋_�:?yx�;�;y��w�����������ol�9ˋӋˇ�O>���_����W֋����s�G������Û�gO_~���_��>��O?vQ����3����;�aۢO�ju;i�gl��@L���C� te��p[��tG�8����L����MeQ0zփ0L
�B%*!���r��\����C���Oq_�9�t��2���1�'~��٣z�r��(>U��ili��g�) cּiN+�'&7G��!���6���7�����R0/1_(3��!��1R�����h�O�*h5O��������~��>���&��-�!�����2Չ��8�LVuƷ�qh��'�W���L�9Q�C�w��'��S��l�)E�q��&��r ��:�TE�[��d��rM7յ�9��o��)p$�c�9
EӏBДM�N�z�2�e����8��#T�����~***Tz�:��ЉV�oE�,0�i�э:WTE�3���H9��(�cJ�E9���Ie*�C�H�`�Q ��1S�Ki	���D�3]!��B� e�@��&�)Њ<�J�[ю��m��v�W]!��M-Sf�LW�������W�G���OGv��k�n�-�ݙ�Y�����֌���C�������O��O�)�߸����^Q]�34��B�4�#j�c�z�c6��	��l���!�(5�\��oT1M��|п���v�-%R{hJ��_����k4%ۈf�B2u�r���0�*B6;��#�,�U�*F��9D�u��B
�Ab�5��J$�L�S	u!MC�-�3���k����NS����_z�Fx�j�Q4K�a�e�1�� Z?q�Ԁ����MC��A��|� ���,�0߆;Oj�8�$X�@Ӝ$2䦥�9�k� ���|F!?�1rRC���(�ڍ|!�FJ
�
P��#�J=����YE��N�椆_�k�@f:�����ng_!��9�
W��L�1"{�4��.�"�	�?Q= ��io�Kǒ�"p�+�2|h�M�L)C�Zi)�B��,���-d�.k_3|?g
Ƒȩ�#ߊ���~M�,SbϨo�"g�Pc[�O��Ӧ�U9��m��WK�u>�)���j�%��pR���\F֢���-�y1�b�u�vf���1�
�T4DR?#�#T���$j��i�Ɖ̩PkT�cN'S�8�1��A3�ވ�֧P� �V8�e����j[�n��D�m#3U(?Ad�XS����P�ւb{�B��!DyJ �!U��I%[�BFaR Iq���δ��5S!�~0��2S��W��D|�(����@��Y2���"�Z�	�t��V"2��҅�^:��-�`� ��mu]����R9Q6:|�B�|
���'=�P��i�|	O��G`��8I��|#kj��L%�,��F��,J7v�q�����q�5�b�/���0���F�\�Q��\���i_��Q�H�ӳA�� ��2Uj�/�d鈖�r��TDH609Y`�i4�I�\�>{�ր\&j�ƪ��(�Z�oĄW1�T(����S������\�g So��	���~���������П��ć�FH���uQ�&�VJ�>�e
I
�=>�&�4 R����j�FU$.
LG-K��n���$2�Ȓ��D!���B6��!�u+���_�Ȕ���.��-��ɧ.�����G��n&��y|v�6����˻ۇG�D�}�vTǍF��<�9�&����C�W^7]z�����/wg��Gg>����k� �۪>����,�/|�n�Z��m��֭�މ�4�����#+��&ْo�.�L�����݋�3�.�wxv�~�s}���ט�>�y�˻�3�������x}4ͽˋ��nf^��];b�Vs�wi�oj�����G��m��m�l/bKߎ�}f����)G���KAȒM���	�,�O�s<dA�s��L�޶��e�7Nj�25�r�L	�k�[9c����%���s���o���@�d^�\F�C�Sn���Ӏ��IJ-�@�j���ǯ�X�Q
�ml��)+�B�G����Տ-��]�7��¥�<�(eH1)t�صS:�d�+�����ġ�	Y�(Ǖv>�&2_�!N�ؙ"+-=e��ʊJ�Ā���T�' Y�rռr8B�1�,"��� o��L�S�Dk��`�~�:䗥�����RLG�dYK�԰~R�Fʸ��`ZL�i��EM�>��`����t�dV�SV�4q:^�&b�s�*µjWYd85�H�QԞ8����O��ƪ �B*��B�NQ���;�5���	I�Li�t������s���αMr���Z@�R�P��V���;m�S�er��" 3����f.W:��s���g=�]�u��4a��=�+��b+��*�b�u�9���Sr9�q�')���G;;ݾ�Г�o`�7A^O,��k��==<��{_{�`}���=�x����'����o?�����o}�_�ʣ?=}�ɳ�w?�_��ɟ>�y������w^'��]�~����u�!x�O�]�޽��{����=��zqwv�Kk}�/R��/������`��=[��e�f`��ѶLH+�j��ιN���A�/��[2�h!�\j��!$Ĵ��W�\&�#���C
��-*�-�%#Y��>3QW��T�m
F����w���Կ��)��>5�Ǭۜ�y��'�NY���Tt��Ԍp�A�#��'2x! Bk�b���H�1M4&U���d#��5U�C֡lu5	��٢f]�!���jIor����t��c��iBu4!Cܿ���N��_��CAo�I���hJ��%�^�h"��f۫7 )Q�RڄE�q&�Ê�S-"9���0>N����i*^z#0C��F����;R�i�I��8+�)t�8��SR��(ڔ#j���K/�����E0%X9�
���@yNI�u&H�he��H1"����s��hE�l�(�*�d!�b�h �=���ӊ�p>0|�Q����3�FmPcpL�tk�,d]�O�X:m�>񍦺���,JM�=[�ӓ���OL:��٣?��Ǉ���\��/���#_>y�;��3��qo��A�j��/~៿^��$6j�-@_��/��n]`J/���i�#�R�b��o�l��m/�T�� B�ҁwDZ;q���!Z�)��O~��O�hÍ:Q����O�����U��i���!Κ��5 Jn�?�=��8)(�ϯ��ڋ ����,��8��{+���@!HcY��4�7L)��T��IE��
0�Չh��S��ɩD��U������'�_-�d�����miz+�đ��)*����uۘ~��@֔&���R!�)�I�%W�p�@6U��ְ\8Z��A�����J������41�$e4b�r�ˆLY��9�LqON���l����� ��S(�,N�t�w���MR�Q�iR�����ouF��nH�m�VVS>KP��FQ�a)Գ)r~��L\��/�l9<�A�wJ��HG�9�Ư��q���������K!.R�Fje���||`]��8D�S0!U!S�)�3�QV��L|J���Ù*8@����6�G3*m�*�پSW��L֘��d��T��f]�_K�c�[BR�.G-xǢ�F���3%"4&b�I�@��/Q�����V�O���J S6����҇G��ϒ�<Y@Sc-qX)�����!�P��'�N��#�)���oK>b?+�����4��#dZ�F���W�h��;H�RƤ�D�4ʪ�����AV�s�uu�2d�'4������pLS �VOP�ސ']h�S��D�*��D�����[/�\����H(�M�4��G�X�!ũ�
�L��.��c�!R"���]8�	�l�V�( @d1:r;{���g�B����8N ?5S�*�_�RR�+��C>�׳r�֘ B��qԉB3�đ��qIpīd��ƚ1�std1�P>e>�ihJ�8���i�Ϫ��q�\�`vO.DJ��2�װ�z���^(��V*�ĲRh��[K�B�pB�rtb������"�
BX��seq�ij�7b�4Y����J��
�O�U!F����l����Jԏ��)��mE��N.n�7�>[Kٹ?�Ǿ��tN�G&�.o����������)M7(u�������G-}������{ux篊}�����������N>��y�S�_?����Q���ߣu�9)pc�n;,G��ˈ��t��d��q��vxrtu�
�[6u}��v6Y�m��N�B٫/��u��>>�z�����<?zq�h>�׫�ǩ?m���ϛk_�{}�'iv���!^G٦�@n3�X��r�u.�lP��ѱ�8�m]�t�<G'5�ڣ�.����f��>������@w b:��b6Vn��y�$�lQ�D��ց�7L�1����%�
M�QA��G.k��L�&��S9+�tQ��2� 8i�w����4^?�U�]�r���qI��p��\��Z=�\���Z��Г+�	�bp�z�C´���r�!bZ�cBz�/�Bs�S�׌�BR�#PP�uՀ�,f�Ck�=oD�4��IA�@��RC��+�����d혺.�YEˑ���
!��p�r#+Ԫ�"����nykh*�����PSb�[����A��	2!���*���ic8J�Dm��ۍȃ��	�5ͯ2��P�S�	MV{+q�X���֡\����m��E�Qv�D�L��j�r�(�fu�$r��-�Tګ�G��V�=�ܩ�l���|���}N�W���/�Kuw?��O�#��nc��2�˚���^�#JHm����
C�u�!�5 :}Ն3��#N�Z�A���y�A;T�`�%�ӛ�v�ׇW~�{��?��gO~���/^]}��^<{�;}������y����/~���v_<9>����=~��k�>�����w�{���>xpz�V��?���o~���>��������;�?��?�ן���7~��t������n�%��i	�i�wt��^>����q_�-�X;)�eI��9�U�%ʢc�((�gȥ�`R��[�ҥP�ԉ�m{�\wg9�\v'�sh�����o&�t��NuM)t��L�*�C-�Th��C��!t"�����z����b�9�j��@
�j�&N9�t�h-MØ| �Ɗ���m��/J�B��7N�8�p�rM��ܴ�jU'��&�#r!#��ak�2�i�`ԉ�����-�r�� D�~j����w���)W%�ϴ��iV�S4�f�_
u�y����p;�7l�	�,�_o�����q�,c�'�h��Y�p���v�M���±��
�Br�H���2�r F�c��)%B)h��������Tj�)������@�'w�jS
M#�J7�e	B���.g���'c�[SO#r5f:��㼭[)V��Q%�#̱���2~�ZGK��,�� g�|
��F��a�Y��
�A����:ڨ�ݔ ��S�?��{����;�����׿�����P�=Q/�~����<gJ�嵕o�����h�b)�KF�N�)�L3��QK�C�UDNn*������Y�Ӡ��b��
�Q�H���P>N�H��.�M3A��N9��i�h�b��s�-�}���XZL�7p�Q��NN���~���myk�@�37�!O    IDAT���,J*~��VT��L��Dei�׃)\b�LY�~�^fm-�z�@�2���!#5����;
�}�E*t�d9^!u8��Rb	BD�Hn�k9
Gc
ʹ��e�'�G=�B=~ɒU�UW�X�'��\#�>�T7Y�-��J��,�N`S~G^n�����ٲ���J�A���������zj@�Qi��ɡL�3��8��r�C��$�Z��-y��^�����OM�����ޣO�ԈF�h�i��R�U~��Z�݋��=A���8����v��� �4bvN?�M�݆3SV�U�GYS�(��&�h�<HR�J�̙��g�Ĭ[��S��1*�r~��Naȝɦ��VT?�:G�W�_5О�5巺���a����ż���D)Գ\�Qƙ�Sj�JN.���[��R���#�9$��@|dF�#a��ѹ�|����lk��1]e��F"�z�/�og8���c9!��\-!���%�3S&7㷫��1�4���R�8ST(M������U�[BC��ycK.k:�P32YRLg�n�c�a9���9�¬�t�����f�M���**J���J���"�T(���B��8BE[0�����j�i����@�����g"dz ����x�m7�sL#�Q�
d�j;|��p2�Z�	l�z�	ep&�BS����H��Q�ғ���)g�>�pT�Z��Z�,.�S�X�r���7�)�D�X�B��<��z�'�B�)��1A+��?4H:3J�["ޣ��h�tj��H���hLH��C��P�)��=���y�W�Y������p!�pS8�(�#E'S+��ޒ-
���e��s�:�"F�s��P f����#�4N�r����K75ڄ��dp_�7��(�H$������CU��nk\���|����z����<������]��Vy�f��v��y}������)�N���כ����r |1�3�ϥ�5��������s�>v��7Þ���O�=���OX�����;�W7�z��ͣ�;Xw��n�;y_U{{�s?s�/����/<4|�t�����u�ԇ/}�탳����G��{���?������x]"����+��ђ��4�/}`�m����W>����l���=�[��K<s�K6�9�� ��rSNN]�8@
�h�eh4���NjU����	r}ߒї���D!j��t�@0Y�8	�����Q�P������9��Eea4]g�v�s'jXE�R���~L��]��E�eO8=1Em,r���T�|�K���LW<�UT�(��x������S9ׅ�c��Z�J;
�ZA���q�Y��0!jh�Mi���|M�3˂W��[��f�V�,SP�Qov���@ʢVa��D�*Z�,[$Z�(>��ф43j�S�B��[N)Դ�cJ�N��9�h�Ʊ�4�a�78#��gus�'ĸ��[�F"-�B�b�U�N�s�F��:]{�cK�d�h��FհǮ�qfɓ�)H��(�I�J@���PVm
�!C��r�q�1�@Hk�sL��*�Z��+��&�uW��2l�!LS72�}�뮘^J �wN�>��A��}LS@�6��x�X�4��,-ֱ)��8F�	i����Ɯ�t��C� ��ՂC:H�h>&��{��p��Z���YU������gO��Oj_���������������'�7�Y��\_���{�k�q��[Ǘ���_���~s����/��㚯..��;_y�}�����1ZkE�Z�������ӽ�8���^!���8`�V-��94Y��!����qD�p
i�IJi"1Ek)��Uȃ�m�v�����\Q'����v�H�[��(A��4 jjE�ΐJĩ����4#����!���953L�F{o�%6j Y�R�U��K/� �P�Q-'�p>��j@���\cQ�I�A�eeE�0�S!��G�Z@R�t0��ۇ���#4��0�D��'T��p��DL%Bd�;���r�3��J�q��k&�_J�kJ�f�8��%�BD��8��(�M�iM�!"�1JI֘����4��0N%��f`Q>�*��5�t�h�H'��%�m��@��U��W��!�h+B�&B��e���	z��JJK��EcR����L.M�D4S>>��c�p��4=Ɉ���1�gO���,�x�A)�c��h�d9����Q!K�6Sγ�,c"J�2E�����3k�(�sZ�4����L�/��/<Iz�a^\tԛjvۇ�UTK��ѽL���V��qzh�QpN-��%j������B�|#|_����5�a�@�Q��lBNbF�����++RZQ��h"p�e"M
�!�WZ	~��7"G����5&�ao8��iFKy�0Ui˪���I)F~��>��l�¡�I��%�d81���f��b"��u B*�����TȊ��b���pLⲒJ|�����@6Q�-0��.5x��1�i�O.KJ��jl�mB��r�<?}Sʵ�gp�'9?×����1���DR�i���z��Wn|!)�J�xl
�_����e�i+�<<�1���fip)E!�d��R����Sb)heխ)��@+J\�(Z)@��V%�|��8U��A�E�`��j�a��6�֥M��U= `V3eQ��e���8L �є�����gu.W�Vp ��&ؔOD
��D���m˄`ƩJ4Rn�̧�1�U'������#+��c�)#Ǭ�BM3h�nBpd�RXuk�U�\i��D�C���s*�rU&dKqG4�W�M!!��CB 
�sh�pz�A�r�6V�,���K)kZ���R�Y��M'B,} ����H�6�9��>����TO�3�$N4q�h�e!0H�|�JL�T�P|��d"	.�{4�9d%r��R
�(Jĳ���!N��������Li>N����)ӊ�pR
AJ��u��q�Z$�R�eT������*+&}N��8��]-Z�|S#N��h
����Y��U�ph��'?���4ߔ���>�Ј��J��p�P
V���,ԛ#���[Q�X��V}N�ȁ����E_�D�1qԪ�j�֏\��?'�T,�"1q�&���z��(\�t�3ٔ$��(�68�'hć��D'R�v�[��R�gyWR.K$ec� ��yuBz�e��fLdߡ0�ji��P3B�Q���ZVE	����H���?���{o����~j�	��7�V¨aS4&� ��-?�����C^|*ӿ��D���M�ϟ��zp�.��>5i鷾Z�ػG���G>�rx�l�~q�{G.��|=���*|y���i�\�.����ϳ���u��w�����uR�a_�$�5���U���vk�;o�ooֳ���Vs|x�[e-�2��۽������\�zp������^�]_����i{�v��ď�ܸ�L���;>�+5���k'�S�A_%��	e����� �"ӿ�lݮM`��4��B(�3��p8.;xD�I6�TQjBp>����Z���L����Q���.G�U��D�Ȋ�!�)Qn�ȌY��Օ6�΋I��ǵt�aR.�ݦ`���M��|#A;�f��#�\)EV7~�U�y� >�Q��Ҁ�u~��YK�ԏ'�֕k/����CcT��/ S��ѧf�[S#�!Y§c�`�9��R�*jϨ:>e�||�b��#�uKMc����9����������Kԧ6:��@Rƪ��!>��g�@0!U�d���Kb3���Ɏ/�_9Q�m,�q����4kZ�-�o׹�o�&M�)N�tb!)A�VTT3ՂpDS��R�KG��ZS&M:B\'�\�c��(���B!j�J�<}g4�u�i�E�رGZA��bTPm�X�;ljϨQ#��شfiQ;��AkT�j+j���{��~}�<��s�=�{� Đ4����;���"��ٟ����������dϾw�+u���_]������j�{�)٦�P5Ͷ�4"xWʠ_�ݐ�lX��xVԌV�&��T[i��p ]_f��9؟�04<3)ٓV;���ڞ\_x|u���3k ]o"�f��cȪ���߫�������a��}5ҷ߫���]H��Zjzq���w�2f�ق i>����+��8xM��b6��-Gg�g���]ߠ�<�J�Q�e�$�;;�{���|^�������V�GcA�%x�k� Q�G�H�*��
)���{u�XS_��;:�Z��{��g����4bfY��[�B��[�g&)�Б����Uݮ�1�Y��&Q�jr���QD�s��h{���K�����e_�פ���~Y��N����vL��^�K?�И�L 1 ��Q;����l���ށ�]�/B�&�I ��n�նgɝ��.�
�����(30*��؊�l�lv<�έ�t����Q^�~��#1�n�7aZ1�q������>�Ua�L���8� q��^'�0U����;kmG�n��{�O�_<�խ~�JU�7�G��\�l7	Z��x	Fƌ���3o�@]�U+�����x��N&� 3&��hX&�/��DgΆ(J^.�
�K�f� �!E���c_^��+7��]��N�����^lS�2I���D�9�.���5E~ޤ�������>g�k\k���y�Q
�h�{&
p��n��go��!V���d6����kjAYDы���ԁ��_A�e6�3
��#����ʌZGa�K��vK�+��<C�P�h��LT���i$I�@�]�P\%�i�E?z�����3�݌N0z�!g���N��bD�=/�*� �]c���DW&�1�>o_kY�cf\��������
䠄�aki�2���w�XC��-��.s<�A��u4�Y�_���×z�#j��g��я�w��μ�0�[h���EDj�|R�x�M��"*'���R���	�Yj5�)����&k�����-�\w�,"��{)F/��y��C�Y�]��.\׊_���4_�b�Xt:v��"��߀_[f�@��=Z��S�`��Y!�Z���:�w��F��mb�b��;ƞ2䊛@���s��{�n�&��^^ތ: m���Q!� �,��GB�ʁWZΗcĢ8��R�]���o��2'�h��4��2��H����R$��
��W�4zQ��"�-N����R&/�<�DEPM@7�ô�{yS3a����E��,kE��E���/�l�Tؽ<$�hK$�4�׋3��:f��N*ɾ�Eß���w�<V9�+ag���2��=e0ԇi4��Y�,���^Es6	��o(;%@�_��A�sieyT� � �'g8�!�A�2��Q�ժ��A߭#�Wg2��(�I� Y+�8]>�"N�lv�L4��ߌ��N�i���e���|O�B���c�P�����8�D}��+�J)���%��A��k>ê����%nN#��#.�V�(�hh��4�e�DzF;�uƥX�٭=g���.w�	�e;��FU\!��ay=JL���|^�G��/g,N�/R�Ꝺ��!�i�ؗ.NΔVI0��!��bO}�4��n�麙 ��U��he��QZl	?-����V�]�!Eַ�y�5m��������&�o�G��6O����������k-��{�ǫUO6��6J7��_�E6�5߫����"4g���ۻ�!!-w�:��\T�6U�\�<�k�:b��t{{��u��<�Y����k�����?S�tR�C̻����oT-��Too���=}�ߞ?c�mc�Pc��3(�û�w��L:=�BqtN6��w��l���D��K��H��c�:��(����'�~�PK�;]��	�-J����mLmh��մ���t���Z[�B�Z
h�'1� ��6N�s��o����녌/�
��{��Y�fB7.�:����{�,�c�A�83��a`���
���R-}4V-U�x൦q�!9*�G���'�K�E�S��U9�0���������5�9��N��E���P�	�]�|���m������9*��u�(�^Y��W�K��b�����O .�T;30��9��,0�_C�Mٹ�_=��Z"Zc�+fH.gqq'�!�ƚ�I�SƻTCq�]'8�ՇV�t�< s~A�]�g�7�9v��R�I�:�D�,�X�o��<��5�b	C.�8��%\�2�|�5[8�݅����M�j�â9^ejJ[����]A6o4�RU
}kbSTp�ǂ�@y�-��nJe�N��i�4'Z�Cs�Qt]�=�[Jj�{i3%�Y��������oa똍k,X�0b�I"jA,<?��`�V��Q�2Y	�@,��<o��}�*�\��q(9.����W����������Z��Tτo����g�cϞ2y?}�龜7���Z�i���Y�u�O�[�����O.��m�ۜTw[k���#�d����o���hJ��5��cK|�;��B�M��Nѵ�������7�+��}�*9���&�~��mx�8�A:Z���|�L�[+9
�̘6vcSS7./{!J!_���f��:�V�_��Hg>t����P)V���m�6�Ԑ������s��5��++jO��E&j����b�3>+W�
PO%�$�v�3_�&�C�p���wb�����о�9t��`M���e���a\I
�R'(�@+v�2���އ]i�fD�6�Qf�b��@��:U�T���zi�������Xe��u#=�}�=��!���B1����VDPUp�ϯ��оj��z�k�y��at�v,dBR�(,D��zں(4�.��rQ���2�~��5�\�%Am��$��䐜�zW�u[�E�/��'f
<�1'�v7�3��{�	�w�[����ի���>�pq�pu�H����"tZ)GE��Z#Gc���xb۝���u��"�	˘�l�:�\���rK�"������+-0�k�B���QHpV�����))p�;�Nh�D�@�h�t;�?I?�W���!�/2�w]�Z׾�74l(,h��5��fL�}���gϥ��s�$�m����9�2��e �+8��
	ps�,K����)cVEÏd�hȋ5��N��*R��V�8����,Y���^!��O�,�Ns3�Ъ�]/@��(�����ⴱWv�t�s����2�:�Vk[�[0r���-�����:P̠ש���̹��}{F�#�"F"��Ç�ǸP�R*��=����zJɲ�n>�2�y������=�*�4��O�9ʠ�^��n�O�G%3M�KU$}��<�����qӨ�x��pe��֦Ka�G�:?�%���jz�$PEw�q�yn�z�*���@����ز�#HSUx���T���WF�:�S}j�X.�����1n,u�E�'v��=zH�ks+U����	��:�m7��S�/�{����Dd,*+}	��[{o�e�� ����F�b���4�Q��w޽يI��T>zȶ�۵��� u)ڨm�>��SMG��Xz�o

�̒cb�cQf^Q���t[�.��ϗ0��Ǜ�6�D|*� ��=ц0�#3M�{�idI�긶y�i��6�`M��Z��M���u۶0�l"��[�t�:g�:gt��cL����GN�O�gG�5[�SwD�1�EM%�c�g�N��N����n�8�B�=���E/�ܭL������	 k�c�G�Ƭ���w{4~}W��p;?4�Y*��G�Ѳ�lN���z"G*�M%JNS��ʔ�^Ew[���V-d�ES������V�͠6J��Lk#�U�=��lʸݔ�/�~q+\p$�Sa��2�@OT���b�P)����p��Q
%6kw��GEwm�W��'	,��*)��3��r&��+-R��� +�v�Oj�:���7.;#�b�?3Ғ|R��%�`��}���Qd����	�}�)N#`mx9]��M+��Dz�d���zM����3�����/3��|�x��Q�߶�IHWU����}�:��p�:?v�����M����N�������Z��S��J�P���yo���+=����z�^�p`��b�=�U��%En9[}��r� Ҽ��zߢ8iK<na�db�����dA��a�=�������g�ӟ~_νRU��.��?-���@�����1Y'��FJ3*��䛴�dv/7�+��'eu�s�b�}q���g�1���N�P��I���+�݁���k�M_eUh�`��`㐕�������O`""��57���RE����ם(z�R��ݜW�ZSו�8J���A�����ʸ�{�#�)(I1����9�xa-��1�oú��|W=dz�^�YÐY�U� ���;�1<���0�(Ot	�	�C0������	t	�?3||����2mH<GF��Xͯ�֢ek�-�X��e����i�B>�b��������yO�KMՅId��.C��#���(��&�ZxS/[���m}/��[  c�4��xF����ZR�Y�3�R��h����}�x����ۋ�[(�AkϷ}]��؏88�q�&�Oܡ^��y@FM���������%%���n:�u���BqTe%ح��j�\Q�hSd�ܿ������u���῿O}��#�4�M͡�xɳ7�
�މ\����҇�݆�6��R~���f�8&�&��cB�3dp�e�w珏�'?}�
WX���R�~��k�N����f��Ϋ���W[;�=�#a�{�]f�O�	�Ħ���yβĆ�*.ȕ�+������ӛ��&䉢iO*����{ �7d/X���Z���-{h�t`{/��&@@l7��,M�K��T�\nG��J��k]|�l���7W�@�pa��Ȕ�c	0
�����YO��Gt�z���I���T�'$�@��}a�\Z��c->p�L^���#���R̸[�}�̅o�����	�f��J�Ӯhh�����%���~���B�]Q@\~�C���xCf>�}�fѵS|�vٚ�-� �h_�,�|\��������K:�a)h���+�����A��<u��JuOCX���{�@�7_�ov��5��rz.y�w�"i�Q�."���3�̣��E�ZOo�Ώ��=��.��e3��|�
�/�2b���4���Ĳ�<���E�4#�hcٲ���,K7<� �L�[�X��9��ک]�Dޭ~љ� � wn�(T�ã�v������.)c�����7o�_߃�����s��ij�KQ�Z@ǿ�C+3n��x��T��o�K� �V��JM��)�߽V���ǑL�o��[��;,<��3?�	_�q9e���\�Zߕ�5:ʖ��򸨖�e�<�>g��?�1�"שS͠s��X�^V����3�}�u|����"��et�U�?T�И�՟�=������GJ���^�@�|�&f݆�n%Xx�� ��va�ɲT"PCR�f��B�͇�;�b�d؝C��E�3�&OT��6بQ'��D!|��C[�	��Hh�}�7��k��RÔ]+eD��IS�ԍ	���h����ބk�k�c��ٹ!�G6F(q�����c!�r��\M�W��īJ��"�
,D�]��+�-�(���1�DX�{�;a�Ja7����|.�F�7.�IS�s=.�b����B��bu
��R�>�sG�_�ݰꨇ�q	�7k�1�(�'V�,F�9����oFCW���e�(}�+�|�.V�:T��Z�w��F��t)�}�߃e�K�$�&��w$�E{#�P��D�.�Ki�'����#���-�Ճ�,�)3��1eT�qu��8�~>�B!��D*�Ӛ�>�};��z��mCq�%W�d>���K��� �<.��+�Ԅ��(�%�H�N�\������CÚ3�8E�������c;~�o|���"�3����
�(	<ʺ>�Rk��{k�2\!�aҒ+�s�<�ș�]�N,Ghi&C��T`X�F�
D �	�:�h%GYl���q"�s�h>}j���0� �����/o���Ԅl=i@�Մ~�'k� u����0��9и�M:��b�y ����.g��0[2�Pn[�^>��#���0�}��J����&�/��/�QR4s��v"�c���5�ǩ�!�ND�|�����h$9 t�.�����(�uϥ���������H�<]��"0˖铘y9�t	n0�?_dL�S���� !�=!�o�4�J�9
�NQ�2�G�>
�f�vmBFjF
����!�1�1�A�y�P�� �/���e]'LI��y|�v�q�� i�O=��KXK�RA7�qp��,�M׸�����:Ci�&uJGo�6���]�Wo����>�x\�c�����Z*#N�!�PL�f��ͳ������5TR���u���$�����˯�����˱ӂ8�wg������8��w���\�~/k����;𣁎��˹H�cj�ҥ�p��w}C�3t� ���?����=�� � W���୼>�F�V����q�����V�<{������Kg�_��I��PH�B�uhs@��8�V�����������|C����t|?&OX�z:�~v�kr�oٺu�	�6��!���0��I� ����ص��!HޙK���z[��i��ej��y���(�#B�
\�2���XF�|�\���?�\B�A�*f�Y�{ǘ���v+�.H]5�(��o�����Q%^;�پ���n%�=�V��'eF�}���
E|5�!R6Hqj�k��������<Y�X��ہA+0�l�W���������)/w�a��}�Û��k��x�8:��Ӻ����l֟u�]�.h��UX��H�����Lݑ��ix
���=�4۱��f��-측�wF�DU�'&�c|.|ac�N�e���V� ��|��ʞtG�� J�9�~2B�u�>����mJn�m[�}�r6] ��7^��	9�����ͣK�/3W{F[H8N�F�I
F�P�^����k�d�<�
P��[?p���D[B l�/RrA(�D<L	G��PI�B���	>��sb��y��}u2�F�9���<�W���E�t��P�@y�VE����b�,�MC]%PBr8�e��Ŧ�X�5
��3r��gK������?��^���W��������-�v�	?��q�X�:�19��
?��۝��vvyu������=x3�����Ř�o�)��߃�} �ۻ�4(�NK�ƊGћ�@�׿߿!�����ֈ�q�"ˬS=�J�k�� 0��T�i�٩a���y���h~�-2�Ҏ=�߼VUE�,~���U;��I�ųXS����R�"O�]-����u%mR�B�,����	$e�^N�ɕKj↩�SX����5$����u�++�A�aF)��׭Xl��h8:��ڠj�'���t�P��G�p��ٖ��U����Z������s������M�CEn!����l̪y-��Q��/�����^p�-�<9�Y�q��W��x�0 O�ĺ�*@�ưjLJ��d���G��Ŧ{�"O|є�oo��H4�o&��숙�Kc���D��j:X)�:r+/3 ����Z9���olW�}z2EPj�ITy�!�#�oD-�XY�YC���b��^3ø@�����l�^�-ށ4�M~ݮBv����Ӗ��պ�f3�Za�YN��b�p��jVCS)��BnJB�f�<��>��^���[�A2)�>�1@�l�޳@�@2b��))6aU�*w+���S_���	*�/D�Jy�SN��ޅ���b��`��%�I��c4� 8��v9�!�L��D��S���iY*xuG�u8�s15�G��ΐ�2*�*;~�%�~�t�1��q��.Z�2+
h��=������5+ZZ�ePJ�p��[��-����V%jAu*+p;�xf�|�I�d�?DrTT���=�
��A������ CA~����|�������6�-u�e�T���c��)r�Ѹ	--X6�$�� ~xK!��mS���z���r��D��X��ŏ���f��l	㿏�_]'�w��&;�v'��ё^{���"�DI^�Ϸ��O��N� OPRvm�2�s�:v�疁���1Y��^��n�����4�
^Z� ʲ�rMi�E�5�a	\D�3ü�	O*��xh�\�JD���uU��y |��c3X��\��D�E�ޡa1²/*a@P�
��粡n&�tb�[��O#q�� ]}}%{km2c�ܭa5L�@^�Cs8�߻�ˠs�T2Vi�&>�՛�f���F�S�q�����!�\2"A7�H��H�f��ƭ�[Q�?���	�|q���L�UDd)L6e�gccP��dY�Y���Q��*ZV�D���
qʫ��;Ō�
�
�6�:�Y,)6M���1�5�0��dk��1.+�4I���hh�)�8�`%��ь��fr;i+M���f�_�&�ָ�ZYJ ����&f�i�t#˷��+W�tA�SR�g��sj��������`��A�����p�����|xG��L��C�	��2���/
�S =�:Gr�H0:mX�X�0ؓ� �P�q���?�5��ZA����s�^�iLܧ.v��1�z0*�����ܐ|Y�'NZ�J������Q#�l��6��H�ʥ�H��Q�A��<<~�e�ݺ��@}C#��>&��m9�Hs����N��+��cs"!u�l���V�i��Ƃ��~l����v�wz���U4�8-�c�|r�N���ß{���	k��0���,;&��Q�1����~��.��.�HG6Mj���ij�H��k��`���e�����=��܍����SraWȻ�M�a��_&����Q��߃0��/j|��|���"�|��v�Q�L�0(����տ��˞��g:o����o_l����+�����M�kÛ�b�I����u����p]�y�����dED��_�P��Ȫ���4 �Hi��_g�xQ��|�Z\�,.ݹ�^�����MYnL�y��4�~&����#+��'��ۖ�:�ueZ
CkEm��)�Z~r�{<��#U�D��
�s�<�%����MT�/��g������ɢ2M�[O)6B%C�y�2-�Dyl؋0�A2,����JEl�,���x��MJ��Q�:�������i.	<w`�c!Da���C�+��B6l�╀�x��bOI?e��
��@G
j��Mu?RG��Ogi`G�ݣ��^�$jn�ݤ������&|+;R��%�n��	�f�8b����$}��[�Y0i���ᳪӻϜ�	՛����9����lĦ��.j}E��Z�;��j�~���P��G�:i���fO=5j:�m��{y���T�Au�IvR�J\Z��A9uB�������Fd�l~�b�.�bk��Cɯ���E�B��M�γ>�t;�}�s'�N��^����r\��o��Z֦���eɒ	\�F�^��:���z�,l��M�^�4�l�mF�-��:y����.&K�X_u^(]�Q��kY�V;	_ߙ��7ϫ�~F�	�ܖ�̨�:��o�j�]�u��;5�T����<$cć��H�M�w����te�k
�(�S�d��ޚeM˶����t!J1o2����\>D�@\�~�d����V�`K��3I�F����Mʪ3����	�_4E��ůܴ�j�aH��&7I�8�H��誔E]��`p��N7G�?u"�lS%	S~N��� S��G���dC�R$���y���׸��BӸ�J����H��Ǆ$��&�}zRKlZ�#���������e-�Iÿ�ZՉ��hM���`�?1wF>+_X��i��ts���#��Vx	��y�S^d�zH��X;h�f��@��@�s�e���`M�D�V�'|��f\-�������PJ.h%&礖9����R�^���#?����K��.��'��y��i&��� '��a���	!H��6'���p�w#�͓���*
Z
_������;	���{ �/�(U��x|Vԝ�����1;c�aQ,ĉk��1���u����57��aPW�:��$1�G jc�����q�L�؀��Aߨ��ԍ)�~?�3��)��M����&�Q��lW�'�[Ƨ�}E&�bp����b&=`N�a����+�]+I�)8�Y�<���[P,�n{5B���j����z��Rk1�T<�h��%^L�}���;ϙ�eS���:���*Mѻ�z��冐� ��%T�F�Tُ���j~l_'*z�r��g��rqu�Ž̾1p����
�f��	�G�>��P�(������=�<�7�J�6s4�bb\�w�nz*<�J�+�Ӱ�Tb�|����Y�8����o��Gš�3��[O�I��qh��n�n���S�Y��)�a�W���5�X=% ��͘����o{��c#�o	���.�*u*��
>�F*g��E{��)�y���$���~\��B!�����͋Z��<�Xɇh���	9�XԦ&��G�����"����
\&�b��X�V���	�(*� ]����� C����|>�ϸn*:9-���6��}�!�'/x;ec��h�Y��cߣ��\������#��xŕ}Z�zM#U��#�nW�FuG�(���_� έ	��!>�[���܌��D��|���p[*��E�����ι��;�X�vв��V"��*�q�nH�WT<�')�2�
Vm;�;h��3�7��h��C��r��ն݄m̊����D	f�	���W����H0�L��v�U0ly���� 虑vD�oݟ��D[��=���PR�3MҤ��'��pg��f<��ą�DѨTщ@�Hja�c��Hw�B𴶖ow��3"C�u�q�{9��F��]��"��#A��8�S}wJ���*���7��Ocܥa�����^Ϧjpڔ�����%����9�w����ʲ�eiZ��4a�
L�0��,a7S�:`�7i�LV��G^{���|]�*���+	�Qݵ�0��*I���^>� ����%��{�G��"��{��Fr��e�=NtZ�8�SEp�Q��Cj	���m�3��<�;�^��K�EFòH�߲�����[a�/�����O6�
��C�v��t��}�r��^b�v<Na��ퟑ_���	`��E��H������ҫ[�i�����:r<��DZbpg�t�Nq�NWՐ�r��Ӟ�T��+iw��?w�dM꼏;�ɜ��B��n�{-��d��N�_̟n��y���)�Շ/ON�l9w��@g'cg]�;�,R�D^
��(X�J����AR%��U�ӻ��KA;�޵�ٍO�w�X����-�8��R�
S�mr�ނ��kz���N���O��V�5��ZG�@����b�Lg�z��b��S1޾g��Ϩ�;U�%�������u���bN�@��7�φc*4�I&�PK�r�1L	�>)zQ%��}�:��	�:`�Ju��P��E9bB�	T�k�¦OD� ����8�#�}]��&�~�7��@Q�7�Rӱ���J�b��J�Gt\.� � ��Z���x�D��:9[�4V���~ �R*�Ee�QOuZK�'�4���T������a'��R���Z���� D=�E[�n��#��Bt.W~�������1r3�.
<5��a�|L���}J6���|�'":?0ۂ�Zį��{(;�[;Ys��H�ng��s�u�6ή�Z:��|�AK;XLUYwh�}���I�h�ҴhG{�OfHVI� NX������	��t~�Mc�slq{T�_�����+�le���w��Y�3����}��1��dǻ��r��d�����~���L�A���H�\fM?h��>?8��U}��yuv7�ꙚHG��x���������[01��~3���^J�h�nTb���mfV�Z)���m���;�C��EN�;f��k�S_��A�)zݙ��G�J}�->&�C��t����
�X�bc1h
Z�qW�1���YYP/�X%2�t\ʞJ*.dN�<��<��d�T?�z"�.�.;�P��E�Q��<�ǉy�z�@���ɶ�	�UfI��?aF�sh]���4�b�j�^X�`w�=A���Na�ꖢ���L_�Sd���bL��i���"M��Q�O�8=�~���Ɩ�'pp��H� pףz�*�sBc�)�.�ev��21�����
�xϝ��ș�����8����B_�Q5����P�K�@�W���H���Y��sbE7}��\�|O���LWj�l[���k2��ɦ�R�~o4���A�?� ;���/y��hՆ4#*�tse�2�'5r���b�HP�d�ɨ��̟M�Pu�}�"@�K4�a�a���E;X�Xb���z���=e"���oS��������\��nn뉂�H\�:ݕ:�2/%�*�J߈,jV֦��Z���n�e��\����;���+I�,H�/L=�A�#V7�'P11���|��g�agfI<+�xn��
�
v�^����^�������F���5k�3�)	7������k�YA�&¿(ia	H����s�c��p3���*-Q.�o�I��Xi���3Y�lS�c��*��`M��N�w��T����9��O�ܗ{&����-̠�����~'�rB-:1�/���d^��6	�x��hy�I�}��#��߂��{"^���s+�f��(�3� .�8�)�fY	�%���1��R]dƷ���y�����|����H�d�F��P`�G�1�\]t����%��Csm ��nX�R�� ��ゖg_��%ou=2u(�'��I0�A�Q��@�1X4�1"<\:(C��Fa�����祉�y�B,�
�Y� jD4.G����l�Ĵ������%d�y>�ϊ�a�m�o����\a9!k~n��bњ]X��!��%�;�������Xx&j��9�1�1��l�|���DhT91X%>m�����5]{�dM��=�Y��Z�Ųb�)��=$����S~ O�7z2Ƣ�Y�������ʃC�����}�a�ڞf���
�"��ػ�t�b��8��Ќ�{K>G�0w��� ��{cO+���y��L�q%V��ը��a�s�F
��AU����WΈ���Z4�q4"l�D�fa��j�(��������ů�̲y���}�܇*�\7IΤ�I��T:^��C�uV�%���z���SX�%s���u���Ff�A�V��t�_T�~�dR3�\T|��{�Z�Y���7����x}l���hg_���9X�9���ps�ϰ�+�5��G$���#	�d1�|�14�up�[l��`��|MhP���l"�q�?uS��K������#���a����KRO�����]ht��k��xa�GU�[��tZ�]E��I?n��(*��
l���F��]�_��*l+O�n���0���NA���Ν�����΢��g��kLv�MF��������4�|����c
��-g�`�{7f�!�k[���7	m�?^`_�~p}���n{�6���x��I����g!G�/3�/���{w��xݲe�2�y�}g����o�[�>�[�S���aօ�ku���>�����_S���V�N��v�M �*C�ݱMK�4I�J�èT�5�;�=�n|�����X��]�h�9��B�����>�ňJ#l��ml�� ��]`~���~�<{T�6��0��b�AQէ�RDmє(��[���	�\����f��M:bTր$�G�,aaKK�O���˿��K�-��v�il ��o���= �|�}�#,	6-F��&�o~�eA\v��{Y@�n�9[�: qyZ��OՔ��k`.�����//�Y���|�sZ.\HcK� +\���:ld�%K[���𢞌� "B����#K9�Ňy��Ѿ|8��s\�{:�O�c��uM*7�QxE���G8�ʫ���G���o7(r����h��8�۫�w.EϬƤ-˻��~6����n{�cm�>��i���@���4^�q�~�X�'Ŧ5F�, �p���5�ekZ	�h~�P���W�N������a��U����U�!�܈ワ�[�"So탷�fU8�3oĊ���� �棛��/�m�͟^Q�)��sz�t+��|�DS����N�s�$��t�������9&��:P _�q�¿�)��BV�Ov>���g~{8\�����������5����������һn����;W��׌Di�Z��G�c��]���
�ҽ{M'�	[�3>Ϥ��w�&w�T���)�L�L��q]��b﹉��PAVg�Yψ�_M0u���I$���9��a�F�G*�"Z�#��=���1|�UEam��]��>�:�^a�GD�͸�|��j1b�a�*��F��'�����O 	���`o׬��M݃r�#Yl ������L�ؘ��m�;Q�����ct`Șy"%xX��(.>�QZ��q������(�@�\_ .��d�F(���.;���� �a78|��T�߳Ϲ��!̠,<Z�$����.t#�{�+2��id)ؚ!����t��	t�_��u[a��}�~mMɚ�3:!�ڀ�/=�붥,�5:{��o�v��&�O�TLP=X��zHW XC�+���Mڅe�>���LU�g��b�f�/��N��J�����(T�W)sP ��`X�n��Lxſ�u�p�^
'� ��+��?��a\C���ti�Ёrs�q�1��r��L�b���� q�'{��{����$ U06��_#���M�}����#�������nފhW��c�������ή��'uN���4B�-]ES�S7��ZA�h�s3�����q�,��p������ �"�9b��-��h1`*Uon���O`�f,DT#�w�G �Y�1p'Uع�t,����Kk�E��������T��V�K\"�;�?T�#���*�ѿȖ	�>�1�/�7��1�J��Jۇ��O��d�j#0^��Q��ye.��܋X�t8����gTC���*�)���#�zNa��YWU4�GZ���DQl����刎|
�k["�o�
T��U��a�]MRxu��T��K�-}*�ߐ9%C��\(*b�(��im���Ѹ�2��k�f�@Κ{��;��)S���[J�<_j���G�_�h��%�J1;��0�{���u��FY��!�	抑q�&�ǂ�,�^����t6S�Ld��R;)�������r╂��o��j�� n3��E��QCg�4V�ǹ�@��y.�n�cM����-�Ԥ��o2Dz/*��Do��V�#&*���o���d��bz���%(�d��y��f�	�1`)��̠Z0�E6�=n%"v��8������o�F:a?a�Se5�
F���p����ꖨ�������)��bq�Fޖ+"Y��.���q@�W�Ți�&�g@P���_�3��a��q=���[S���."�j'� �ID�h+z��@��V=��6z��9��v�0�O��1 ���NO�g+j�m~ ���a�.]ɁV���6�`½�D�]�:�(Q/�f/���4�JPt�w3��o<�ɩ��[^n��v\��A\���*��c�ẗ8��]����;�����g8�K^~a�$"�/��*����,~C����M~�+� /'���hw�b�3`� KOv➖��>'��ܙr o�Qӻ�{��3��lg�=��Xr)@��7���x��w�5������ZB��wO)���/p�0	o���qP�����~����҃p������U/���������T�l.�x6���ŏ��WwL�����ԕ��ﾓ��/,��ޛk6q�|���L�����a��BN�2�Jz���0�˳���:�?
��/�Z6�a~Aa��f�tnU��꼵�o�����lr���j�2e�g��^���������.7�7��C,C�L�>ǟ�R3,N���!�7غ�R���o�匽2b�����%���P�u<�1��qegzF��i���pԵ������NP��0Ͱh�NJ�����p�K�����������y����v$��'74؜�>�8�?%��!�Lߘzrz�L�ϸA���YE?UY'��@K�É����@�0%��QR�����f7vY��!O� 6@ɿB�#+%��w��=��{���3G�Il�@N����|��=���E��eU<�ҿ3S����
�&�K?G
��o���ŧV:� ��/��D����������m�1Vd��[f�6S�f��D��Z����ZBT >YNjȶ�&���?� ����C Q��#L
b*�mR<{h�x��ӱ)�a���1�g��Z�iC�#�F�d���/].�ڍ����>��{���6��o���%0�����>�����r�0u�k��޶�_���\2i���Z[K���"!�\=Y	_��Ye�2Y���,$�OAJU88�8��s`��P9$h:�hW�G�]�R��{�_��W�1���`/��}���� ���=��3[i	��[DAna�v�³v���i?�3Ć�Ud�-J���R�
�h�B|Y�j�Ŷ9~�S��Tq����_5�\K���G�.��6,��ڦ��p]�|����qH�)�I*$�DD9F֪���
�G�)}�N�L�q��3!��D��@3�h(�� ��1V4�����E���B�B�J��Q�G�'�rSº�q����{
F����u���9�'��jՀ��J���𕮷��g�����k�5��~8L
��PT!c���Ke��B���h����1C�ᗥ�8MK��3U�`��VG��9���^,[�\"U���6B���2ẅA�2t��t��^D�U��E͝�,�qp��Q]ݤ\�ե�f=���ڐ�Ez n���[��2ijD����*>�Z4c\�V���1�O�*�������yܺ���ɕ+ZK��iکB_jɂ��Iuk�)ڭRH���t�J@4f*^Ι(�NH�GE!U�+y{-��7!�~����7���j��D�N�jŧS:D'e�~yMD��j]|�c�B�?Ƙ�E���}���"P�럏�^�Xd�@Q��AnSHS���~!(�	�����g!)��fv��6�-��(D2ͷ�B���hIID�����TW��7N?R�)A!)��J�U�쭊>ea��@aH�H�Zƪ ei#Ӥ󐂺eՉ)��5N{�D-�8I�9�L���:'Y��?u�5�g+�
�4#d�GN��ժR-�lN�JBf3�G�"ڔ��$����1e��'�I,�>3'r4>�����X!���_�Da�h8F����!F�Vr�Z���!(�Q�B�3'�N��`������&�2�j�2�@�������pR��DYG�4BБX�p�j�n�(M���s���"����Xc��� S��jUQ8��
!��g>Z�D���1U�L"k:�R�LKG����g]�I�� �cd{ue*�7�g���	�I|kᷓB���ґ5���C,�r%��25b�V7�����JW�`-��$}��!�BYE�����s1����4��8��~��%NMJ�S�ǁO�i�?!��ț�j�O�-��r�:'EqDS�JWT	8#k��P�����Y�r��)7�lKE>Gé"��fZωK)ʉC��+�m�='<�}�t8�ĺ���)�3N�H�D	���h"vX��/'}�E)��i��Fj5�=��JD��f���o��O9��j'�*WKj�4�VdR��cg"J����ob+WN"_!�"M��+mf!|�a�"4
�Ek��W�T��|��,
F~m�+1VN����&�C�Æ��lISJ�NL�駌��oL�B>���)�À�/%��}K���F)�9DD�/��28BQ��x[�/���A`���r�;�M��`o��$4=�H���>�i���+|L��֙)�R�!B|�f�[4�P�Ji�7V}�]�_�" �E��j5ӱ�E�&!�!��R�|6�2˄㣵![���2P��h�vꞝ���?Z鳌>�yr|8��]^�\��������]�G'N�����Xj����rwzyz������1�}u��_�����'�7�G'�7NFC=}<v��YA��œ;/`>�y~������5�]M>?�?:;=�`��_�<��nw�Ka���k������o���J[�ӧ/��ݽ���o�<=���󝚿v�'��x��7�=���U?�]����o<:��~t|zv��t��A���{_���-����|�h�)Q�n���h�A&?D������D 12"8@ǚ�[���/�l���CLG�Br-�?��i�Sz�?������M�o��f��۽�����Dm�Z���j4��3s�h���f��XWW7��\;pL B�kTqѡy3\H���ԃ�z���JR:4.�����!޻L��K��%8Rz3�����V�8Z׸��%ȴg�(�`���)WF��]hzHA�h�/�M��a�,���%�r�צ������D�d�]]>Mj�!���,�#����S�unE4�K���C�������"B�F�Ȧ������|�+*:��,�L'ݞ��Ж���BBȡW(AG0|J�R��qZ�^ut�9z�I
��-O�&>�FQ�`�Ps B����t�IyT�w�Z�Dd{詼'bޤ�裏�r��Ŕ^?@6[�WTc'q����ѹ?��*�@"����?��>�x&�m�sW(���r�0'��Zf����Dӥ�������G^�of�$6J�Xg
(�h��C�u�:�yd�+�J�� u?��S������ϻ���n�l�I����}�+_��{����|G�R���/���2�n^��wϻ�Y�6�j�[�B6ZWJ �+�	�nՊJ��!"�q��Hw ������!��g�j�>�q����(K�E# �$(�ְY���+gQZ*ĨiF��}�s$�����N�6߈F��A�g��+�9[����\"0B!��u�rRƺ���U)*$=�����@|6�X&)k�{�j�������A��t�/N0�ܚ��t8>f4��k�L�r1�	�i����$�֪�����}��-G��C��dMYQN�v���m�?!����D"����&ί�+B`J8c34N|���PN�(J����5s
T��jF֐)�1�5�OR?��M�IDV�e��B|d!㡓fkq���<m�=5��ءt�S�b�χp����D�;�Q�%P���AHEQ��|��A=3d:B@��`
)'���t�^��+wV�^�5�����~Z,>G	��������я~�%��V��o��������$��U��h��F�b�g[�:�|�v)2_��^Y5`�מ�r:XvD4A3J���'(�!���1,S��GN4
��y�������J#7�A����z�Ӓi+�-r[*š���uˁKLӔ�'e�r>&C�4��FѦ֨Vd�6��oC09���!���,%B�F!f:��� E�LV�~�M�M�D��e��@�B�M��ҍ��i��-�:4�P�#3���L�Ln�ē�����?��]�I�)H��;�]M��qЌKt�m,�H�J3���֘N�z���PQ ��t���3<ڬ'�=:ΐ���b��r�ő�T��c�"%2��A��I�(Z�ړ���,�����8�NiR�����B�':��.p��O)"�r�kġg�%ұ|ʪG3��e]� �$�Vuʅr*�KۄH�s���C8t����=��CtR]N�B���X���8��R3&Һ�Rj�(�BdK�

@}r�
1�������L�2Y�K��J+Ԗ�3�5Ӕ�+��Z��� �@"M�ҁ��`6�oE�(ږ��W������:t�-�N-�i�4U��	<(�A��<��).�_bdS>Q~���C�B��F�t����M9Ρ_��Zo�*B��k���qT�CL�50�L�CY�R��Ij|��95�T��1[�h �~���%� ��J�ČB��_(�rM���i-����SW΢t4 Af4�U�gF�աh�cʏƧ�f!���}v�*a+�pG�Vn�j��B�3pR8p�����6*����__�H�M��!􉛆  �����1�?�R0��(�Չ�+�*�F4`~
�L�r��!ڂk0��"'��1f`~QY4�@c�5	��2��%bj�hRo��YNYS��#qSY9��� ��p���)��F�%7�H���fE	�C2�(!G�o9�:li�Z�Үr|��!��_�LWS"�ѥĒ2J��%�������L�9@�?=G6�ld��si����gs���8��O�ضT�h�<[;�    IDAT�1VQ#�pmX�ߚ�c��*FM?�d!�9L�J��̺D2!S)B�c=���I�ҵq�a�G�>�yzqzv}s��Q�׫�.��n}��_z\�;l��1xr~���uw��j��=9u�.���?�V�靿���~����zwz�k�N�<l��N_:�9��ַ�>\\��s}���7�Z����<֧;ϝQ�'�P���������>�כ�3�g>�������;�={t�q��ӫ�_|rwu������N?b^���}6��Ͽy��������3��=�����7]�=O�v�����.�T����҇/����*�2"s�E'C��B�w�A����t�O����\S�>h�>��Ip�����������:a��V��D�Ȣ98�8@%��B������WהÈ�Idz㓂��)�B3��#��74�R��hڕ�w�y���,@v����N��Յ ���b���6*�
�(�� �-�t"h��t��)%q��=�R; g��e��@,� SFǔ�*S#D����\E4��,5��@N{�Q�t��?�1RNH)B���R��D�egKM˥�S2��h�#� ��1�#�+ʉ#�o��p���i��%%W�F։a�	t��Ƕ�3)l܇W~���4��&��`!Aʶ��_�.s�N]���D��Q�C�d9��R�C�4��wD�Q��lB�F:���Bޤ��˧Y�%�g5�P
6J��8̹��*���ՒPc��Z{g��������)#�o%;�Ub�`�j��n�2�t���r�,�t�ŤϏl1�Ȥ�����0� ��=x�~���}����{ϱ����cLQd���?�s�q���w��]O�=��q!9����s_Z�s������kژ���w7��[�h��!2�S�Z��rZ�2[Nm�9R(��s��(�}�Sb��B�6�#���)K���IP��c�D Vd�^'�=�Pn!�=u���3U��`S��9|Q#�u!��X]S����ҍȢr��c̲�uh��U{��i���D�a�ܡ��}S��h<�ҁ��9R
��sPpHmen�D���P���V�1��K�O��(�)�=!�tH"8䩮m���8Т��X.)�/��
ZR@H������v��9��
��i@
|���:g��WX?���T`d"�߆F@�irЦUdVu�G��/�?ԏt�Ę���ȚJ7mtʩ"b��1¬'st�;���i�%/K���65�tf��k�n�.>M!H1r��D0Mi&�b� r�V�y��#�Z�n��9�N���F_T
_禥4�Rߥ�� �~"-�~}��-K��6�w`�N�-����S�� ժ��[{c4%���[���+!tȩ=�2�d����Ŗ��dMI�rG|��Y�P|U��h@)�t,����,�&)�P�)_�^����~p��M��g���j��V$
��s��Թ,&e�b���H�D
|!�:䳔9��ȱަ)�Tn����5�#1�1���r"ɖ[�h���8l��3�|:��!�¯b=�W�O��I��lL����c��A*$H!��(�t��>����2J�hN��I`�3P�z@j�i�5M�rq^*TcC 8����)=q�� �.P��ND�75�(>��K�)�n��mic�Ɩ_c3�S��ATB��(��r�,�(ę�%%ډ�Ǟ \���@�L.�0�%��Dp�U�ڃ��|x)��b�[��XN�@Q��
q��	�g�S3*�(Kl+Lۨ�;�P��č	&N!��C'��o�8�~8���O@L�tB-D��7�kX���#^3��Bu��~v���Y/4���#�y�6���u���	�2Q\TFLј�HE2fBp)�p��Ed�74�Ԍ�mڪ%��i�D���/Ŕө��O���r�2�A ��h��6Y�8�s��j@
��XA�)#ԭ1����#�Y�)2<�SK)��i�%��L:�Z5,�H��hB8�
5�S`�C�O�K����,f�ш�V-�.FN�#ة>����8��g�S-R�UD���жP:�[��95�36ˁ C�L"�n!`�qR.+f�%Va����0`=7�#ʁDS����b�Ig��)n�I
�~f`g�hG�4)#�V�-!���ʗ>���B�BJ	N�t0!F`=��DS��M'�\c��-N�)@j5��h����i ��K��a�Y8�B�m�#dʟ5�S�1�)2�T��5����P��:��`ʤ{��wUo]z�ϯQz6-Ө4|8��h!Y��)-�p�h��D5Ӷ�рhF�5mgzeT������]r/������z:%�]ϯ`�ޗ2�=1j�t��+ZW��k�h������V���}Ç#c&��X��z8|Zѹlk�l��<n��7�O���w��㔗�{	�9���uŜ�<�)���������7^={݇h���C�����G�[��z�̫�����w��#�9��4��7���즧�'���l�����Z��������*��w)��w�jԷ�nG�ܟ�]^x�����ke=
u���D�V�v}:�{���>����h��ݿx��������羠v-���?��+�V��^�Ho���RQ&,�	��f;?�[�d���=~��D:�RF.=��'t�{ ��3=�M9�F<�L�F3b�$�z��*~LS
�R�iR�*'ET��aNQ��\�)8'6Dbx�/��q�c�҈�:�.5F�TQo�r1bz�L�fpt[{V�'�&�0����t"U7���)dd�{C�&�|P��@���t4���B�I����#2�E��F�/Ũ\�8��j!1!M���Hd�h
�����K_ct�� ��CD]�E=�AfD(���ʮ[q��hMEsVx�k,���������B��n�pf$xH�,ǈC��*l��[��R8J�hO���ȔM%*ǷQn�N�)/Z?j���r�q|�R�Q�NȦF��8�V� ��(�S��F&���v�CVB*�2�h��*!ڙ����&����`ӌ޷,�G�g�y��?���'|o�����1��(_=�9���i��}`*_����׽��04�D�3S`"j	�!�RR+�h�A�
�����6T���y��/��/�������lkDvW�H��C��W���) �?Z{τ!�p���/K���K�{���,�ѪQ!��J��ڮ�B������#DS�N�L�,f�D�|����ӡ&� ��@�)�l��hs4@�#N�����±��GFQ�u�]�Y)�����t��u�h����:^cN[��2q�K�[�)�����Q�}��3�)�R"G����9i6"��S�4=d�J�-�*��(!ZFV��dQ(d���\@�tGa�qfEL�q�(MRL�%G���LKkr�g|L�����sH-0�`�8��F)e5�P��H�r��l�_~�(�2���㪺���M��4���B#�NH�*(���*!F�,F��m�����aь@"� �V�i0I��pʹ��p�S�SWk7�����#ļ��T:5m0M?���������aV��z�q�k�I�Vn/J�� ���T���@��)��W���F�S�^)I�R�-M�bm#��{\����7�{2�ƫ
�>� _u
n��9q���5��X�ۆX#�(Y�*�p�M�ȉҔ�C3�s��n����0՞��)�M���&M�4��O+��M�`��&n�N�B���Ѐ�Y���-S�tUc�b�4�*p��%�=o�֕�,L&�����,�YJ$X-#A)��A�)p����B`���VTVx��O%�ř�J��p=���q�h�2����H��+|`k䌬\L�V���d�45�G�G�@}~�z��i�0�B|8�x��jJ�(
,�$ǔ.��ZfS�B��M#�W�f+*I95�R���Z��V:�.�����&8c7�.�6�4eY��@�9�qd�8-g�@=��:Bp�6�b�ҡI���h�tLkÈt�)RQ:9��r����	��iE�h��|�Ʊ3�h��Z�����[�����>V��'�t��ڳ�L�KOM.NS!N�qH�qZ\
��m'_E�h:�`
ę=A&��('���%TT"ˇ'ޒ%����)�$^>Njr%�!M�@(E�]�~k���/]"8'D�|�dS����Ac���"ʊs h�1�F��8�E�N�4
4�g��P�\H�3�҉��A��rX�M%�Q�d)muj����FS�XQS8���^]Y�2~:��prE)DKj)nO�� �Pb~�4i�%"q�k N'��N;���J�Ǒ��d���d�;)�b�2��a��E�M��V�Z��i��Ҁ�j�neW�8Ei�e��Sې-��%ŴNRh70E;= �.�J�aJDHGȔa�؎XE�5�HM!#\�����>)4�7�Ⱝ�Z ��6֯��j#��FSmCp4`ZH'-��Rf	p>�8�S6~!L�*֫P�� �nn���V9��*�7m���b:e�s�I��\Z�D�L�U�T��aBM��K,"Ѫc�V�8�ژ]���hd)�'�@J����&�@ʫ�m�k� �?S@8�p�
A"P�s�od��4-�������CA.K�_���/�ʕ��ˣw�-DT9�1�2ֽ�cZ�@>�6\:_E�C�8B��q�n���C��Zz�j=�w�-�*Z��_���_="�Ng�/�u���=���']�����������h����d�ɧ7�wz�y}g��w�W7��_�)�ɣ&=�\�4�{o]%�lz��Nm�`Z�hs����vw�>�is|@��M���3�[�D������w��ԯu��vwv�q�ףW�;?{�ړ��'�_���{_�{�><z������}�׮/^���'�>T��W?���?~��]y��޲`�g��v\:
��wۼ����j�-��:���H�3��/�đ���B8��ѹG�����폩��+�W�S�F)�n᜵��%����hƺ�ԡi��8x�pm��2���6mՉD�k������.�ޔ�Í�]V���J���+U	S>Zׯ\RR(H�	����#{�� �����VUo��@��Kט��'�nzt�����{����6ŁDa�%R��$��dL�(	ql06O� ~;>�O�>������Iʵ���Zk�{w��vw+��\�W�ɽ9c�A�7�j����/|oXi����g4]V�
^m��@�y��e�A�+i�@�53 ���I1 P!|�NIL\$"��<�tl��(08�N���N�{z�Y��"��1�����ԫ�V��,R|�@�=X�Kь�+XJ��yl�Fj���qq��7�);`{DH�w��j;����M@�I|��|WmͺIշ�9��N�h�^A}y���!ā�Z7��������%�L�@�R�pjh��b[ै �N��Q#w�{�+�[��~TY���~�S=���;��j)�ӻ�q���mOK���L�,/LPK�h� k)˶�Ug-euj
__4Ȟ��L�Z*����������������b���fI95W�����Y�����Q��?��ClB"�&?�������Dr#��1�35�~�+�;̖�+����q�Ф��ӽ!b���&���ږ�s2� ��#%VH�&�R�D!S��롩!� �D��H��Il���]�6�T�5ݛJ-|��>�F���A�!Z�֗�SP�1�(���0"�%۰շ1��g�~Ol�����I�2�Z4�5/��2OaH�dGGLY���e:���=�RR8�_�n��._����@��l��m˭��U���М�P��8��8LjzIC�Kn�ƓB`�����*e�h���od��kل�J:�v�<D*I3N�@}N�%�\ ��f���YCƄX�<�rI�I�̉����5��Rb:^��L�IUNS ��`{�CH�ٳB�((�Є !̣L�gq�d�.��R�~kz)��eU���Xj�v�#UFrh@(P�W�ǦX���vڵ�E �4�j}kEӄ�g���H"ZKE(Pd@]��L�d�A`�ā�8��K�\R՚���j���2v�\Y�4z>�҉��hZ�W"k�dg H�Ӑ¡	QU/�>8�fj��@*l�<��IPl$M>�XSjdɖ��3\�;�IT5-o	~�!�c
4b���Z�G.K8�ɧVkY�8�
�PJ.Vl��R,D d3g%<��H��
j�N������wn�0<|��h�E ����qʹ=(�	�?)U���1p&P���13s���Eh#q��Y�y/pA]l0|uz�5'��x�Pk~o8�������٩FI�v��M9Y��b�,
p�����W{��IДx٦�jGM��cV�� qF�Rv��CLEJ�T���	"�\�JIY�pF�d�&��C��(`�m�<@��Aw| �vR5jpK�O6�Z1~�pMҕ�3�y,#�S�,gd���Rl/�Vy��CS;YAV�Fp"�>��[S�8��PU`}�1��Z�GS@����#"�+�g�`� hħ `�V��;���3M-�5���&�S��u�
:gٖuǱ�D\ �QRb��؉�Y%RcPn�,�`Z�8MFGXmY�}�&G��lUʁt����x�6b��Sk��v\�
�^sC�A +���NUR&�)$�s�\,�1���-J��Y�z��]��lH�5v�Ia�e��#N�`KR���FHn�a
�g��3Y�x<15�o�B6~NVU�ATբI�MyHU��wT�J!���Է�RS�x��/v6e�8��֪�C� ��)۱tژiV�n�z�V�w2�8)"hJD<�U��j�-���fP�����F��s����,ܲ*�� �w��Q2�T�NMG�r��@\���|�2�=^m�qjZ�@P�0����4-�Q8�m�!�;�ٔ�;}φ?˙����$���Ս\k��gu��A��u�A^���� }��W�V�z?~*[jz�Czbwtd���݂dy:RDf�
c�,��qX�@0!����J9��mE�����J|�򱅟�ti}鍍���i��G�;��������!�?�y�8�N�ˋ���/�O�nO�������~���\_�����<<��	��_�x{D�$���8��d�{��~�ҷLG�7�W����W~[����BO��>�\3��-�qѵ����S��?���j�_>���=�[��Yӓӻ�S��.��>�\�-�_<����w7��գo���7�xv~��#��v���w]|���g���qy�����,�D�j�@
Rj��9���#@�� đRإ�MD����^uI�d]e�Vy'�?v#U�����j�ut�V6���(��Tk���Q�61B��L�2$%L\@\��w�m�s���l����/ʽ���%k)����`�!<��&�B��a��;6D�ti*�I�8��F�,�v��.kfjd��3#�M6dA'&VE�y��E���������Vۘ�Q6<�H�&�f���:m�gmd�� �����sI,@�8�u����Z;�]G��D��(����=I���M�>�M�T�!�K�B"�@"mJLa�RS+����-$Ւ���U���:ڲ�۩�%�_��Q:j�j���C
l\�����W�(+��&0]x�N�fUË	��K��d���#V+i �k��	���#�d���W.�М��yÈ1�7���=o�[?�t/���;~��ɴ��9��u�'>4��K˔z`8DҚ15s�h{�6�-0"2��+o���0Y�p-��e
6�Ћ���#�b���;Y>)xjo��F��?�3�KV;�t?���fka_%���7</0��!���W�`�>��#����h�c��V#ҏ[*�5���B��rޥ@̃��[լ��{ ��Z�k׉�e��ua���`<>o�,~[��@�iw	Z�Eꢪ���7	�#2�,�{F#UR�[
�x.0y�b�����޴F������e�9�R�C�ZD��2`K��L�����+dƫJ܄�5�I*2+U���d�rL,�i%�6I>5LK�B}���e�'����3�    IDAT����A�8dL�h�$ kf&v�
��v��!��R
��B�^j�2��%(�0K%
1���&��4�.R_<
�c��J�p7"��h���b/����c��`] ��b�Ad���R#�6�Ę)��MaU{A�P��<s|�������š` 3g�����{]�m�k����;�ڹ�SE�רg]ô�nj�Y����@�HyD{�eɢ�1�M1j��E����p�(��;��!˴��ۂX@��r�j-yL�@��X�8'�ɦ֓VV	B�E�F����(q8�f�k,3)����p-�.R.o0�jA��	�.-)��sQ�,�
�i!��Z��lw�8UUҜb�DJ�K"J�-6�C�����b"C��=Y�,D��T\���h�8�U8�K���b#���Q��8ͦ-��fR����0�\n ���]8���Qtڣ���lB��N��:q�!PP�t�7���BK���#T.�,�)���% f)��Ԕ�.�ǩES�S#ղ-�j!�G
�|/�`�-�]U�@�^�p��*&��3W��TEJ�J
L���*"8b��fCF�C���БZ&�x�ā�$�N;1<r� Ǒe�j=�3��'�WU���l�u�uY���l4Ӂ#�.���U��,2�:�|S9d�l
�
�
n01DV�����+^9�� �o�a�qj1��x�F:�(��xRʖ�X�R��0;�z񌾬 ZOs���� P��a�D�.*�7� (f5h�RPañ#�&�c��Z�Y�c��k6���e��8&^e������6A|�����S_Wa��e8�*f1�����������A��M"@`�����xˮ��a�*T8�JP*�Z�|�ʓJ�wE�8��a�6_�QF�M���Y�Gk�����*�Ɛ��W��̼F�ӽ �SN0)�U�Vj�����THJ�zUU�g�M1q%1s'HY��be�I���9�l�8�o�/@|��t�`8B�9Ɛ�b%�q��W���#0ĵ�2P|.e��V���Pe�Ѵd@ن�ŉ�Z�vn�b�f;8g�A�F3L3�T�7ƴ������=#f�#��q���pjj0`û��U.����	�;���C�b��X���Xj�մ*#ի�)o���"TR*<e�i� ����u�1�Z��'e�~!�p4gn�1p���⮀Sh%]���$8㍈B�MI0Or�TY��ԺǐS�d{NM���e�RܞNI5�ZAq����I�Y����3An��U�����*-��>��i�?��F��^���;��OF�\яU�YM��4J^�>9>9�g,ﮎ���6�~(��r��X�����o��P���~��o5oN/�����S���p����Q��S�s�n}Ji`�C���mt���3��O��8��!a���M��:.ýz����>]�����OjN�r~����7�txuv��o�}���������C����������pk>��O�}���g�o���t�S���4����KgG��m�~;�u���h�gjIA��ێw�x�ym�؃BU�������C�m���S�]_Uc*��a�&�@9f_U�0J
	Q�z��{�o��Y6��d�R�6���e7�,�~�֝	��>�b�D�L�K	�	*�YM�[ztxK�X��r"�v3���"t&��r-t����w�!�,�ڗɽ{��J4�i#ޫю�
������@L:�l@��<e%	J��N�w��i	�D`p��5��	���!��~}Р#�ٴ�P�B{�;���������f@x�N�bA�_8V ,�4�8Zp�$��a�����Ů�Q�}l�Hm�*L Nctts�AGY>M|Gm�W�<eG��Ŭ���V#H�T	�\%��y:Z���PwU�8b)
&k8P��ٜ�͌�>2���o��땥Ӵ�Y"���p��_�H�1��o�r����~Fs}���I�0��MH��.�����ڏ�T{�u r���Y���B:��cVc��!�e��S�2[��#/$����߿���8�ϧڼC�|��W�W�8~��w}�6�m�8���yJ)Y[3'5�x;n�;�a,�2#�:^A�"�u� R�zZ�A��H�v��Q"�4BpDAR1M|�,c	���t�"��޽�(�5�axb6
8�80\l�-�r�8��<�	��ZV;d|)�����Աl[����0� �g8�J���� ю[���R�#��%�����r�!�'�.f�J�*h*f��R(�A �:�)��L6������m�����!l˯g���b�jmG��6)4��Fm����j4�e�e�R�!�&�f
�N��<�.b�|���R��4yHLˎZVl��"�b��H,@�T�`銘*�Ȳ8��t��)$�ϗMV�ӻ����xfS�� �NC t��r��N�ZV+6�'�^
5�q<��:�5�OYR�C%��u] 8�/�
1ь�9�qd`�:�M(�kY��"���c���ी
,�`�����4��r���Pܨ<)��	Z�*X.V�)?K�!ڡ�/�}�G
�Q�l��x�o�cq)��vJ�g6��tix���s�1���:�UL�I!�H5a)^��_j�\�{��Q�!8���������zծy �|��'�ӏ��ޜ�4r"{��`�8���Q�&Ô��[B��ۖ�L#�y�!A����~j|��p�&�fRR�z�~4A	�ٴ��*�h��`�J�K��I�ۚʶ�Ԥ�9�X�O#A�t�L�KQS΋eC����6@C� �����"��4��2\s<Eq��j�.FߒxYA�5��`��6�3�Q ���T'�j��[V5
�y�U�͌�K� �Q:#ސ���|�O�G�p�1���/ol�4�!��r_^G�T��&q�vʛD����y�Y��6A:I�&ewEm B%�Sm���Q��eUM�k��������iԖ�IP@GgR�,2��i�@nNK��G�	:��<`�M����'+�!|���|:
�m�N)���5�,�8�6�l�����҉�3YA��,�"
��S��'��9)�e�P��J�l�p��1�f ���&�� o�h*�!n3��}�'V�oS8�h�7���-#��jy��7OH�G� AL�.�gϐm<Z���K�x�{��0[k��^�J�
�YG�º�c
�Zj�c{��%k���1	
^�{��o������mj]/�6%[�Զ����k΋�x�!����fR�Z�Bă�	��4[���m��IA�Xd!��(�����+�x�I�.��e�BԨa0 )�v)�xj�l��%��V�#�W���U�-=nJ��ĲhL��@mִ.wA�*�p�X��%|ZX6mc_;q;�ѥo��%����2��N��8xC�pj<�@\!Dǔ!U	��V���S��f�lht�ڎ�w`
����?{� j;���4y
����>B�-�v*@��R,U���	I�����=�!3'S�i��B�!A���Q@�R����� ���Z?y|t���o��>?���{qz�ƻ��CO������ɹ��<<����������յ�d�oUz>k�.�gsWw�W/zS8�?����g���A����=ɕ�Ťt�����\W�����������'�t���O���mD�'��G�~<ӯ�]�y�����W4�A����9P��1�㫛�o��~�k�����/�_����+��~�w������/�����׾|�n���7>�}���ˣ��ѩ�j���M5��Z����-f�a
p~Y���8�N��m�ˑ���a��ëi�Roh{_כ�d���C0���`:J�ј�1�ZA�of4٤V�vC*L�h�4���
*l S���B�������nB�/� :@ſ�(D�EJ�AU/X7��k�R�Ǘu8�b%�Hp-��צ-�q�I N5�1�i
�e#�o{4�	�l��"��fk��h>#����v&�7$Z����j�8Rʥ0���W�xM�G3�e�H���GN
�a���^#ٯlRfB���;�i��!�ꟍ�d!��S3Oc4�����Y� �J
�e-�B�K10YA�Rm�6�g��b
���"�ƻ��:a�����%s����b�t��8��;^ֲR����zE�ES���1U�J���SK���u'H%n<�*}++�T%�c���v�]���7��.��꼝K���o�z��%B���O�֔n2�jHKP���;�����lIWU�8JL_m������8<{�H��Y&�@$N)x�DP��DVU �*`]�W��������5��'����/��MJ��������>�����*�p<��|�M�g`�&�ކ�qfh;8�q�c�!�dԪ2����e4岆��l"q� ��l�cZ)
ʩ��v8K%Ȫd�,���.7�G��.�@�2-�����獇)K"�׎g@�^�[f�B��%����I�� �Ǭ���&�#�rx�Ǉ#G��OPS�>�/ŇC:��jiVR�Y�4���C�q,�pJu]�����*3C�i�� ��4��^�d��1����d��o��::��R�/��ĳ��M��į��h�Z ����;qYj�(�![G�!��3Y4Y��xx
��AU-źPS��!5�,�(a�З�)UŖ#" *"���y�ƋӷM��<��T����dKG���O}]!K!Y1ZL1Y)K
b]|y�$.&��e�"	1/����[Ʃ55�b:��y�hb3�:�{%E�,&�T�x����6����B_���(�)D`���R^��*N�1�p�����We-������إ�w]�B���~��_ҋo*�;�G�7-\;牟�����(~_�c���5<��E���%65�#�V�r�BKq�(P��liȗ:&8):ͦ$?���袄o*�e�ũ��<�<�j��p�\���e�k�e1[۫i��$��8qE���űlK�pR�e~�$~���l"ui1�Y��CT)��#���Z��i�J�#8j��vj��� ��UYf)O��b)���!�-U�7qR+A _J�a:bYU�u�ӑM!�dȪ2K}1S����j���bY��"w�����4��j�++ŀ��b�*,AH��ԋ��%�^ZNGK�̂��Qd8i��W"u$Ί�X��ti��+W%Ƅ�U�ޏ7�����"�+i	�J���-�4I]pd#(D�i��&�1I�S9�L����U���ۉI��$B��:4_G|�5�f�R_�p^�������R��̴�����Hl�|:��#�d�>.n�%��Xf��蔅C-�8�|�lZH'�/fR�ǒ2d����J2�I���(F�O?Z1�^pH�U�;:�Z0H�?�ZYWIG�K��ŒM6N}�R�UY��U�+���vD��Qh_<NF3�����Z�y�,�*��NWPm�8p{iw��)@�\	�Z� �&0���6l�!�.�'Q[U�Ml��S�g*A���*L��� �t��'[U�[vL��&����c4LH���c�)H��Lj?��^�,Y4��,{��u4y��
5��.�+o��]��E�B�P� ī�V!� �B�8-gw���0Y;�l���j�����wh7p�X��iJ哢 ����%�����e.eB"��,5>�t� � 3c*Ls_U/�v�SG~z	�4$>�h!��U�,~�*Mée�@� (�d���uq'[�) �3H;�"�DڻYֵ��N�8�DĬa eS�H�7�W�@�-Ow�h��/eG���Ŀ��鸋d�A�@�h U���L(h�:2
j!^����i~4_O���]�K���g�
����0��Qo���/�������~������<9�{����<8>��������O��.�Q���kz��u^;�9�v���/��_�\?L�����*�n^�ܿrv��͛��C�'�����	�88�!�8�ׇG'�~�ү�������"'��'�G�����W�w��!^�^}���ͯ���7�%ruz��������O~�Ga>�6���嗿�ç���k����Ƿ���~{�?O�?������;�кs�im�[:X���l���8Vo�v���-�*��ϻ1zt{��C��.�85�b"������ �U�^R�)$��</%� k�pq֨bC�gŖ���Z��4�81���9�B(�{ux�ɛH>�uD�K�;��_mw�o�5�f84ٜ��v0	B��ہ�[:(/:&�GS�lM��{C����(�ё9�^�J����Y-)���x���`�����ͣ���h�*�L�(���eUL���t�9mSGR��I*�ե�H5*}|��I�9���,�~f�֕��HS9@�Ȧ�MM���%�	��Q-e�@�ً%�
�Cx�)�g�-eIa��k��\�lѐ�T^��(ߛ7�|��6��҉UE�!U!�`���.(��.�*���d��#T�֗��"Ҩ4]��A���Q��u���m1ܨU��б� ��Bw]M����]d������&�� ���%%P��>��C4o����[�|�{�;qK!�av�%l�����:�Ę�
ڮ�B&��A��<5%fH�QC Z
x�<�R6k���Ka�F��Oy���w"^���o��O��O��G�����h��Ц�ӷ��2��ׅ2�/px;U»Z� �9��#L�͉#�i��Y��;��}܈c��Y�h��CpP��=��*19C�e*� �� 8�~�����fY�M�9|A-��7�*]R"@ A8/F0������t�b�,��ɒ2�@a��C*�PɈ��)���z|
�Wz����h�<VS���\�+�IG@�y�[
XL)15&Fx��t��R�2�X�]`��-�X����(0Y�+ix%:Z�R�٦\�8M/@�%dqj��Ë]Ix��T�M.%�e##��b�uAce��w��Ӽ,�-T.�kM���i�p1�g���ʦ��\冔o�u8h̒��AidYd�K����Iz����j�)�5������W� ����ղ�7]\tY",2�T5}�閈��F#��e�BY�.�j��"���&Ճ�Z1�9��&P.�?F��Hd�^y_Gkݥ�/��O_#�ֱh��B:b�~���Ѵd��FV(���� �0�r���K���.�x9�7�F�Jگ�*����
������b���k�� ��9k�dd��DV�8�xjug8�׋r)x�p��S�f�gd�Py�� ;�����	l\-Z-mDV�`�ę}I9F^\9��p�oǂ_)L����X�]�AF�*�u��QEs
#+ҷ�h��)L��7g.����p	�q�g�Z��p1Ϩ�i�?j8���솗R�0�f@P�R`)��,ծ��v����*J6s��,Y1�lJI��R��^�=���x�2m��3G��c<K:�z!0���:�SF󖲪4
fx[���	�̓���u��*��)��ŴN�F<Zw�C�9���4!3�� �t&pť,Y���^���;@)��x�H�i��)G��٣i	V�OVv��'�T�HxM�Fx�ؗ���UUwR�0L�T�F��1��y]pjZ�v�� g3|1o����(��bM�u�qtA 6d{��*O<N��yR��d4�T�RF�(d�3'ВiǪ�G|�L�Ϊ�Z+�d֮!8|R�F���l�!�6:b�r%puݾ�t����:áB_��/o)�ә��L;`SMP��Q�(�C�A��r1���� 
F���g���Z����B����|��FCP�{�x�P�������P@������έ�3����Hi$ �.��;%d�
��t
mM9�f:U��K}�o#!Rs��<����%r' h��R�J�>����ҁCxF�],)X����G` �v�ę�V
���8Ē	*(lw��'?��:F.���9#!��pҬ��B��%�3ȴ��Xn��D#�cG��iGh��/��H[�z=Zv��`�j��,�2&��y�p4�@J,�7'�0����d��ӿ�����ᤀ��*��BpX�_���0�}�}    IDATQ��)��X��^-�R���?⚡��-��f+a�!���x4�F�L��������⤿�7���2qK���\�m��b�ok���D��	��w6ׇ�~,������������/�e�����kO�_;��m���W篞}�_�����?���z<������'�/�����7��ۣ�?�������~ ����z��}���7��<�]�{�xw7��[ϲ�!usvrqt�nٯ��Σ���2��|����=;���W���׎�_�>��!��������+���q�����������g��w���޽�?O?�<�=����O(�!n���v�:I�@',�w5�U,�א8�u[�����m��^j+��qJ��I��BM�>��MA���oL�}������!1�J��,�$���ydRk��I�����f}x��$޿���#�[(����N�ƽL��;v�DHy���FRժS�Xy�˚S#�V
��lCv}�qCG!��I�y3�4C+W�&k��<S�fl��Z��Dadeq夐e�CT1|~/R� �� V�f�/HV`/��hę (@�]��! y�*l�.�]Pfj�4�CHA�	H�	��k�[�+~`�K�Z1KO��Td�	lGSF���S��sP�G��ص[AU��vvL��q�q�c�.�%��]�N�.���0|8�]
W"�R��#� ���'�~g�W&SX%f��f����}|�z�� �Z���|��>=%�oNY|��-��o�;��A�����dm��YN�S�M�L'�����h������Mֱڃ����+�c�vAx	I�6bVH�R�im<$k����6o;����?��?|v��������;�k� ��j��jeIi�e15[���1U1�4�o�0]���l��Ց���n��[��u�XWdƨ�a�����BJy��T�ɪB�
�<�0)���{��ik���R�>�0�i�
I����Z��, "�	0;Ld1.�f)6CK�A-Y%�x4q��5� R	M[����
�#>0�(�R8��q�R]��M�K(.Ҧow&&쪵/�iݜ����խ,Dw`�P��qJ5!2} !M".���Dfk
�L�D4e���R��mm���"��	�b�R4����U��.��<A��!�`u�͖6%k���T}�L̒���	#�J\��*��e��ow�R�,���e���4��s�p�|��ҿ��A�?�6�=��Ⱦ�!�=��zj)w�v���I"�U��C�&:�=�;%M"��!�̕X����S�chRju�Y#�8��F|WM�C����W.cۋ�٦l��y�M��a4u>U��h�U6@)|1)"L�%P\�ow2�R���/�/6$CT�̤x�+H͐pK]d�Rу��#OPl˺@�ܒ�B5Ѕ`ΰ_� �(t�{g�T��F<�eL3�� 3	qʃ[��@�<)L|�b��g���Cj�VmL�s'.��(�4yÈ�9}�-��gڶS�R
&Z��ۜ��)�O\�*}���C(XV"N3�ҙi�Cd!R�6�өҭ�QhL�
�,�ۋXU��H���,��U"�P�Zd)�.j�LVw�Y6@>��(۴RB�]4���b��h�Y�/�Z�LH1`je)�G х�Lz������1�.��!q�~/�u�R
�4�,���Ze���Y
� �pjOS��+�<|3 ��0Ӂ�fX��_"��e
�Yꮋ���l�^�bH[�V
R:��	�#�'�&�jѾ�3� �p�l%���N��đ�Kjh��8�3�g�Y������<	΃-�M%X-D�r:������S��Q��I��X6����S �����j#��^
n���೑f �)f8l�z� ��3\kK�� f@�� �XH��ߺ�Tk)��ġ̶��u)��̀�,n������ �,�#F������BK1�WG)�,~�`����0����8�h��:^Ab�N��˪w�u�E��p����01C�/��D^�n��ǯ ܉���r��v�,� _,���0�Ym���D��p*ɀ4cB��LJ#AݛaK>^ҁ҉�OA,���N���V����!]�=��^8��&k��?q&<�r�y�@���TK��J%��āJK�q0��<V)1�� �eY�ڍ`R��tԺO���V�[fM%���j�����û�T�(馒B���C��%���[Ư{���fi<&��-��i����:f
J�%����ה9K�a*/��ҿn�O��Q�{ãY�ji�b�F���R`S���x|�Ӳ�UGP����zi���Wm��[L���g�ĵ�#�g��:[�#'BP�`����e�t��V!2BY� �#���K)1�����n1�t���o�=_o����ݞ������>��������yM��7����������p�Tc}��?9;���A����mO]3n�G�~f��n���8�w��w���?��{ì۸mb8��L�C�G�����
�؟�\�G��}�;��*���&�/>$��o���_9<9?>{�����g�~����/?��׏����'g~�������������=|��~��֏���Tw{���VĻ�] '�r����k���;m�!c�R�i��4���6��e][߮][�7� !��O��T-+��g�GhA�;MU�KYR�	�d�lYJ�3U4ËǛ�[���w��{�=�.���tWզ��fG�Re{� +�����������ѻ1q��ON�.M���*�!�?=��(��N�^4�T}������m��
�"�� �7 �ݑ�Tew�4q�M�6�'k4����*�� �D1�%FЎ,�:��v���<v���(��q]����>��~#)Y%m�=*d�y�� ��U�D��GD!2A�����-W2<B`�a�&f�|_�0�4�d_jDֹ��;or���"����yT���~��m�"��Üp
z��.�u{��Q} ���~�O��Oܽp��,v�պu�MJ��T�?4�^��q�ִ��?u�r���L����{i@d����k~?-\V�����ۿ}뭷:/lrN�)�Cc��;OV,E�ɨ7+�����W�B4����5<�4�C&aZ^��&��e�����������Kb����q:�����v���aML�%[_��hZ؝r)j�mZ����7F�@�*�*D��&dp"8vA_V�kT�8�ɉ���RE��@,��t��v���b"X2�<�r�N���]k���Yc����`��lB1SBV�Y!#������M�	d!�1���jS�Yvz�MYb�D0���]��Y�9y%
����e><}qFB��`��D���M,`�ϛd��J�0H3�!ȕ7�SB�=D��	��<,���ܲ�SkB8)��%%���+èM�/�3L%h��B�TR�E�b!���hԊJ���l]v� "+l�)GD�Y��b:�<K
8��UiǙ�
�y
-㣵kA��5AGWʄ��G�x���0�,O ���{��=�p|���ײ�6Y �׸'��W��8�N�G���&�����X,�W'f��h&a�U`LU:b�aNR���6��(N��'"0�rdY�l��?��/{=e�4}pP6�	�NJk1O���.8�����H!�N̒l�ZX
���Q�cG��?�p�侜�^I�B�xS�˒)�_��e]��7�8	��؃=>�R�&KD������X���քD�DS�~8#)�����ɠ)�32�~;j�u�,�Y�gp�=a8��Fm�
!�R!�7߄q�i�B�u��G�JUE�w�0M d���$!��@�7Kq�6b�4u��sv�t�|��Rk�m ��g4�(�m�kђ�t�52C:�K^��U�!(���Kz�U���LJ-p����jc+����'g�E!)x����äc��(�wqO�.�c�&&B���D���2[�T!R�%�☫�6)��Uw~�)@V�C��)__>/��<�!���?�Z�/Ԍ�x��! w{@�����$�i�R���m��Z×�S e�G�@k1��N�+�lY�IB�!�%"���j�$n��F��Gf�  �i*��crK�2�
S���iZƱD@!傭n�W����M��P�j����Q����!���#~~�h�lR��D�Y�C�
����>�>Bʕ�d�b�W,�u��VSA��H-�\�]�UA �J,�߃@�g^/�gf�dfN
��
.&¤�f��Ѩ�NVj��
���C�`1���%�	��\)��I��ر���e�f(6���ٸ�C
.l;`�+o)�Kx��*��ɛ��8���������d߄�M�̘��:�M<�8�a�Kwۅl���\	B�������Z3�bA����F��~�p̦0��F�W��eUŚ*5e��+�o��R4��A�v��|�uG�0Y|4V!�8�eg�j����ͣyz�jڨ,GߒY�3��d�1� ��AJ`��V��G0��Y)���Ȧ��e[�]�6?/f�^��)�]c�ʻU��85��B������Rv�k��~��S�l�lִ3a�IA�d;x1��e�����bK�fˆ�i��i��B�;��
��AUW!�����ȒJ_���lG���X�ұ3~���t�g���O/���}�p|~����;�>���;8�;[?��w�Rp������G�{�w�^����<q{t�>�<{r��5��;�9�a����/n}2yx��ʦ��y|r|p��#A���c�>Fuͷ���۽��|qy�W���������<y~s{v�}+����Gʞ^\]{t�=�8?<���;Z˞}������}���/��^�ϖ�ˠ�U�7x��_����g�~�ԗ�+o�����[ݮ�sE��$-]�+��.N�g�x�M/������=�<�KF܍m)�g8�#���/hbV���Y�)Y�4M+�˲6a�pA`�BRZ ��6�,D�<�%_���^S|Aw���z��w�]9��`w�*�>�<��rip:=�6�!
�*��(�2��T���u(�%K�7�eG�c��|�6��]�S��Wd�?T{̲i)($����b b_J�:�o��,e���?�7A�N�� ��B7	O���,
6ei�����5<��i��Yܜ=i���AW���Wh�޹bp`��tU� �pc4�e�"�V#�&ćF6�%�P�_N����WlS�N��+�;.�tX�L1KA��83o��/Mq��,\��A��rڹ����v�]����.�ݴN^�K㾅Hy�ԴJ�����o���[oIu2<�<M�S���0���pĐb|�z��xR8	*�koM�-��i6K1}|�-�:%b`ȉ�̊�'B(�I���Wo��bY��� ����cd�� ߒ�����Rb^
��Ҍ/UI�4Fo8�S
�y<5����Ë������_��'�d���^9e�*;���&�L�Gߙ
���x��8���ʺ�h�^&)@`-uG�o �L�b��9uq	}��n��Q"��"�`<U݅�#�Q�oK�Jq7�����܆�4�G�{�A᣹�5U�����!�ķͭ+�SG:K48DʴME�����FΓ%�G�%5��]4XG
�l��8t)�ťR�&�%��4-�Ɖ���g���P�6����TI���J���;X)q��;R�p��:���*�tiB|����ܝS_K��*��ަܜ�F*5���)T[�.j��A#.�&Pć�+�1Rօ�Rd5�Ӏ�3�Ԫ���<��R�!̓���YG13��&(.+VK��I�F����C�/ ..�����G�B�1�Z�%��'�}���C�	I�($�J#�U���E�����k��*�e�LsIES�0-|Wj/@4�bU=�|�B� �!��Y����H�G�k
�
fP���3�%PG��-M1�x�2�u@��|g88q��)PS]�<>e�v>�'p"M"�m6:�-�ӠcI�UC3�X T+k�d����b� �Xz9C��q�ٮ�kmY_��	��4�4�D�R�b��d3�Rc[h�ł�+�'�W�.1IY������ �d�Q"��/��$E�R<��Äk�f�#Raj�z�#Pp��f)��L��IA������Z12&�h�r>�+N�,�! �w�HQ���Kf���μX!MH|%i��̋��%�nTK��6�����>ô,k���;����Jb�E�10�H+L����!���&� �!�L�J��k�$��/"�#���JA���܀x&���ݱ���R��F&[*~�j���p4Us��:j�Y�v���hi�&;�(K��&��0�bZ�b��ojM�)�mNa[���̽�)D����b	ʶ��'��.b�d#g���jT�Wb��������Ȗ�UL�2��!�)�����Z�Z]Jٴncˮi#Y�J��
��S�����!<�Y��+�j$���eԀmD��T鷌9�"{�]
�k��m��(�,��܉�ӯj:FV�s�2)��_��8�0�jR
눠P�Ԧ`f��|{T�W2�J�*>��F�3�e�PdM�#����tc��T�t>j[�|�YUk` �	�:
ڋl#�	ʶS��B�-f�ZW�`Ɉ+G�
�A�n�J�%nYМ�z����\V9��#[��`��s,&�W[F��w�<D��,�D
�d�d;7��f�&��v�J�^V̤
�OU� ���+�[�� �w+�K�V6�v����/�ܜ�N�NKմa���l�&A�����/5UX;���r��X!�J�,P����`Uʣ)X�3�JĘ��,��,eY�0y��r/�g�eY
ȍ��%��Q�G^�ہ4�h��V8Lݵ���?T���)\�������g����)7F���L���"+��X�Z�gr��4��0��@̎H�rA~�Ha2�M���2}�xwrzr{w�O���x��������+'wG~M�������/^��بO_=?x����/����WϮ�?r������3ws�v�gW�7�7���w~��[eM�7����kރ[A�q�����?�����^�	ч�����/�79�qM?�y�D���1�7�)���s�Yy��Z�{���������������~ݕ�9�������ǿ=�蓓������?�y{t{qr������x����c��]ǥ�`n*�,�.(��5՚����%��l]����l��DW�i 43�]�步j#H'3��"�fj��c#��N�HMUw �.8��O��!-d�[��7���u�ؔ7Ih�{ѹ�#�Ļ(���W��v��'��:R��v� ���1�R�Y-3�HZ��n��CJL4`���&AvJ
�X
x��Ɠ�Nʨ�jM(�̀C�fc�W��5��aA#�u��!%@�M�
КY�1�}x�^��6y�	��2��I��Z�'��S�A緩)����蔌u�X�],��f����R�(4X�:�����#�� ����!b�6��Yu��G�^�L�R5�rJ]hAWJ�vE���NM��������Ϗ��R�)37����W �7�����(~�����D���,k�z	0U�nH"ݱ�D3L��ڦ�n��ǌf�}����:"�^�^8
�.\eһ����/+w
O�^V�;�y՛o�	��hu�53_�Ҕ�� 3���[��G.�b3�p�M3�휗�4�,����v�����zź�?�я��3������w�y��k����u��������R
g�^lZ��H��Wv�� Z�)��ik!� ��؝�%C����bW��M��UG)W� qwmo1�#	)�8�x{�;1�	ݵ~�!F�����F���Ay�`�C����Ʒ�� ���
ِg�����A�)�@yb�>����J�������	�O	�d�@>�p����t�p>� LIY���3K�d�n���^�ө��:�,����#��~ r"�D#[��;�C�ebH���J5��^��/q%|YAqS�+ߠ    IDAT�VӤ�oYL�B�l����[���P�9���jo�����������&>�v�F�������dS]7@Rm��4�0����#�A���iLг� r_����r�o����Fl���RS��N��DHMG1��/���g|
�@L�}e���a4j�Ac
�<�̠�%)"�"�*�xT��׿�d��DCƔUh ���Ԁ�/U�M� ��	�c�q ��3 ��RKVl�
mV�!8v�<����
e-G�Hq��i�� K�F��Q��G`#R��}EP}8.��O_7̦�N��r8�lNKqYjj!5E�\�ۋ��牗¡��x�&	��뤏���L_Q�'���8M^	�f�6B�a�aJ AW3eY��!���m�K6�	'%P�fޒ��:�S�fاzY�A�L媔��ԨZ�&�%����~��.z�|R� �Й.��Q�D��dʣ����L��L� �T[��@�:1��bg��P@9}
�^�u�SpCv�Ȕ'+Nm@�a	�H�v��(,U Ɓg�S.NM�j�Q̱P&e�0�1�5gKR1��l;���a�`,�-\\_A��t��,ML��9��8�&�K��Ň�+��YR��APX�D�i"�59�-��[� �l��.����r`U�5
o�bg�5'@��V�gZ0[��Z���@���]5��l��j吙��S�����W$5����)V"��Z�_I�z5�e�<R|&�;��T��Pc:�u�-y���F�P-�A� � �j��Ęe!�mV9PmR�挩�Q`�RUő��b�r��B"<�c2K��eb�e��&+@��h�QH���E-��GP2��d�Tk�{�v8	(g�Ł+a��B��4I�8^28�����H�2�
q贜֖�i��PGH7�B֫U@�O$���ս�Ț���̪uh|���A��/Z�,��'����x	$n�-@��}a�[`���k���a�U��ڿ����T�� �#b���̪��Z%
bM#���b̐��!j�ģAR��� !�D�K	X
���2��L|�#H.�ф�~n� ��B&��U���B<�k���� �<��M��h�y�N�o)��*@*���祀&Vŷw��h��Ա�����WBA Q��uh��,��p�xoU�3I��/�g
��,����őmK[X*O��C�fBx�x�F\����ˬ�KHk�#N�B
���i�iF&��H!�(ёc#��KYMR��E�Z߸�?xL%�	Z"O,�z��QH���>���=�055�w��:�D/� �؂DȶR�x�ٝ/Y��߼�`y��pџ���z�X�._﯏7o��.�/�o�o����?|�#���O^�����;��^yW���'�ƾ�����������j�/vǝOo5��ߝ��4�y��*۝���;}/��\w�]��m`;�{b�u!����zz��z������umo�|b�{��y�xu�}��x������������_��X��o��~��g?����>�=wׇ��V��M��7>�?���}V��yRv��p8j~�C�c�Ō�K�0Mj=��U�^��5�,����:b*�o����
��`���BU�&8�,����L��7v�a&h�j-��D��ĉF��H9{�$���5��{��^��ĕP�`'�PLG���Up޴պ��.�gT^�!�ȘL��>��k�i�9��qH�Dx&1!�E3�����C�����f�))4Umv�~����o�Fb],1�"h�H����#�Svh�d1�b)f#�j`-��<L�����o����
��	LS� ���I	�Q�ڭn23@:��R��_e[aA�rUfF�\���,�d|΂�@z1B��wڲ�Ɛr��t���ű$.�m��F��}�l�l}���}h���]�5���gC_��W}�L�Y]6��@�}W��������vD�m
�K	o$8D\;�4�����_=��<v�~�P��>�4������هzf�([��z���dW���Ь�՛Y2����6�bf ���D���.J��y:R��4����@:&)/f8[�z!IVV`���E��?�s������,ۄ�Ш9A^�vӨ8�){�\�3G��@ǉ9eW���6�Ia�N`��N�x�k��w�k�&�`N8�%���s�}�G���Ԕ���(k'@s��8ف���1��=����G!q(+��fl�Ӳv8��!�
�`��L�X gKt��|ڑ*��%k�h���pJQS[#����ú�)DP"`J��͐�CV�M����v�DK$�r����m�����R++�HgA g)7<)�]�^
ޥć�:U����Ni�Ә<ڈ����%�N'o�c#J��I���@��d)��!<�
�ܒO�S�b4өr�$+5��K}����ܮ�`�h�|j=�����2̆�(��6"�{�z���ȒỈ�@�A�l &� ��#F�4@)��e�x��������%Zd�L
_U8�y?Qy���5U^���N����6��H�^���@_V��
I)�R��$���U�0�#��W���e�Z ����h����+wPx��JX:�)V>-q�tX��L���Jx4K�tgz9��pRLP��Z�B�F��;&�{����
��B\��8����Kx{?e*W�0��i8�l�, ��`�^86>L��O��;A�u��Dl���AL�	�L_K��ITE��U�4��⼾��"h�� p"�Rm���� _w8dj!��g�Yֈg��,�<��vV��� �T�S`9�l;�<Y�&\ͶۉT��L����p,#���-)H�-� H�Es��a*�4��#AqD�	뫄B�c�t�A`�k��1¥pt�:4)�4y ��xU���)1��#�E�DSŷ�ȧ
���g
��^��Q)�5���ѯ��eʶfi�
O�ŝ�*q��aT�
��Y�j!��"2qs���Ň�[�Y|�Ȑ�#��<Kw�_��ŲSbI$D�,�@��e-y���� P,�*��8�S��P̔w��M8�YV3�`�!n�=�[b"ȶ�dRJM�X��Є8!C�o�:��Ȭv��;���ɢŴ�!KŉR9/e�)4g��2yUhvJ�E�H1�Tj���y�@����l���S��Qhb�Ԇ�r�>݁�k�o�4�x`/b�K-�)�Jx� '^vZ'T^ߔ���i��X1K�� DVUd~RS+�P*��.�7�r�i���5��
yx�b�?}���B7�`������,f�h��W)��Fk� �y4\�R�`��j!��S�Q8Y<�p�%�H������3[d�RF¬�֚j�Xd�H?<?�d�"��Z`���P�k'�p�b�.,�$5���6K*2Z4d�pUp��
�'(E���F����ͬ�x�>�`�&H�v��4���7��6o�j∧;AL��{���GoG
U�o#�L�<��ݔ�oI9�s�J�JP<K�<y��PW����
_ʖ�R���52@38RK�8�)֥8�MH�<@���5�h�e͖�h9�S��.mr��F���������/�p��$8�<5A [��|7�:U��<?��|xy���=��������7ono|4y}w�oƮ+���ʟ����|�;yw��C]�m�x�?��2�y[�J�����d}cӷ0�!ه��L�uM�ۜ����Q�� ۏN>�1��پ������<�'��O�n�-w����p����뎽���B�;\�O����?����>�߿u��{�EŔ�G3|���W�~������|t��Ս��g���sw���٫����՜̉����lg�p���!�@8g~p��dh�n�u���ʲ[K �@����Q�x��C����\���*�G!��Ł0�ѷlHd�x��.YS~��d�u\��Y�_�ٗv
<���3 <@ÿ�)o��������ֹ�����WK9�I6!�B��QB��:d��=��%4�����'¤�x���Q!�8�,�ol��Dp��ߥʜ�0��}x��#�����25)%f �l}F�l�R8p�Z�!>��u&�q��ʼ3-�@G'��B�QLJ���z	,��&W�`g�)��R�Ȃ���60�$p:SX��V�,����Jy��h��D e'E��*A�/�;���Y�SpS!kl��]#LY����*��$�-5ro0W��_��4e�S�,C0�6�:v��t�q׉����R�i,������?��C7�,C3qCkrA�l/}�\�R�lw�g-��&�sV[pS����FUb6�J��r�%�'�>�t�v�IۡTC4�2����g�/������O=�QK��"h�����hh∥L�Qy`�-�[���mM���-}����ߍ����/>�����D������S�;F�5�N��w��G%�ۄD�5�F��FNH����x4�l�-�c��@"��
>oGp�`���Ȫ��H=gi� ��8�r[�l�<j!��k�Ĝ�*�J`TRN[�uE�^����	*����N!�N��͐�Ô%>�xJ�׷	q,�Uh�$fb�@�`HKd������S�Ԧ��p3K"u/堐�Q�C�	W�S���KC�0����d+?��BN�<%|-"�j˪f�)#@���L;��jGP��
ˊ��y���ڍfUe�oR�FK�Q5�7��U"p�4��g8LJ\ߖ|H����u�hy�@�zYvYe�3� C���K! ��e8P9��k�{��g$?Fh��ƢA��<�1�'!%�,����,2�χ#���F�4��Tbkz!Ȫ���3�'�Rp��R�6ES�&GFk����o0�X�� ͐��	xn�_��5zL�]���|Ty�s>�kљP6Kc�H
!L�8����f��O(����!�)����#+@p�
��4�oM\_?�:(]h꒠b�R���h�!�D��R�b�t"H��ƫ\�T� ��\��!�I�qF\ 	�TN^#��K5��PVL ��T%�;.�8�u��4!�L���g@��l��ҒgJ�Ju��<��P�YyY���d��p5�� m(U_1��G;K k$AH�t��,�tN=����@��h����7*�N�᫲�e:b���S��� UՋo_�b�%�����A�u8ϔ�B ��-�p�{�v��A�)BS�%E'Aj�R�$"��rHÓ�����	�01�����Μ�+���-�(AHgd:���SIg�h&��k6&�䀯v-1YAj��jC:�D�Y�R���Xʪ򲧛
\��L�Q��8#�\�+@�^�F\�����*I��A��Y��pè����)'�U��m���u���Z�7���D̺@�F-�lU�_ã����hZo*GV.e�ɧ)"0K?eYqc�Q�o%ʪ-N��,#[6Z�]�����d��2͂�Sf��.N�je�YJE��؝���Q��Q�&)����XŪ��d�y�L�n�I�j������H�bx���*���i��R-eY^!��*qf��(�K	�Z�&,�ǄTe���y�5��-q�]A6x|�tdk���BT2��V�4���>"b|`�c�'�7*O� �+��[5��ױ������>+��03h�0]�M�xā]8�B�� �ْD��X�%��,/�&K��鐵���,[<-���rq�F�G���ĝ��)(�,�OPؾ �4Վr�̠s�~ڬ��4���m���m��1�%���4ÕL���ѪM�b�%��F��f��or1�/Fk�D 	���(�W3�D���4۾�l�P�{P�1�&�em$�i���ԎxxL�F��T8�_�`UR��=)���%����#Z�!N��c��d��^*d���>m���Rq�ho�˦� ���o��w{_��ͥ�{?���'��J�n��W#vչ�����̓��󳇫���޿���<��9\����������Ǒ�����ݛ��h�.��.6t��_���>[?�W<}'�x{t���H��g��UL�.���n�Ӟ�ޒ�*|�켿|��~�r��p�ҽ?]{������z�����������_����>����_߾��F�7�w�?��r�|������>�u�^>����։l��(z9�N�v����]�8����U�tu���L��������!��t�C��;xʲ��R�Ѻ��{1e�$��C�<f8-"�G�#�ʦ9q�@C&�#��1�O��{U`����܋π�wDLaj�M��L�FM^/o�8��c ��zW�xL4"�8=��P��Q>5 ��(o�����J	�7�l!}�6�KM��*\��m�8&�׺Á[��DpX1�I����Yu,b����q��])��YF�͊e;���|�\6�:����(k0�||�Ĳ��&�@<�,e	ҩo��Z��� �ȖcpU���j��CH�h1ˆ� ~����ZS��
,���܁�*�c�wi�7x�о�����I� ��oi6����:��Y	���e��L�FR�А@�*�\�_��+�O\�i�+D��m�-m�RN�[�F���W7�W������?��7B}��$<'p�E��9����f�
['mL�=i��4���Z��j5�~��+d8�j�Y����;�R�� �Q��z���	H���X��cr�g�Nǥ�W��4�q,�h�]u�}����ҡo;�0����i9ۇ��;�X�����
�*˻�@H�\�����1�Pʒ���sMO|���i
��bb��B��Z�c;7��Ƒ�w��HՋ�y�6��*���d�m!0Z�(K���VU�
��Xj=�C����
�)>�eD(3-�-�H6&�e�D�-c�i6g`
[�u�dMR*rj��J���5EX����l�([�B��vc-Z�`Y��@�M�B%p���R��k*U@�'�V߆�"9�րI�pK��:j C�($����������Fŷ#:R��	�-$^��!y�b�F���f����#�P	В�# C����-����� V#4g+e_��0Oh����V��P���.�=�9�
=Ƒ��9e�i��7��ck8)�y���H��XS|]�����(K�N3ۅ�'��D�WJ�j>�SHM�#�L���9h?)�1�^̀��ֳ�UNʖ�a�N��m
AR�p1�2~�:�m�u��8M19o	��ص�Cp�$r)L)��S$��1}ǅ�v���Z[�۩3��;P�P;8P!)8�:�� �@����d��R@�a����!8��[J�._ߪ���;�d#L4~ 	BZR(�*IA0�𛖈��0ө��D�e�<��|)~Z�� �X_dA���9:@���S�Z�ř�U�j�Y'3�hR�8��dq�K���U��'5��T���� -e#(a@�I��Y|�e;�DS�,��C�˖����%Z{o��iJ)!�0kd)�N�,g;jM�T)A>�7s�=������&H'� �m635H{G��T ~d) +��) �-=	�U��nI�+.f3�r)F�	*�1_*�H��J�_��δg�V!�pMU���U�lØ�������p�&�)
�j�8)�����m�=F.���0�#k�)���#`u��b�2Z[�T�Q�@h?3���oN�l�@K�h��<�G�?j�uD(F���b�q�
�E
�ސ�tl���I����aʝ�]?u^c�g����J�i�"�ĺ@�R.k��b�q��F��pnw@3���`��N�C�Lߐ��Ț�8��HʑtV@jL��͖�h"�u����Y{LM���V� e)�E3�ʭu4~�+!H_�@�8�QƏ�Ѥ��)�1@
��:��U�}|4��diZ�Y*i�	���Q���4�%>�%̉ܝ-|uķ�of���FJ	��������7֢�����񳬐���
�ZҁtÄ�����@�[�E����l���m�i���H52�UK9r����\�&)ƴlk��SasvuhJ����n���g�24��UUL�2
@cpHA%��&�(��%.E�@,%�T��������	!-hbx���1-�i�"��X���8�N�����rRuĉϋ{�%����{    IDATJf��mG�?3�����j��l��F��A&�ꖣ�
�^x���~�cp|��W3����1q�6p5ؖ~���FY#�F�w�2O��1;|�M;�Ђ��kH�d)lU{٢���|ވ(vS���@n��g������O|��~}���_
��}xs�o�>�7[gǻ�ك?�zp'R8����jw��\���>�<��ǖ��Qv�x�k������g}h���������������?�y���#����k�j��u������K�7�_��D�pw���:����|����G�g}��a���������ވ��O����������o^�������������˳�뇛������s����aM�9�����12�i��I�]�:ϧ�w� U!t{A��K%�4&�t��l��2f�8��+,����?x�DX���mG����с�!"��o��*��V\�����N��*2�7��y����^M��u�y�.f͐�PR[�8jk��h���^ކ����ǚ��&O�,�	{��H.�/�lIG;F�.Ş%d�K���a��֖txRm�	6C��K��_�R[���hLj��o)��Fh����m<bH'�%^��vJz�Q#��=�6�� �����3K-,����T[�F!�b�D#�"������*���Jk�U�'2�!-y�?�l�f���9|`W�Bp2A��p��]/GA*�x��I�E0d�&��"B��G�U5
�tQX-��z���oj��������D-Z�����uab>��h��>���V�;��I��vu�R�q����ٟ���a֍NB��ۈ"j\ٳ�������!�F0�ʒg�:ˎ�c��h�X�!�)6XY�e��
ZU�&������S%m�ы��o�����;���?��?9���3�s���e�<�<ƀ;Y�2;t"���,ۋ*�t\^_�μ3q��u�%�	t��o W�ǆ�����i�y���+���z9�č�`�w�vd082�*K�- Ťw��R�)�&&%�,��CNH-�Ș�ZTd���&D��0|�Z��eW�fpj�#��I�R^O� �q��T�a�4 pK&0LH���t�p��bZ�e�t����ƙ	U��!�k�f+�3
���ٸ� "� <�A
�2��h� ��E�W�o��d��i��KQ`��8snJK3��2���.��2&��l_R��/pƨ�W���@'�&�
���R�H1�R�Ӌ�@A��Ē������)(��Ń7���곘R�Y�B�ӎ�t��LL)���"��d�U��j�0���A�F0{�B�4Y��'4O���3��٤��>�4LB���JӬ�����7/�����"�m�$4���,^&�"(�'�\l�l ]�p���m�I�5~�9;�hS���>$Ц��kԎ�Յ���W���,�e���	�T�:=��W
��{�#������f#.��o_b�rV\m��#�d�>d,��ɆWRkYA%!t
��.h�vJвa@��u��K�#'{:����s�5I�*%DGH���q�b��� �Z*���j��A�{5�FI���Q�0������N�����hZ�b�&�r �
�.e`��:\��p��n��j������肤�ќ� HD�ڎe�j�j!+������UE��R���G^қx�Wbf[HAm4�N_�;(�!���TYHW�!-3K&�\G�I���]C��Z4��E�������]���v�
Hy����Gk����}��Q�dy
�yHKq�����T0LGM�1,Ų͆I��B��W�%��"�A�x��;�ȩ�i�vp4`ݩ.+f��pfx`�AX���]�
u\ʒ�j :��r���:�A�PyZ��&p�k=%i�CH�RЩ���L��� ��SRh��&�l��T\��"޴�kAL���X�eHLy��A|�S��8��,+�w�Lޒ/�ؗ�$��p�l�m��F�]�d�Ml�G	k_@yr]��<���f�tK+������������!�4ϔC,��& ۨ���P40� �@���L�����*�M1k�t����f��R�pV�VO�`h@��#�>�Xw�,&$YK�)�G(�s�@�,M�Y�똖�Ap�J3�������p%!�kT`���5�Bx1��֤<��ܟS(�9�Dᨩ��+Nd4��8����iM�<C+��nD��6�@}�I/m�WJ�,�Y��4��1�{lh&H�OVM0&�F�4j
1q������H���!�d�,�c'2%-+3)މ	��A ��%�wE3C0U���	����V+[�v�4�7�\&��!@�4y"�{H&�>��Z�4��*
�V5��>fU��� �-;@�8��сLJc��ڥ?�˗�4����Om�ϟ�y���.}�������.=n�֗3=���wc��p~<\>?nAz���O}Q�w/�=o�n��Ԭ��x�%;�\�'-��1�W�{/"��e�M�L~G���z��A�)m�^�����]9�ſ8��������z�x8���=[�xfw{����(�g�϶7��v���uS����@����<�[�4�����k���\��w�b��ɶc\UC���pUY:b))�l��״x��v�`�̻݊�)��=����B�g;.�,+�W%�/�L��^���R�=�ҩ�%�v}�I�o�}�!&�9 x��{;ȞXT5|j[ݣ�ȁ�Hu7����<f���5�>��-���[j�͙���f���d��kg����w{L�[a��*�4"ŊI����Bj˯v~�Bc�cFn&f�GV�B䪀�[��N`Z��B��t�C3_��U�HY�'[!���5X:�fC0��˲Aȩ���E>�@���O��������^��$אGa�)��vd���:fR3���ʥw��s��b%�"t��f$�ƈЎjG�xu)���P�>Zj㻚�n	��_����.3��jA�Q�� ��H>M�P����}�v�-�}]of�;��پ������)�b�U��y۔J�2P��F��L1	�P���a*��#���tx5��\ v�p�ݺ�	�D�W��,�'('��\S�������������������;���_��+�������n<��~Ԕ��)hA�� x2�������۩*v�5R�@��%��V�Yҵ�)�8C"�5{B��MJܵWhw����1(t2�6��,��c<)�|���p1C��S�|���r'��e&i*�p|5xz>��?�������pM�l{T(�g�m�Βf)8��C 4S+�����K9sY8�ԫ�u�$�˞γz<=(�u��������3!��p��1U����%5� [�6����4%��ϐvJͲ����J*���j��tZ��8���E�4��b�#2`Up�㋁E|K33^9�X��0�,h#�W�������Qؐ���kOO_
@
�9iZ��H�T}�K_�Cp{���$�r3+1��r��c�O\�U M*e�@�����E�������H�S�vp{h���� E͓$�Z��"��lq7��f���F4M;:��X�ۿ��/���x���T���LH�Cڎ�N�����cȘ��&����^CV��Ҝ�ñD�B`����fc�dJ�����"���~��@��iG*�o0�������U�ױ����1�����.�~�]��T�v�1s�� <gv��궯�o�94M�l�R@R΄&$��F�X��m)4I:��c��_#��ő
�ܒN�e)3���ZLǨ�ӅT��b6a��m�2ZM���68RV�J�B�KM9\��
��(}YH�-��#P�V*YK�VU�Z���\?/�&�&� ԋo	�Cʆ���]�2R�ؐ�MgZl����,q"e�d���=t�@j�!��tᮮ
R#��3�y��QS� ��Q�����r�EnfȘr`��5B��u����+TB�²��#��m�!��<�RS�[�ײ�f3���-4F
��SV?ܲg�f��73ZcW��s�dk7�Ȕ��6��h<�E��8	Fh��&��T�����	������ _m3 %(�M�ZC��_�o[.[S�챽�VX�z����,q
e��c�4!62�^�^��]O�y��zMğ�T_�|�ŉ�D�T���Un)��t4!SiZdqCFvS�ݔ� ������q����kY �((LDP;�f@k���t��p���C��Ҩ-$b�f��4�tGcp
�6RMBd�6KR�Q��
�I�Ѐ:V(C�j_bV<�0����7��V�
����Bh��U�d��b������*5�.�!b�����x�_;�RI��rY&K��r<�2��[��c��i�z��&~�G"xZ�-���^&�9���#t�*l�1%�Jh� �l8�՗�M�!�պ.��X��[�rӱ�$��JV �T\kA��"e��M�e�R�x�SK�b��·�id��^�R�e�	����)wK7-PId���n�~���_����3�Z&�宔�t��� �I��S��T�L�B�5�v�e���]�������L3�~�rP~�e�(�ƣ �н�����LG#�8�_��Rۀ넛��-ٚl�-�����TGK�W�4���uL�Ť��羝��S���wן�=[�ۣ�P��%�����'��߾|8�E�ピ�~���/|6y��;;�_�<�lwsw��?���<�/}�y�������y��Ѯ�y����hB��kqq�>X�/a��^|s�߸���Wh�9mİ�{�g/^������ӏ.�?���ʻ��-O��s�������?�hww�O/_�FQ雝�xx�[[�ҧ����z�;^^�^=쎾�f�f|��x�=d��ױm'��c7�3����Tb�\Y1���VK$D�ۿ�D�=0k���`�[�n'4%��D��.6'3�.@�< Sۦ�
(ė�Xpʷ�G�Wl*�^�)KS���C@���%fb��b�h�5j�q� �`qI9�6N�#�7���{c�5x8��f���� 4*d� Ɛ��'�!�S���8�7L��&��ӡٓ� �]b�v�ぬ �,�q DVߎ�C��R�!x��Ӄ#�2@� zuh�`�^RUy2�Y��b�x��G�If�f�������p�*��SΆ�� �m���*
�=�c��e�+���g��Y�0}��q�9���Ǒ*�jj*����,�(4e1O'�x����Rsidg;1-��y�뚷(��f�{�.qjF����$R
Y�k�Q��[�m�Kg3�0 �Ix��W���������������<Pۃ#�A�R7�l�X�D��c�;�l��4�(T�i���E�ʑ��p�����`��ѐY4��
1eq �Һ���P#����x���.����ů}�k����	�,>�1zo�q�))��L`��du
�^�S|+]�8����֑�1�t
(�p�.����df�f�`���,nfA�,prD�[*t�iMߣQ�Oё!�2q^��C�� &"�d�c-��͊�VVr�U�@�m�9S�����6-_a|�L�A� m�Lǲi+�����jg®��e	�)4Ub� ��k��œ5@3@��8NM-S�Q-��$�%�F�fz��>/�V��#ߎ�������RUE�S`���u&����i𕧯i��_��T=�����=v`<&��.������g�N��Ԇ/HD9B[�X��Cб#B��� Cq�|��s�,g�I�� ���2q�$P��1n0�*��Gk�nc1��X_y����ǐ=)��#��j�J���]���+i`�tat<7���\73� f��g'�p�|�uN�����?��Ē9��вQ��d�G@�L�"���L*iS1�R�/֗u�%���#kT��v��|�������	�y�N���ˌS�L�j�����̇�ǯ�7R4Y�#RU��Gɚ����e��"�Cs&R3O"�x"���v�L�A����D@V5W*o���1��N#Kd
MX_~���MA�!<kfxdUS"������He�,�2N4K��o���F��ֽa�#�X����c������v5�c�Յ�R�V��;�S����̲�И��,�� �!4�G'NY���8�C���L'��Z&B-ک��t���D�쬴&t�!G�,�T���� �xc���Z�A��h�8�����&a���IAJ@m�+�Z��dێ�T�v�T{��]*2Y�T����������3�e�D�uV�LlH�@I�������ܨ�h�
-y1Nx󤦵%_�zI�w�v�pF��}|�j6�*8�vR&)Ka�b�*K}-;_�SO�_-���4d�lyF�.��U9��݉�90oI����R�i��tЈ�@�L*��/.K��0�Zօ���N����B��h�H~D�@L1��v@:�l@�T`�+�uj��뫑%�fk*�i6*�����mv*k��1Y��mu��1���vѫ� ��YM
���(�ԝ/5�����ڑv�LG&֋���7 �H���4	������P�R��`���RjZ8:&G���Ӳ+���;o )8��3���y˶IY��S��7�dh���� b��5�Ơ�:m��+��I5���p���6{!� ����Z�P(%(eIJ��) �;`g§�97���t�[&+�K�x����qZ*Q޹U޲FD��x
u�����W�֩��l�b&f����!�2Y~vQ�j垮׈P.5��Q����h░�d[�	lA�R���U�(L�hi~�߼���[R@�G%^#�H��U�]�0�S"ԜI��:�9�D���&Ē7�98�r�p������Qv$��R�_����f����B��Me����!�&D@�g���3�e{�WL*��wM��TP���><\�3�v�����;�����a}�x�O�G5}0��>n�H:�F���+�~I&�_������q������xw���yvs����_�<�����p~}��wn�������c۱��>�nk���k/�����[��.v����z���ȁm���.�Iڋ������0��\�\y>��d�n����F��xs�=\\^�ö�g���k��{����\�.��{����G�v��|�i��qx��3tT��6��]���~�.�H���ϥt�m�Ei��w5�V��]d6�txo�ͧ�R�y� y�23t��:��5�e��$��8f1�r|�cRj-;K�I������Ah�[���)N��S�Τ��Ua�ԼGԫ���1�I��F��:���Rs��� O�5�1�*%�&�>�	ښZ��7��ۤ���\��v��Z�bfS�@�A��B�VG8qS)g�<_#%@%L�⍾n*_)%RUUN��h��*���o4J:ykf���
}�&}{�VM�Eǖ�@���)��)��!����/qfڂ�ȶ,ş6��+��`ޔ�^���T��C��p�t��X� /6*st�nK|YA�<�邠�9��𖘂����]����?��?��X�4q�����%q������f��}�p{į��p�ZȪ%�}��Uy��?�����i��;P�3��WC(n�<-]�S��$�Ĵ��T�שQdm�g���pT�-�ui�hn�L9&6[�S!��>f:���T�B>B��x{�{���w���/�������>���O~��nOm��P;}�Hل����C�s�2�����9��l�a�eG�l�@�f�v]��b�E�K 0(t�l�TZ7��<t"X�iA�v��"(�2�����g�Q�mEkM��v��N�G�Y�����TEd�X����]k�	kG���S+�/o	W�eM9&��&b�e�ڒ�	o~��ץyxjI����W��&.���U�2
�bU3�iTd��i�r��V�lR]K%����IY�d��Z����Lj��T����ʞ��Ň��.�B�����حK\�&�8�ڭ���-�L-�4�
�g)[\�i�S2�@ʕ�o�� ǜB��3ʵ֑gD���:z&pl�    IDAT:�����0|YkM�B�C^��6m�c�O=F��K������6B�D�s�7$B�<��i���j=�m�x��Y"���N�BǈO��?����_��Wȶӿ����+_��e����'<kiG���M�H�F�g�v�)�7��׮�-LRyޜ�㍽i?�gw���B��rÐ�΁ǷA�S��I�gf�:Zv ��6���"�B�O�%�a����W2}�@('իL�Ry�V�/FS�� >"3^J���Ȇ=��LҐ��bJj�M��S8ܲa��[�f��R�sp�u�PI�����j�����q�Bt�̚Y�Ʉ�;U��,�!C0��E@�M,@Ա^tX䖥�L	PJЎ��	�-�2|K�;Cw�rH"	b��t�sx�X1� ��~Z�rzAq���[
Bx���,�Z;j)ˀ��cU<� �ii����-2ڨ�̇��[�2CGAߖ�9�(�/�vJ��=�<��Ш]�F�XvY��<�w!zԄ�5p��]�م���*c3C��e�.���$۾Bx�O�l��*iw��k����1 2�P�TAUZH��ŗŁ��0�)�!X��
�GK���pct��� 1�,�%�l$1���83L�D/�����4'U��j���ْ�`�&�ϼ�xPK�T2�d!-yC�rLdY���v&@�,��H>�Y��x�że�6��ދ)K|H�Z֢ \,7��	�N
�=7��M8�j(F�B�r���M-⋕Hš OP�y(4Z12���B<-(���J�,�lNm����N�,��Qs2�-k$FsiT)ѥ֖Rb`�d�(������h�|�0G�lx-dVK-&�Y��Ѵ������3x:�e"<Z%�4(3���RD�|{�ZeO������AF ����_�US
m��&e������;�||�9s�5�6g�G��)$8j�b�n��S��<��>��ԽBY]2)%���g{��c�BC�&��n�On3jjDSյK���vxU�r���P037	π���=�X��Fȣ�Z�pA;JPIdA
�V��(U����Ӆ��QVk��!�������g?�я~䗻f�/2Nd�r8P�	t�K����+DWՏ�ťĂ�"n/::��J��[����د�5�W��Q"ʻւ1[X���⦕U.VN_
b).�Z>+G�!#u�iF���-XU���/-ڷ?벊������p�>�=�V�4�bgx�u���g��%no.�7:��<��W{�i��^������g�g��<h��;�T�>%�����g�u9���}��{��6��E_��gR�@������t}�s����gz��Aڛ���?yuws����Or��=��i���Rӻ����~�s׏��?��/�Ύ�߼���Z�ɞ�Ώ�o��}�z�O����]�|�dG.q�e״[�S�L�T�NA�-������<pY��T)�@���0jb���o���b#���8�&�n�K!�T�nc1�
�d!�)�3jb~��Ad�X	D�����(G�W�CRֻ��U*�]4^gզ��k#�ۣ�UEM!\#�B� �c�� g�� ؜�~z��	Jy>)�C�FJ��,��-{�	(��Ӛ�J��Uh<|����W��zH-f�LI��#��p��nJk<��̀�f��C� @ �Xyq��,e�jL ���=��o���%�2��$/h��g�3�1��)L	|��Fb���NKf�Re��p�q%sڶ�`N� �v-)�g\����u��e^��n��㕅O��#�S���I��85݋u�v��P�?��?��_�E;"��ja��r��m��;��EFH�����ޞ���M���Ǹ�2��(��TN�Ɖ��_���K��IH,��T��7��݊u�GcDy��,&����O�����m������U��!)[2dU�C�۝8�Q{1�7����{~��z[�`��o�������j�կ~���U�N)M/p|������F��D��i�W�n��A����k��<��'i�*���
�< j�+�ӧ&A�]/؄����1 h���ͪ�hJM���(`��G/�x|-�D����u�y��l#���\_偼%��TEVqK�1�V��j��Y�C�v6l�j'kI$eޒ,>���a�[
����Gw)�mGJ�l-&q>Y4�*��	�2�Ṱ�:ϲ�
y�B �r �1����h�d�+��Z���L�U	� |1�*֩
��Cc���� żB��,y] 񉄟���SQk4�w"��C�S�����i�T�*o�#� �I��uV���Nؕ�]S 4��p�0Y�b�q�x=>�w.�x����#���y[-���p��(�@�$��s�����$4��.�@Ok�� okpR���/��7�����5���I�� �C
2w�Ӛ�9�U�̫��C^�!���/�����<����q%>�6O��k�c�e{�hgr]�ƶ����"�3TB�������
⸤_�5%����9�)5�1xV�X
j�y���@G�*��R��i��7����<�;s) ��$MY��u���.40���Ph�D�V�,Z�@q[��GX]�s�L-�0-�O�ڐd����pѮok<�-�� S�f�);7�TY��u�X�&�<L
sC�1*��Dw�h<�T4�Y����Ưi�o�r:�@#*�,+�_�]�*���dY��	L�T���� �����8���)[�ld�f����PeDH�������l�:��d��Y�����b 2�I�֥R��=W��<b%u�3
 '�$�`&�#)x4�PJd�E@J�9��c�X��6H$�X�~��=��z$����&��KqM�l���K�j���$[�e�|a��|*"f�%YKj,��T:�hv��3��m���G�+��4/%ˤ��晣�B�U��b�ݪ���V-Ĳ�HY�!b�S����`��n�j��8s�P�(�fN(�6��ۻ�q�(������m0^G0��6��uo#g3p�FGm�fVUy{O?2�Z|f��VH��!!��׷Z[��x�2)Y�l�4Z۝X���=���h<���Yn���.(�ɦ�0pԊ�b��y8�L�3�)Ac��5��L�C��jy̎�T߲�T�0j�������P���,��W��o���`p�?j8t���1���NU��W-�l)�h�r�Rs5�#7�&�����0r�R�y�:��7dR�n��-k*�D����n�Rb��;A?�^_�٣H�3-�SU�3�� qY"b^k'#��I���4f1��»"|
#k�u�RB3#S"����x��k׍�(�Y dt(A6�g��o�ڥ��e�E�1���,S �Ln��y���/���	Z*�Ut������t_��ũҤ�~�&�R
�j�'%hH7����O7*�jT}�[�l��t0u��>����Ȳ��9+R�95��m�%����ĢQ.�CX�U���_w��|����뫙ޛ�T����^n��}��������g�$��;�և�ެ8��;{�,m��ޗ؟�X�y��K~r�����G���od�?�����������{X]qv��^��'����iZ��� ԋ���ۛ~���慿k~��P�uۻ����ޞݭ<���A��=_�>���^^�ֆ/b:�o�������z����/�R�1�o��[t�L��z����k�KUW�1c�3���
����Pwi�����wOƯ���FR�р�:��^PHs+zO	2W�o���ԅB:D�5������.j:-&�pd@
ֲ�d��D�AaH�yx/ڛ?��#Y��pz�(wV���G6�%�F����R��Q�n�*5�&��)@ꂀ�C
(�異Rƨ
�����ْUn�
�.�͚J	8�Gy|���?&����&AP�{;��U5���%G��d�y1��]����r�"3�	15|^�\6�t	I
(�g�B�`~U!Nk�{�{|jm9��IU�x�J1{��/o�Y*A 9@ƿ��Z:[H���v���t���'�ә�����ˍw8��=%p�8D�j���w��j�����/�kW�W� �h=�z�u���:�)S5w�%�v5u2d͉���vJӗA1��ۻ����}�����H�m���o}��_��i��^�Y���N����8�K�Aq(䁬��pL�ע���>S�D�M����m6)M�wi�M�/��ۿ���Q���V���.���4����Gz!�W�s�_��R��A��`Bd���M�u���a(3d%Z˶A�f`�t�J ����W6�m?�:�޻�@AS��b⮺1 �틦�����L_�a&&��#6�aD�m`����$�v�4m�e��P@SV����^�R�|���	٪׹�# M��!�l��3�����<�q� )��7^ٺ��kg�����q�S��h4��e�i	A`J���K!��S+L�W�� ȂQ.V�>���!�d8A�4y��K����)֔ƴLo�Q��(l�pKVG�!��wK�#�G��owR��&����O��� �iw-'5�pf ��y� ن�9�-;@�t���3�'4W�󌥔���IlY@�<�$�@���'1"h�~X����Ӎ��.@O�j�+�m�H{��ާ�xJL(E���S����j�H�iЋ���=�b�S��!C�㓼���eM�����پ�R���Q�#eInF6f�ם�%��A��s+N_S���Dm*FбH���q�).�+#)]pTɚA�[���Y#�_�>\#���8�Y��.��Z4�J�^::�����Q���B(c6 <B�i4M1P�d���T�p��m�i�e�:�\m���B�`���0
�,�,As"Ñ�
)~�>n9�OY;����8�@Ni4��;��b�Tq���i��4����l�Oy�ƜB%��y6K䴅����N���Q;U��1�Z0�6�:��tb*!.�*�,�g&O�>?c�q��؎Ti.`Ԛ�X
�f���֝-GvY�!�ɩ4Oe��*SY�n��z]�(k�$�&���&����@���3:�.������}�s" Dd =����¤��j8!�@�T���<�w�,ecֽ%BU���۹Վ��0!�Q�t���V�� �ï]�I�:Z�<����2�J5��]Pt��Ԣ��ӷ �)d)��L�$�<)�)i�ʁU�AM5wfU��B����N:�jkR��e������f��3��Y-�\*����Დ�C��EjR,|zY�8�&�adSn��:\k��N�J�T$��(`j�r�<��ƫV��J�#VeN�b������-YGݥR�$H�-q
 M(��� ��O�:F����Fj �h8����A�j�&(�"A������)q���3�3}�l���.�P*��:���p`H`qGMG��O�HJb�#�/L�+��d�m�U�?��t8�@���>�PP#�T�)�d�!)���H�e�1񶇭18�B�f�X`H�'XlN�bxL�������ď��U��FNG���C��qex�=��3M#Xl�����c��q�H��s���B7*�����	�'n�'[k:��j9?�t5���T����	���t<e�.����`X#MJ��
L�<qĬZ�)����E��#A'�C�BZF��r;������?�OZ��iӢ���K1s:��~��SN��M�Z�����A�����Bx�����}�FV
�';�-(g�8mYМhU��;���(�2��*1�G���o�G�&x���8妣|j�7H>#y�{���%Ow����Ο��y;�{��{?ҿ����b^�ϟ�O��n��ߜ������<[\��^�>�w�z�ً������t�#���nγ]�}�˳S�ғ�w}�#������5�Ո�Rǽ?�iZ��Msm�9z�sY�P�b�����M�����}ss�����u��x�����/�=���z��׼����?ן_�N���{�������߼����S�NO���܋��5O�޹x���>{��o�p�Ԝ�N���!=LJ���X��Ȗݷ�ҁ� bGb���Vޝ���-�.r������F���vL�[�G�좑4��ɯyF�8��懋�6�Xm�&LJ����#�Sl���J�Xz��"+�L�������#N�	����,}K�p-TE���i$��XFhbF�xL%Lm��3 � _!��}�T��<�Mh�݂/�Ԛ�g�;k_h��T	D�,�� ��	�-Y��w�mj�d�UɊ��2�u1s]He�E���������W�x�pfr�&��[ ��e|
��X-'[m���-���`<���FAj�)�3��K0wuLK���Rm��ɔrP�L��'�بM븘���|`���b�Wn�Z(������n�Xw�)<C��f�S��@����Ĉ�%�� ��k!f�ߨ��8��I��f����2?�>�b6z;�G?������~�����/Im�{ZT�Ob=L��&Ѓz���˶a�"vR�?��@�NJK�JĶaz��Y�1� �&�D&X'���lj�F�Xy̪����mVl�v:55I- �b���%�e��@�g�A�OE|,��.�������>���M���c{7pLY�# ){�u�t�hA���e�R��[���|�;^��a86��%�N��y���N����R(�L!�MG
����w�U�����)dżl���R�������ډ�
J��%�]���Kjv�.�.�B�B��em�Ԧ/�j��pH�lK>}�i���hI"v�0�IV5�uIv&�4�cA+�W2��Ѥ�ˌ$�ӑ
��b��A�-eIY�(o	Xj�G4U��D��1�� �-�X%f�p �k)���و���B(+Q�k��y�,2C6��`�ʪ���a�@LKq)Ǣ��񲖼xJ6��})�M� �2|
4����y��)�C\�9˾�#e��@|�0��mxK�Τ�T��j�s
K�FenB���p1>��݉`�P��C_�':��� �7����ffZc���)���[���fK�����_�B/�Lk_��Ց�	�t���ѧɳ��@����@H��p�QyY���iTL }�D
R����B����8�A�� 2�	⾎|I��'?�	���9h���}���^8C��,[PY�	ӡo�v-5+�����bZ�Γ&S�V��x[r=�lG��O\j�|tR�V�vd!���RD�ƀ;ᲆ�i��J���<NA1�lX*���bV�#�'��ٲ@-�Ѐ�㽧܉�E��F�X�2�N� Ϝ[|���ձͦ��4RE���ZV�Z[��A~k<1�p�76Fd�	�3M�C�5���-��־��N���&�A��w4Up]X�R����J��є3���O�R�"�V�m�5��)�R�G��%�����o�q��
-�L��g9A��3-�S�!13
Ȧ���Ra�3v|"�y�Ԁ�e���L��ӆ�k'NA
hɤx�<����yR=d �b
*��'P6� NC-;��1����E�%�'� ,��&�x7�IS,�&�i1K�]P�/5���Z��BA��UV����R�%��|FD
�d�M�U�)��-D�#�T��o�)���(�/�\�W"��%�x������B7L�&�xG6	��!��" �0e[n����l��c�p N�k�;�e�åLUFGձ�E� �µ�0��!,4���2���H�,ϔāԋTx�*��D�_\v�?�D�%j�Z�$�=��y�1㠱�&
��@	��ƛ.��R�o)�a	�AI�q�Xʊ�@��W%�Ĭv�b�lˬ�(��);1N���.�!�8
�(�ؚD9�w��4�����ZWmN^N���9Õ !��IАb��w��-��W�a�+��&�jY"k)k��h����D/)M���gp��c�Rp�<Z�d��j;LK)j��~� [ �����"������@^	�ڶ��~������M
�2}�JFM�u�m������㌬���f�'�����-Ŷ��I�����@f�ت�C��dD,�0�~�� ��x4u����*�    IDATj�mBY��V(@c��D��	d���������r���/��w����%�0�������ӻ������������峇�u��vޭ�qvzu����/~����~��������k� }���w}�&�>�7/}@�����:�y��S���d���Y�/��a�~�s�k�ӓ��fQN����a���n��#��7��� ��՞.�v�w���6r泣;ڇ���>x�Go��rxy��p�r�*�����7��ޟ��]��}Vӯ�=�V�� �z��{�렞.��4�A�������Ku�@«Ap}-�^E��É�u���>=��+�o�'LS
����i����H8�<��5mk��b �-<N�J(��%A�Cs�p�^�q)�BౠE�� Xz�'�jS�/з�K�k�mJ��%�T�ERٚ6$)L�3s�Z���� ��9�:��s����_/"8)�fq�N�7|���'�vAD� D/Ut��wf�Z#3��k�ר^�fChBxR���e^a�j:����./X���������I��M<Y��^u��	�k]jh�����J�Ώ7�Rd�tڅX6��or�,܅H"@��Y"�^��&����nH�ց{�;�>ˡP����3�u�C�MJ�i4�1���@o�������b�=�]U�J Fm0:�L�@��yjhZ�+�v��)����5^_�0e��M����|�0p����?����5U�������m���/��&���XD�[ܸf��I)�X9Y8N;�|�C��u�JQL-�,�����ȶJ���G(�� ��`~cԝ/�Vk0d C�j �
����=�4�[�bXz��vt�91&��3רZ��^���.���i*~�����đe�p���:[|f$^��*�h��2fi���I����G�FYo蒲d�´�yR��q��Y�u���#��}�8L^������6d�Ҩ4U�N���S��V_�I�3%p"����!cR�U�Z+IG9��+%��e
�!|���@0�5����������Df5�);���bB��k�iI_�BY]U!7���j��cPwJ�i�T B��ઐ�Se���Rh�*�MGJ̗�?0e|GG
�3׮.N�63	zL�:L�y�U�$[��	(�T%֨�(����5��e�sQ{�����d{��b�@�����g �>�y�S���̦#�u �FR.�����#1D���Ŧ�Z�
�O�5L8)�hC;���<OJ��tQR시��Z(�Onΐ�������M�f�������/�$5��!ND 4!P�7O�+�6�@c7���q�5L�����ܼ�4�-חTLM-Y��6�#���ʑc�6d�'E_@ǥt�,mX@�Y��ā�0����F�T���k�� �[��C��uz�)�#��-�^*ā�5�ӓ �T���	���T�B[G�JM��<$>B�|U�۝=ڗ%��hY-5��KH'�f���ʊ���BKӪ���򘖘&�Z?�4�-Ų)X�K�Y˔55�0�$�X!�A��3�1��v�e��2)qS<�6PS��
}��<N)&05q�y����سP%<�NL\/��@�"��RUY�:yA;jY�<>S�xA�J�b��������i����IM�X�eSi�N��p��4�&�#��8�&��+ĩ�vN~��'�,���3�^���_I�ݾ'�X!BS�'�2�bAC����1~L�H	:���q���1�2�(��ᕤ/���d��ڝ���zI�;P��p�/K�52��)�Fj�w����<s�/F��,Hpdu2��]�X��ߎB�����^/)%�*)f��<b����-G_�8x�����3��|��RFb)�#S�5_V5K�_�g����O�lK����Jѷ|�Y	)A��+�ā3����^ h�F���0e�0;�|�"o�70��d��)'�nI3��,;�y���KP�Snmb��G��j!����yV����$9���U���Ų������G+}YK���<;搲�׮�Q�sj����	!U��oxؖ�͒I�t��h�htp�:�Zt&�ᘝL��Ch
b��!e嬍�y�}%��F_[�o���b�l��=�XV�����V5��l�D#��1"X
���u�<�K"s���GQ6��N�Q,���Ɂ��@�҂�з�q�!�5���F!MA�)7�OF~|"{$
���n��1����(��@��9��S#���,�3%ȓM!A8��㨢@��yx1Nj�rr�ľ��}������go�.||�ȥ���!�x�������eT��ϼ-z��Ho9�]����=�ڷ��韾xy}yuz��������6�����������2���Ns���n���y/�K������la{�r{���u�g�"��Su�pw�l�qw�|w��h�3�D�'����|wz���g��w'ן�����wΞ�x�տ>�����]�����n�O]�������J}}�������Ϸ������vJ���u��ע�ş�br���I�6R�*�"T-�u�޷/=u�1"�j@"���h�udԔ����ȥ�gP��,+5�Z)�D��	R��b�@;S�Z
�CXU||
�1��~�����2��A��:����E�gZ��Mu�:�Y4�]�v�<|��N�v,�ȼ�)��1(��4�B��7����j�I�l`ug
�=9(d��&%<e�7v���c�o��1iB���5mfY�Fέ��@d���<{�����o}�'�:Z�]==5���TH�QP���ъy-V��겚m���:�R�'2�1)�y��I��X �e!�ᴌ!.P��[��̮5\�.��C��K�5���l��|
�<o����2IA(��^*D����_�'&eT��\ ��7)�K�30�1�N��FhIcZ�3��I��:$q�]7*o �����}���U�����|r4���v���3��&��%OEK�9,�� ��\	($
PC��B��|���΢�U��tQ�cy�J���;�!��4��ڠ�����e�?��S��?��K�ĉ�l|gbY���uo��Y�t�ڠ%r�d���.��3�{�K�ݩK�H�hG�Ů.Ц(#�k��	�
�y"��-�ISw�ti(����B�ۊnD�č]�	�l@�,+Тl^V���@2:F��T��/���;D,�/�*~'�5�]#%%�+/K�R a��l�6Bgb:H3��M��+7±~"8l�x�2o/���j�lw��ttt:p����י���D��#���M� ��j�.EG�+Lmc-״p��.�2��n�N����p�V���0)^<�ȼr���˪�<D��%�NL�H%R_�R� !hY��aHѩ]|j!���C��^uQHǗ����
��'�S%���mڞ%�4-=�	�m��?Y|oL���Pm�-��Z����z��7����
Y"d�3]z��gR!Z�y��O2Ȗ<��gr�����0��e��0�]��i��X;�h��I#���D���<!��c�Ȳ�����9��1�
Ƿ_d ~��DжY�7����?[�S�"�b&E*/���4-A��U���H�o`Y	�u�B{����U��yN R#���ow�C��+�*2�"��H��V9}R��^q"yL%s����4�B�gvDY2U�P.M4U��L��e�A�+��U�v�<� ��;
d��_4���Lpj�x��Dn��U�K;�C*N3����NL��v�&�i�v�C���4����!_��#O���~
�F��@���,l�<~�AV	��r��c�a��$�����BK1�mfPI�6l�Q�Zֺrq�8���e}�t?��a&�.W��U�EJ����B,��w��z���y�����te�i�X",��aؖYjm$�ʫ���O�q�oNY`(�m����4��B!)��坕l�!�/%�Qc�h��J�($+Um��&K�R`�V
�aBҙX�<�īcj=6BY���U�� t��l_��a2�l{\�̀LM������U����i�B1~]��Id�dgZK4��-�Kp�����*��
!�ĸ@K&�-�/ N�T�<M��kW� ����/�BK&TH�²�Z��Z')e�������l�8zɊ��[��"��0�f�
Tn��1nF���*�*Y�%C((�͉i�G�u�+_қxU��)�l��QCBR8��ZH�]�:��_ o�/��^�H5[~�/jj��b����r����q����!K���'0q�5X��0]��CSb�f�t-{2� �ֵ�@�8���R�e��vx:b&�����w�<��N	Da^ �\v�_=�����v�$CңrȐtzad&��d��?P��`zE����}����a�(-�:�v�P�.�@�l�L�T�եBH�,>���l��7$fG�rq�� 4@]��xYU�GPBُ���lwq���x/� |%�BHOw�����W���Ԑ��v�3;ұv�W��Ց��ԋW�ahRP����P���3'�~�3��I��؜�F��b�|K~�B����Om��M�ޯ��-o����t��ͩWͽn�3���Uޝ�N|��_��̧��]��^i�}��:{}��̧/������������ݻW���ӋS��䍿�y�?��ݲ���A�K���'$]���_+�ѝ�i�����Ü
m�!��4���6�ٟع?�y���� ty���߸~v��?�oP��sO��ӇP�w�_����/�n�]���������}}�9��ù�7�����g����åO�]=����we�o�o��Oc�Ι7H����rE��Lk�m)`8��
� pͼ��l8P�N�6@���;�`���Ջ�]RR���5��m:�.z`�F�n����7g�~�3�3��(��<�j�Jd�G�� E����*/A�ŕf����3�݉�Ñ��;1)x����o�1����Z��9Y��BYЋQ����ȒY�@�
	J%��5�,�
�Z��L-��&��᫂8.48A���@َxK��BժU����
���ϔ�b��b�f�JQv��)�7�z�O
�)ΐ��r�v�S�,Eb��-��%�.�#�`�%O�.Ų�,��őSh���L�i�3�pf�>E`��L0Rh·ע�yK��C�<��ZtM}	���'}X:Rq�p:�N۫�t��PKA`F����M�j��ױ��0@�(7UwN�J����$��{�z�ʧ/(��r�!�0��F�듲8M�����?��ϽUg˞���O�v�FE%v;3-=e��b7�A���dbm��S�f6��OZ˘۴��a�R��B-���T

��CT�GH����0)12��`;�����|s
���0����AW� <5�N�ִ��6�6�+����{��!�tu�a�b94d�>��f�bdK���'Kv
������;���Oʝm)p�~������2Ӷ
��6 ( 
��.f�D(T�Ftw�#��H�@VU�����	A���W�2/f��c�LbB,�TU�dq�3��pt�RI�m�/~K��6��0|RCH����`'�0j� ��frH��3�e�e�j�Τ���h�G-m���Bjk?O6�5��$�,�^��Cc�dcB��_��B��[��;�q�� hB���g��|��TU4�a���������e���6��G���I�H�$X��DL�#8%�b��0��a�hz���H��C<�y4K�j- �%5%�M�G�N�h���<]/�0�G������TDTIkU�Rp�ھ�*Ac���%է	��k���1�㫚�*�}��%@/-�85R+��Tu�۵�R	jdB4)^\*Pk�r�fP�s<����y34��2Y`"����p]�.2D� ��0��ID��G�
�U��B30����vW,��M9>D�'�[�J|]@6U{�f��'Ư��i�:���Z���h� g���yl?/�R��h��� L�I
|{l����t2��Q�(,����W5@Vﭗ�(!���`wh5J�6�$+;%�g�J�2�-�8��@V��;ޑ�47�z�"@Ȧo�{g����1Fgv�������!I�+��ҝ�*N�Z�QD�̇� ZR��uzp13��*UI�X +E�Rm�O0Ȉ@�<C�\H��T#���0Ys���D�M����%S�ǒ8D�<�D(�7'��R�=�uK�112o;��-���5����jZ��i�<8�4m�hZ��8�J�ad�n��D�"`u�m"�Rl`�M���W�0}�8�Lq�@J<� ���b�����`�@>|�@KB�lؒ�u��@F(5'm�Z�Y�O7�0�cU�Y }���0"��f�+�Ǵ����I��)E�'�Y�3KY�<��wv-��`q�\�$���n��	/+hkUiA���u��\�:N3(��/6!	����oz�!�u�ԝ񐲍!�.ÛGl ��ȥ�����!Ù3�/b)�&H\�i�MK. �&��)�%ȓ�S��rj8��ΤFt�!��}8�H��יd�2)�9��Z�x�}O���S��Rs�i�l����B8�+�^V0��N`��|:��ŝ�h���Y`��J�����,�Q���#H��4��#&�C���S@�,�u�!@f �!+� @)�S��H�7���n1dƨWUp��Z㤬o���]�c�eUUH���lG�f�d:��h�h�oŉ7�H�?jJp�(˪JJ�
���xKxχ�B��te#G��T�p:Y�3"<P��J^y��N�<N%4-��WHA���Y�\f*/���k<q�i�h�CS@Ak]p��7I�I֒���X�܏���)1&>�]��2B��E�R<+�<D	�BL���p���W.ON�޿��e����i�g1>d��rw{v�;���}�W���W�����������^��\�ն�߬��?��坷,�>��Q��\����pr����k�H�G7��[-�;/���"gb"�i���|�䫄�m�˙��UYb�s���;��O|���߽����óW�~M�_���s�~�ߒ�~��/o^��A����N��zE�p�??\]�=�>|z�/nJڭπ�Q����g�A0Igȣ1�䥔�Y'��Z��Zڣ,>�޽�����4x���� ����R/L��RS%���0�,�-#(���N�p |A'&��'B!��
YY��R�,��qa8Rn�!�5�ۦ��ӰYGD�c�w�R�LM�f-L�P�AI����N_9��)�-��4�'�ғ,>Y���W	���I
���55���ߋ�F�(����GH��t8fC6	��5���D�ӐDTa�&ըb8�Z�X!)��'�/N��p��G���T�����5�g���&)���₲飥?�
yȔ�Z~�M�����4�I�z&�$)��]#tb[�S{�bR���Sե�r�Z�(3gUp���%9�Ԥ����#�d���$��2�;G�@��`s�C�[K!2��d�ҥ�P������b܋�.��O��Od~��'?���½��%e��Q�̓�	m�����{�Xo�h�MA3i܆-��v�&5+�iG֒!3�mk)�� $E��XS�,;�������"�j[6�h�޵E�$b�HѺ�)w�<����R��$�#�������"�A��O��W�Fkc�w���{%�cڎ���q�Ԁ����;���,	�����,}dC�RR�(��?l�]��`f�2)o_mӜ����[��Ij!e	��0�t��?�8p�B��%�g��c��,�0P��h8��e�ȺX�#�[>�Ii$����l/�|�9p�����M�a��GKD����lY���R8bHjeG�����&��n���3�rʂ.(�M�kQ�X�-�bU�n6�Ī,yv���p�8�
SS����$��G����.��TR�.ʍD��+����m�J<x|yyp!#�j��7���Q���N�%>2�(�ϋ.������z�2�g|&0�z������\�Z4��px&��)�����    IDAT���1�־�!����g!��h�����8�� (aj����i�7-e��ڗؗ*O���
�� � ݉�
W�i�60B�tJ4��q��hir�iBG-M�u9]\)d�`��@�TR�y,��T.N�N���_7�e�hͦ~__Z&�c;��(��)K�m���Q6'�h�!�*	��c�kq�tMM�l�V���e��A�����%��Ա�����l՚�
���
G���gR�8b�(v�J��1�TH>ḙ�څr�z��Rn1�:0\w�� � >6�ڋ� �Z�5bӂ�%�a�
7�z(	,�����y8) !�8�@����0�s�@�?>�w� 1Fd^/�xm�l�@|d����E�����Iub��Ǭ]岍�7���z���r&D��I�NҷL9���Z����<��f�+4���t��jZdc���Tb��q��f���ґ��3c��G�N��h�8��ё"�f{I�x���@JܲZ�@:b��l!�l�`εH$���zCLyf[s<]A'�&x:���w9�|���|�@{���������++%���#cz��Y����.t�f��U%��U�^��~Rbj���#�/_�W"�.�ˀC��)�!XƟ%�]C�o{�aJ,5���U�Y
MϢ��$A�/͝���)5�h�gh����x1�F:>�sn3O��є�!T�m Ū��li0L�L������\w��J���|�i�*W%�P������w�-�h1�-����;���>�&ėqKRH��e� m��� ���*ׂ��	��-�$>�,\�R`��]A ���8�j-�p�,P�J Y��}��eÁ8b�ǵ�#{k8A����vjW"�4X���Y���(F�"�ɧ���Ui��v� ��ų�R!�;��uL�{	�v*�bF*Pв�!�CSk)?�LU��X:&I�c� ����L N� ^w���I	��6R��l�?1��~�H�W�#���R@��;Z}�����Ў����%?Ȕ%�/�����]&"��稦�ze{�p�8j�jq fc
�J�x�ٴ���&k�hhD�GLD���6�* �E6$^�R�XШ(���.�NO���<=��)��Ý�Nw���F��R���ݭ����_�@���ts��ܟ=���/s����pw�?{vr��9��׷�CT}z�/k��;?�ˇd�p}sw�[gr�p��J���ޟ��mV�Vî�e�m�������ML�]�W�7�^_�Y{pE�oo./�?��[ѯ޹��>Oo�Oo_����߼|����p���|}�F�_���}p�olޮG���ν��l��tw����X�==/u�0��i�w]���Oa%��R]  ����Ԏ&0Nc�����G �ḋ�!N���@��t*�-���̘uW�C����0݁�R�t�M��q�c-�6�ѿ|�Ň 􍁗;���?���*�^��X�u0cO��r�� ����g�f�)7�X��=0�b/�lcd�x�F��9���0�tBL^V9\-A��Z���R��8m��td�-~�5R8D�� �GG@��fD%ps"SvUT�`9
J����2�\\G����^0����¨��j�O�`�Re��/(� � c��,��ʦ�T����x�`Y�`Z�>5��9v/N::�W�Q���F'�UV�r:�NOU�MU�@_��g/���!��Ƨ�F��ƅ�7��!��M�@Y�����x�C*(3�b^k|>��yR��fp2��5d�׫�:��9�B�f�|�	}�P�xt#�������̧���fRTi��7E�|	q������-�
T�m�h�b�v+h$[`�
y��F4=�4�Wgh8v��p�b�Ƴ����k��U���0L������&Xj�-h�b���e��ej�n�x�]_4�Ԓ��.��aT����M���]#1}�C���C�10����ͪ���H�RUM}�&Q%0-��0���ݻ6�ܻ�%��Z*�d��APwA�|U�዁��LIVlwZk��nix�5���5�DS��mB��;&Ñŉ���r8�O�m3KA�!��#�.��D:��)W2Mi��==Fp�U�0B�L-Y�|%�[�ㅓ�$�-�N "��"S�����
���\UM��)�WK%� 3Y� �h��	đ�,ե䫭�X�.je�����B��~Rp��-�گ9S�I� �.hf��A�?ǥ�s��yF����씒�S[Cl6;J_wH��S�`����5�F�r�S�%&��G4Y|��CȚ�wc�. ��x�a�b"
�<��G3��/W,d)�@����6^�~���Ahr��+$�(@�g�9��O�����,���f�lwR�Q!bY�V_���fZ���ԙ��,iZ�P� BL-X�Ȧ�ݺ�G��4���(A�U�j�\JU�K���*�����2eY��Jx�(0)��Ȗ�;F�r�y��	��٩�N���k� Rj���2K],)G��J�j��V�g�&��!�SF�@y#�ǔT>$�ikh��*7�B�lGAD�O?A4� 8�q;`���2��]w�-13H����B��5�B�8�%���#�W�J�ҟe�8��f
G�	S��'��U:�b�m�6@��1C�p�%��ԅ5!/�B�-��~���,Ŭ�d1��1B�#���X��Τy҉����J
zNs_Y&�t7�i��6��u�Dm��š 9	yT���u$[!Ϫ�)"��]��03D�.I���������"�Ϝh�/u�B�q@�. :�)��40�f
��4� 3C"ʁ����(��B�
:Lq)���ʥ��8ͤ�HP`�r�
���RjyṶ�G�$�&�~K�xZLձ�,�8p��6F�����R�iˆ���x���pqK�!=#���$~�n�F��c� ��R�v��%_\	D	�dj-��J�!�T8�]�ÕX
�Lmׂ?��e�M�l
�O!2�И��`ik#i��Ek~dr3��|��g�;0�t��f���(N� O�av8�W�@Y��<��3�T;R���t4
�C���O>��"ę�ǈa���55� ��X �@)K��x:ֽ�f�Ya���-�G�`��t׷X
��MEH��ey1�����4�5�����?M)��@
�<� h;�l�Q�Vyqc@�M@��E������l���S��H�6�7�6M�h�G�T��вp �.�����4���)V�L-M�ZxM@�b���� �؝���cZH3 	F��X�i�00N�|M��)Y��f�8@K��Kgބ��HI�}��䎞u�h����,Ɋ����+x��|�Xy-z��C�f/8�$}�%Ah�j��A/�jA'�ie��
��
�#΢�xYUц���>1��DoQ�wN�.�l���=�V�w���{�߼�<߿�����~5��A}��/�]k_�-�{��'g�.���U���Ӽ�.}�r}�ӛ����~���A�s�=�ك_I�p�]��\������\?ӷ��m���m�[�]�1T�ھ�G8��y~��o�}��Ëg�����vo^������������������^�ϡ~���{���߿�F�7y��C|X=���6p]��o�&���.qS��y����%�U%h�շt�pTU/YU&�6��L>����&0LVJm�e3X@��wC�H6�NF�	)1Y�[õ#H��	�`Y�%~,U�y�x��C��w���QL��}�gD�DR���@%�b4��#�ϵ�S����-����{uJ�+�>M��X�����.]V8�r-4��	���k�����d��d�$#"�ԣ�����Դl��������r��L� ��?ܲ!K�� J\&���~�W�o���F�d�@���1apAU�֒g�*�ȲS���?� ���`�ゴ�߲��6m����i�HLK��B$�C�)�ŝ�Q�*�u�4e㴔r� 1:m`��*���h��x��dq i��iJ��"WՐ�
y`� N@���������0��s�.��	���%O����E�2�W[~���8��|�;��y��0!�Q����x357B��C�O�r�s�4�RJ�h�XS��A�l�=بgh|��	��
W^�d5j��m)���6�z*��w��K_�@oZ��0�oHM@��Q_4d�^��d�f�6*&�^��x~t�8D��3?��1e��B�֮����w��@��1;�1�yx4jް$δS�#k�X��Ԛn_�d��B^-D��e���#��
�H�c� f�ʍ�i,W<���Z�M�1�%��0��>/F��̦&7mUbU8�b^��j���-G�d�i��+�L
G���ņ	AD��!P��\J8r4�� �����-�1qf)v�� �Y��hh�F��#���� h�'�y�s��r��q�D@�IM,E��XK�1FN�&�� m�U��"O�^��=|<Z���1�x��!�L-2<�R���Nڸ� &�T˺�!=��=Q�)H���������҇[@��� H�2��c#hb�|�a���<?RU3�C��}�ݳ��
��$�F�Ȳ��iei�S�-5���\/"��Kim��D|���G�4�g]��m�`�����@�᫢��`�@M��pޒaJaz���N@V!�5�*>�C�G�R�EI''e��PK^J�ٺ��3D�����PȀ8Ū�L��0�S�D���u8(Y�txL�$
O��(h�RM�gr
��XF�;"��7^
<D���	a�*�@0�Fn�U��#+�*�J�j��@����#X�M�F�<��� =�T���X�0��Rd1�l�u��4pd�LZ-��LP_�^	B*L�*�@:�!r��jy��y8�g�8�>F*�^D���\R��d8�.�l��3}�o�i��l	��f��y�-k�7F)^�Q�,�~<	������Z�U�FH��Ĭ֫l�"��MU�����$) �/�˲@��!�E|��
�o�R����#4�q��Á'HY��[Rdu)�|39��I ul��e�I�Z�S�2��8��|`U��U��J��4p���Z-���28��c�gѪ�/}�84�*�A�o�H!�uQ��D�|���Gq�'8j�\_
8� �� ���(��Bˆ�ᖘY:b��n1�lj��$���s 3B}U��D��
�;��vQ*N"s	�?�T��@	>��H!8�q,V% �+��z 'R-~���N��o_]G���h��3)�r�$5�-�W#Yj�l��%D_�p4q���ؐɶ#)�\)����q�WU\m}�9��R�Rb#U(�[Y�.�h|��7	Z"��8��ex[
<AӖR��8�.�* �������.����ن��dU�8��@M G��I.�ͤ&;�����.�
�U�t�x�-TE�cw�	J*L3�!��C�e#5��Χ�y�O��	i0%b���8�t3%8^
YU�CJ��	IsNc
��G �Q3�rK`�����r��U�9:sAj��e-���dY�DB���+�;1�,��E����9Z3�y$��S��g�!m�.�&5�!PHS�U���S�~��U���0)F\
A��t$�Ƕ�8YL�If��id�-�%���0/E$�Q�o�}�?9���|���G/���Yz'��/]���_�oOή�!y�=�gׇ/<�z�i=�]�n/.�NW���w���޳ӛ�����g}���z�=�#�~5-�;����L�W���L���j�ǝ����{�6�{d���3���_r�-����n}j��̛����ki�~��?�>yzw��o���N��ݞ?�^F���y�w��p������}����y�_��!׻��]��[���T�6hr��Y�]lϐ���@� A��	@�u@�3���,5��.!ʉL��B��C ^�裏^��������#���to��8�T�b�?�Z��`�1�e��p^�]l��s�No�����cE^�Dp�=@j���G�G���E+�j$���,0)/�;@R��I�R��L��#��ug�qy��W�;��hZ�:[3(Ѩg�:&H�T�����t�@X[K�g��[pTU��d���	zzC4�4��lfdX�b�J138:������73��N�X`��`�@Έ�o�#@H?���� ���3_IK�b]�*�q�r<o��o� ������B��B#�v���>�FY	X��⎋�tEh6�9�;sD���ZG3�Y���8�0e�3���
tiS�6�x��-$��]���8��	����0���o�)y^�&��9��XY=�A���-��*�R�=^-߁6��W	,�O�d�	"ৌ)+��i!��\���!�:_qCv���%�w|jj�e4�d��ˬK�^�S-��M%�(d�3Rp�v=����N���E-q���u�1$ĜnJ����7��s��L���mM����g����f�>e�[D- ����l8K��aZ�����eK�1���q��!(��� -G\p\U/s�w^�1������@%bx��`Lm%���X6�b)U|�h��?���I��R5��R��	Rr6"��p�UM	B��~'ٍ'�WJA{O��@m3�����D�������:�nW1���D
xRoy�u�b��`i�F�9�L	P�Z�t9��ㅘ���Th;=!Ѐ8f�F�m�i�Q- 
�tx%8[�l� ~�����$|{�K!�裏~��zb�h��<94-�����4���Q=�-��ĺ{ʂo��H��+�������I��Vh$d�Z_�|X���uh��{�[KS��$�Y�++������t�կ~�����w4��$�Ϛ�]ډ�ubZ'��l',�Ѵ��uN�y��L���	���������o�ij���Gvh�|}��&T"+���}Up�8X�����������Z`�J�����2����A������ǁ�-��p&��sk�!@p &�$�����8�/0��UA���Dfm��}�Z��OD�%��f�gԥ�=��2M־�b-р8D̓e�ѱ��k:B�`���i�B���/���q4q��B3�e��苑łڅ���,��ނʇf91����ɲ&��RUm���<���F�x�	��lH��QF��8��A�o"b�,�)�pJYN��Ԣ���$���NFG"�7RIclH8á/P�p<?�,�_R�@��y �d)�L�ZHd�Ѥ,#����*>/�P����)+Id
o)hDS̻�J�GRX/;��S�<q�֮�!1G���@}1GY,e$H�s�����@ҡ����"F����jT���f�,�h�OA6/�����ӄ�TwNC�q3IAy�uC�.fpV0�B�J
�y�Y� \/�jb��jimj��>~C»()��mS�UQ�(ӗU.%��Yv�	��"J�Y4���剥S�j�A�jT��4R�����u�LU�	
���]�}kQ-��S����]�zż�������4�Q@�<�~:J4����<P�GP�8�8s42I�4�X-��`q�v��,_d&��m��
��K�e~�_w,�����Ԯ,��9A��8]/�qk[��ܐD0j�7F%�h�ײS@��$@U͐Z�թf#�˚$q�D�H���v|
�!�����	Gc��m�-��bZbZ�:BdŘ��3�j�J\�tO0���"�,�Fd+OJ��-egkR3[ʩ!��j����@F9�l�1�R=֪j$�^�Y�(ıٍ�������h��3��ɧ�x㕐b6�V�`�o�0��ڋUIY��&�.b�H�y<2K:M+�i �����G����H_�z��~�u�^*�'��2#���KS�������N�8�g�mؐ�ٖ�5��q�ߕ�.m����;������_��?sy�89���___������z���-o��̳U����|������������ğ�t�_�����>vy�xXO��^{H�@�?�>��~�����9��bSxx{�]2�    IDAT#��s��?�x��m����N�u�>����@|�;~��u_��w_ܟ�?�ͳ�W�4^�/�Wv�s�����g/�}�����{wvy����׷�k�X��`�s(Ev�O#��(�[߮Ї�eW��+�{�,OǨ1��
���_^J�5�vM� ظ�/�㸝��D��ů���ծ��xj�[&����K1_I}+<&��U�&gR#���+?t�b�^т���Y�d�B����ᙾ���Mʋin&���̤�'�C�H�}O�1���[����͉���~��T��3�f��P�Nbk�hf ��J���3�{	S���V����e��ehb}՚��$��d����������cIYֱ	�M�������MK� �?0�R�U}U�ڷȖ!3�..eY;��ۯ��@��6tE �m�<���vp�X��M����,5���q��рZw�	*1!1��]"�1ņ�5��
�FƩ����23 �h�d���L�s3-��K�}�я��_�����<�ܽ��;b�x���S��r�!j,kcyScm" �M�lm���J��A8��2��k����)A�#�4�]u7�R�&A�
eC�(��Z�wv
]�ްc��ΡB�)�RhB����ހϞ�7#���w=�40��:�4��(Y"�����B`�'�~Gǳ>��"���A$�Yw���9�,Y���\����}L�i�/H�!P��@)F�B�v4^�.
�
T�3Ӣ�7OX�8��g��Q� ��<uX1�KUb�0Hq"8@�LL|Db����,�V���$���]y����ֽ�H���̬̈���p�-N�������Ux6��'@BB���š������cD��?�pۄ��-[f���Y���-��![
�ۗSJd۔f�	�La4U���e����l8𤈨�&���1^�z _;�5�'��	�j$֨=�n���B`�WKm��ִ�Ҭ]}ӯ���1qR�R���@QeL8�T���B^�ND�hj� jy�i�Bc�ʳ Z�zY"��!&�]��׬�8�����: �8:�|��4��Ŧ˚$P Ĥ�3c+�;g����)�pY)Sx*���5M���Q=�̬�F0��>��\��&4�/o��"�rMڣ�A�"Sf,Ӝ��>�h���Y�,\m��# 3q�m�Z���� ey)���0�1Z�(b���Z�k��� �gҎj`VB�W.��IJ�@-XW��K� ǯ�`	��8��dh��Ȝ,N-�����,	��\IU��(�S�m�ɥ�S�M#���∕L���.1	Z��t�ʢ)�0HY��i+A(+��▘,Iձ-�F�F���F#%t݇�-�&}j5�Cjm9j�F� 6�
�A�1IY�%��jm$D���YnՌ�Կ�L�\a��F*HgN2�he���xd��;��%K�GV:�6
�v!@�W){l���R��N���&V������պ�h�d���95d&�h�$�SH�8~H�T(nC}}�$}�A
J�NR�I����v8� �.�ΧS�eM�}
�8Mh)�k��eME�K��d�X��(�,��+�TK%�|�r����iw�Q��!0�Z���!����+d��:��3:Rx�b�-.H��M/Kq]�2���v�u�;U'fI�W��a�̀P�Z[�D�/��z�S�[&.�G� ��P�9@K��rdK_�*� ��0��L��-5�I���m�в�f�`��B_�q��ěs%��H��4�fS&�2N{GC�፧���N����|����9����}^J��헵���-��M��^p�p�@6���\���ץ�n����*<r�_���J��ږ�&)혥v��Ԇ[6� ZH��ґe��VՅ3�-$��B3���vY-&!��5��`-�Q�<e)���/�J0&B�j�34Y^
�a�Z
�I��A��y����u�-�w�Ʃ;P���b��Fa���̽޺�Y_w��JAw�DD��76��+h)�<��E�P� �Z�|K�Q�ҩ��mVR�H�mɏȔ�#0�Ϝ�B_I-�:���k�LaALKWR�-Hi��M)^ܵN�.�`*�[�tx
|�]k��Oi�T'�N{�%���S�.��
дn�.�e��QP+����-��L־ڎ*���1�)�5�I�x�
*|<�j�L?���ú7������G�>XD�<���O�=햯5��6��>���t�������7_�]?����xv��F�N��|z���/�|����/�=]|<�3����_;W\_�}��)΅����/�]���'��zo��{z���΂[�\�ݝ߹�]��z�ݢ��]�(�������=�;�����k�ǗWw_��×?8ݼwy�t|�?��}q]������^yvmˬ��d��� R�V�j
Y� � �3�nw�h����Z '�ӕ��.o�V�)��F
��4��-�	�$`eՊӄ� �t''Gc���adŐ
��x��)u�C�1�'}Ui$۲�I,M�-���^#|�
��T�k�� �c:�NRL��K��R���* M.��q����@�K KG	�G�ׄ
y"8�e�WD&"�R+�X��>�Y�A����(��]�����x��
u��HDU���?뎀��@J`x�G��?���x"�y]0[�b��b#MJ��,�ᔂ�A�9��&�mi@�Ri�k2}��,\k���l�~f���m
����87v"s�:d�9ժ0)����t��s��rΘ�����4 ܐpKLY`�J,�ˁ��c�:��(x��)�*�R�Q�>���_�jBF���ӟ����?���g"����u>n$�-��j�EhX�i�,��Lݬ
��)shV�J`2�qU̖<�;��:G|�@������I�{���4�M1o��R��(�#H��)#0'B_ (��Mv��>�� �!(�ڒ׽	ќ��1��a�}���&�"Ƿ�닦J9_l A��v̮=����FyHӢ�N�������F8�Z4��ۯ��H�Q�h4�J萅��N�m"�?��hJ�Z�dd�_̐y��S��F�bN��K��Ϊ��� 33�r�0!��J� ӥ9���E�jqh*I|;�M!(/%pEx��y�bL��M��p�Ƭ]�<Ș!��/K������eM�`-g�Rh��]}d�QK"h��x���鮶y�c�!Db"h*+U#KA�Ȕ���f�cL�^b4�r����&�3�B&VU���)����EC"�ƇG�dR�Ԗ룟�I��bLj)Ǳ����SC�z�K�5n0��o�u�e=�kJ�N�s	� ���#Ł0]L��79N�Z����ƇXz��XzQ{��
�����Y�lwTjs>�-�y��#�q��:�����L.�����
��%d5��p0�7FJA☤Z�t�	�$�%�D�����81�|��:ľ�ۦ���T��H��r��λ��!�B�}��cB��s��������N�Z����*K�� �0
��W�g�f�Q;����?�6���*H����0�D�S� ���<2N٦j�ZWM quFç d��r�d�i���5X��	;s)��V<}S�d4��__>��q�ӡUųZ� ���Kє�䁝RSDVep&e��Z4�l��%M�^��0"�Բ ��L3� )�͖�������*F_�F��������6�.R��	X��� �G��k'�0�e�,;�%k�A`@���N_�?NH׮��ʉ	,��R�!J��{ѐ	�L�U��n*�r��WB"��%��f](h
2q�J,I�AR��Ek��ķw��5��"�"qK�,�G ����R����9�-�d��=��F0]*LJ�!�ZfuĴL?A0
f3`���b	wh1�$&�Y�OS*�v��
����9C
�z��b�_9¤�-K�.��YJ)/h�f~��W�3U�5�4�\���~�jM���5Iy��^�,ĩ�b�]j�|�g|qw_�UY��!5K)�v-|�	Rk���(,W��<��{NN?����1�e��#U�Ԉl��B�H�*π��DFȗU�f�QȊQhI�3�e)��u���hh
�]�#����B����ǁ$�)�CR�G*5)L����}u}2�"�t��G_�c�j!��WVU]��^q����h�ܦԦ&��6�Мe�"hMXw���,�����Lw�0�����^l$K 0Sۉu�IM��;�pR8N&BRI󫂳I�5���*h�@
�Z
d!	�&k�J���?���)gz����k)N
�BqY��2xA|������3��Ɨ��T�+n�"��8m�uQ�k\���l-�mY��pFj韜&2��lU���!�;L�e4}}�7���9��G���@�_�RވkB��j��X)]XC�b�vwj�Cfs�
��4Id|��l�O0�g/?oy�,�>��ڼY>����������B�Å������=p�no.�W��6��*}�;ݟ�������|�����'��؏�?�;��|y��/��{}��?���x�_�~J��d��oa��~�,����O���-������:���7ޫ:\�s���aip���wˏ��/�	���7'����_?>(�?�wuܿ�3��{�_~�Ë�pzq���?oO�o�����v��W�I����\9(���9�b���Z�H���������A��z�u�uc�����z��"ԅ�zk<z�D��iq/���T�BR@�i�)�	�VU�p�9���Y�QX*T5c^�B-����xuxk�s@�����,�v�[�Z3o|97��G֝���++��y�����T��GҳB��L"`Jd��1�!�{�(���Y�����Q���םH�e0`k��x�:��s#ː��7���hG����	�YJ�E1���Q(!H�UP�V\-Ħ��dD\�5�y��	Fk��<e�Z4��e�!���T�X2��`�S��XV_��W"��8��CJy�;����@v�c="K��u�h�L"
� �䵆 �% �tQ�MRw�n�h�]qDI��rUR)�+;^�f � ݓ�)���{۲F�� @33�tKx;�w�a���b_��}�`�������������D�����o~���ҤE<�4���f��L�&h��+��mt��"ź�.-&��A�Ԋq����X�ב7�R
��T�pT�Vl
�f��K@���S�����jLG`����~�;���z���s�D��+�K�g�#B̖�BqWר.���hڬ��j:%%��dq�R	1F����E�ӹA�3��{�汔�޺�F�կ��,&KJG
�n	��ru��;~����ʻFZ����vHDL˪d�8�O�@��D����1|�`J��/6@L�zY��^#�
�a���VJw�Ù^�ӧ9�(�i$���>�r�3�^��pj����.��@	Y�SPӖ�F�F����1ŉ@�$<�)aբ�_����	�Ɣ�qRۑe��Y�8� ^.Gq4��e�)!XJ�Z48��YU�p���pAM�l�X��c�ki�����k�̾Z�/�ƶ�'���C)2����-���ͩ��0Ox�"h��_%������ G!}��;w�Z�r���r�@q�bS���~���?��c�v��$�|�	4f�|ݑS6� A�����8�5������Q;� GjR�����6����Q���<���}����ɺ"���1y�.�A�n�
]n"@[��j�+���":U��#��u�b�F&A�Ĳl�BK�(���FU[s������ے�1R�l���Fu�b��yUņ�[*q����?��o |���BmW���i��7��-!ΚA����01��� h!?`��
��X�F ���;R!_�����H�1{����#�Ph/�4����Y#q�ӝ�XJ-S� ���#.�R�o<�R�u��"7!f1�=�*ox���5C�Ť��*��l�RS�Z{L�g� _V03K� Z�
����[z�*T%�yИ��0��AT�\��@����bYO�lo9���/[!N-,�l85�w�H!�3�Zc��JdӬd����X4A")���M��
@��	����Ԩ���Z޾:s�Ȥ��.��K�2��0����5Ň��0��R��U��kٲ-��cRD�("���d;�8p�hRD�XM����b�nN��Rq�L��9q�U�I!����9�L�^D����8k3Z�f�Y[HS��-�������4��
-x�Yn��Y���n�D�p˱����(�_�����t!�F���*��� )X�4U:�o%΁g�!���фcr5��c3Я6�g�*��ͦ0��e[�PRI���[�����˷�L�r��AR�� 7 0��!J�#o�R�(�hqlV�e{�X���i|�����������!�����Z��,�_m��HE��4���;g��@]���<ek�&`��F�B^	B���Z+)��W�Y�Xv4,]YK���o�SH�BA'�!Se	LM ��3�(W�r�TB
S�T�<��pL6�d�K!��a�"$�ǁח������r>!�;�`x�9��Ưr�r>S+�U-s�9@K�Y΄�^�'���Rh���ZH�����1�j#� N\�B�������D��	=�d����`�����Z*d	�*�7a�@� ����.p}Cj���{>v�+Z�}f�_��u�N�j��������e��>��N��w�xw���5�����_Q�t��b^v~���K=.����|z��9��~���u��݅���_�n?�y�oz.��^x��58<��Qͣ��9]�T�с�8�U�.����r�Ћ����^^O��Av�s�/n�7�Ʀ�i}{��S���\�������ӕڼ����v��/�:\=�.�S��s��{8��O��Oo����u�.����q�Jd�>��0 �^M˥���_����ɣ�_#�*{���r�͠�r5�t�>���G�� �*���m�1��W�U5{�.2�<M��<������(@X�:����jx(�F�!�;A�W��o��Ȩ����N�%)�G!_�J�X_�� _L��w]�o9���D�#���i� #����-�Y�2��b
��Z|�NR�	��_w3'�V@�geO��Xʳ�R_%�,F;x[�bͯV	Y���@�{е��_��b�k�]'���*~�[Z%2o_<%��KMa�[K��X w&�:54.�W���J�PK�=Wy�G�wz0�Ղ:䪤 ₲��0�6�W
��y�)��l���U1dY�����sAS�W-�&�D$�^�эAD�%)��_����ʴ�B������9گ~�+~نǜ/�T��S'�Pw?	��ﮁ�U%`
���Z�8�·={P�Tb�e�L
!NA!�� �i�$�|ͦ�F�m�.d� T�����dLH͑��K��2�X��tt`��mH:���7g�<����2�9��F�8�BͅdZth�iR�����គ�?��Aj=|%p"�A�Z@���$��ah~�k_GP�(h��eR@����]��7'|RS	$X�uHU)��dR�!�B �#7�s0yKA9C�M�fA
|�VJa�� R-��q��&�l$�1�-K$.&8�� �,�*
���WU��+��"�b�b>��gpMk� ��jv����e��4$�Y@3>MK68��vI6<�v'l<qc(�v�]ԑ�$�c7�9٦��*[CH?�X*N��H��{1��2�X;�t���� è�j�K"���/M)�b��W�3���$Oj��������$+�Y�o�Z����ʘ��(����0��̂J��n�R-� �6�j�G��K�ȒRE����c�V�#؂l��
�'�`���*䩡ե�'<�rF��4)�,�����59NY��|�7��71
�,/6��%�%�3�Wp"��/�ifU�B�E0sc �j������
h,5;R[�t]��n.    IDAT0�&%n>Ȓ�/�
/����*1a"��� �l6��5$���׽ֲ�Q�%K�FZ�DÁ�+�/`�#�%�J�<)�y��
����n L
��bq��Ƥ�a�!p�p��0|R�RnK|�H��*NY�.�94w�hij��Sw��6.��T1L���g��r+%Nd
u�d�i��S���B�Gk�|"��\MU]�O@Δ�!L�HM/`LA�Df�@&frd��	�#�y:7KdMעgg����^ȝ��Ԓ�Y�Ʒ��Q��)��g�7f%�lk�:*�1�YF\P	N����.G ��Ln�F�J��:;J�f~4j��T[��-�� a����94q���nc�h��8���69)N)��t����Y���EG��)dD(�
"�3��LY�8�l$�L��#�5��m8�M���U�5�A$[���X� KYJ�(th���J5�別�Ҵ�u��ܴ���T4L%1��<<$�Ė���d��1y�6%�Z��r%��Zڦ��8S.���u��e��:1Yje!�83@N
�uxL1�X��x�f������R0]�
g)��FA�~uA��Ѝ� �#�#f�@FG��v��ƛv�,��H)�5j�l^U�!K��4�����1�%UI�р]��4�Ap�w���Ty�8[Sn��N_�[o�|Ub`RFB,�d^�SRЎ�q]�'|J�m#���X�'@c����r�nZH�KlZ1�O���iY!��ͳh���#P�_�M"K5g��VG`�JUa8e#,*�))d8!Z��#��&a�kY����T�D�l��'��Q@��.v]�{���_���R#b)%<�C�"�+�F����@d>C��
,��G���E�iT�b��Z��)�)�ΤC����p��ia�{�����Q�4O}lЮ��Z*>� �ljqL���_��tr �)=>����hl����w^\��N�M����� �?ryy��:�=�������-Ix��j9	���χ�s�tqpbF�����J����Q>�!K��K��W����ox��y�_���H}*yu����[!\S�tT���ώ����D|���?��h�?�l�o�<,�q���tw���}yx}����������������3gw�����������gE^��.X��u��<�����4�,&?W�K�cV���U�iʎ��*q�_���񡦥����S���� M�O_�q7���7^ی/7�rU!q�^)���&X����{�-1���q��6ޣ����?���?Ѩ�|�{�"Y����y{!��3�T�A�HY���1j'% "��q��A0��%?s��e�k��
i��-1�<�ʉ�c6�;
�RhNo�u�uU񤤐�W`iN���舑yQe�<0#�l!,�e��-Gp���]G����-�Z�ϧ�F��	�/sl��k����^�꺯ZD�ve�
�5�Y�#�磹]nK7��k���	T�l��s��N{��6}1Y�F��ײl|��' �Ժ�M�ɫ©|t
xYVwK�&�>ВT�1e��m3"�}Wh<:��9%�xkכ�n��g7�
:oH��Aw�����}Q�7������Cu=:�v���V �j'�&fD��Mo2
�h����q��-��31�����ڪm�l�s�t:;�*����e8�� c�!�'hB1o;Ƚ܍�������
�B'�	���p�.L���*����U��ź�x�� s�\H �JĲ>�ŤRV�� K�JM�e7�XSw�6�]ڂ�X����� )�o��q�Kaf&k_����b��[
ⓒB�,%X���iT����c�o#bd��	6��d���tO���^d-�o�%(֮�	�!��$ß�C��m�d�_�e�.��	�֗Ǆ�%1N���N�>�o)q32��6+��c:�}���y��	�B.��e�Ș�B�)qAGsj눣6q� �
x��o�(C�'�JYP�p޲��g�5ؔcJ�ߨ��+a"��OAmWG�UnZ_$,�� !��XJ�W�k����N��2&AJ�2}�8n�""%��<!��uRb���:����U�)��zQ�h6_�>��߻��/"Ph���0��u��ɚSʲ�e;B�BLJ��Z�RnZYw�pfY՚Y6咩�^/�oӥ���/�	�/+��-TBӒ5 Ϥ\5�����릗x����HPm�8j�H!0��t���gm��ׂO�o�[&��6)%ěs;C�
�q�XG����k�I��NCy12���!��!�TR;jDTűT3�6�$|�B��W��4x�T�<N��d1�N����O����#1�<}4���S"�`�Z����r&��]R-yC�kqA���P>]*I|A�R�9�L����Ë8r��i��&�@GHvbA�) �.�����©{� -��(R��C�^5��TE�c
ꅆCM�2��ʢy�6X�fC��oY;YH�jQ�3�N��vF�Bj�V��lb��qB� ��g��T��4O�)`dH�ƈY�h��h��H�Z�R�-�Z)�S-A3 �ѨZ��p2x ��QP�rqx��iq�Mg��b��F�� N3N�p�3|K��V2YNYg2#����&�ި$�hź04')�l $�SՅ�$�a����2�k6j!h�Zze-���F�
=�V�����jH%�^�X/ҶO��]�<���3 3/E��R5�������dx��]��P��4�TE�X�! �@[k�{
b��wV��!�Աm�-YF*&�5� ���o�b�5J6)��U�ٮ�vYd�I� a��HӔmk�8�D�/�M��gSRZ(d�j����,�Z�a�]��|[��bx��U�lkM�o���5UXmUţ�F��µ�CD�8Y8'.F��k��aR��2�v���������`��,˪e���M!s><0S(HM0�qR�w�S�j�zs��A�d۝؍G
�����2Yq�@���S9)�%B��J��D�i�L�XֺK�Hp[e��Q)�n��}�{~��/~�_��ף\P/%3����6.`J�����3��I����+8�QxD��R�ֱ֖�=��=O��z_N�a��e6)�J���=3Ų�׋���n��4
h�� B����lq�R�Bp��u���t��xyX6~��J/ًk����q����_�ڧO����^���Y}�oj������;W�/���./}V�����q������~�r���P�����O^^xx�~t��u{-'�|ֹl�$���#Z���N�_g{���[�������6w����p|��s�>�=�?���?��>}:�O���t�{�G�������ڤ���j�w�7/����=�]]��g��o�Y��u�����6H����B��A4
K��ޒ�,��@6� ���o��?��+_������U�-�x������|c��L_�&�Y�I��+A��1䢲��S��ŵ�xD��;R|�<�׻L�,���zy/]��7�eMEs�G�oIVl�� 1�d��Ad)dY��c�l_hp|�zo�[�z�!M�o�)���iJ�Bg8�Z +/h*�u��,Céc�b�R��U1Dk��B8e�*��~�E�m鷾%��Y�˄I��a�GA�tZ����f.[
26�Rb�[)6`4. ���5Uj�CxKxAUCP8���汬P��:�\&A-���uD�
�,���Μ2Z�H ��I\6>�Q��,
��R���+��ă�q
�ŧ��!gZ��1Y���֭��<��#x!���m�����kܻ�LS��=��c\^�
�읗�N���:9����ǟh�c5D \o)�fB�X�Z�Z�]���cT%R�΢��l�N${3�]- �n352��\b���E7rx����o=k�1LjS.���u�+}�� +Wk�����b����� bx�P��y��.eI�Z�w�ޯw��8e[�0���z^�@��/f<>0���i f��4uߘн������~4��*���+bI�c��Z�uK�7_���*�B�jq��2��}��>-�����6����hi��'�H�� 5@ʿ]�)c0)%S�x�x8�F�R � %h!4�B���F�dp]�"���,�N���Y#�#l�!R��.�d!� (�5����`����ܒ�AM�}e=��M��l���
`+,���9��g�f�bh��T�t,i��)��4[YKL�E+Y�x��>%MH�ˊ �C�F��pƐJ��р,)A�y-,��0"qh��Iyz{]#��=�
�BG��Hj���O
�������� ��DU�� A�3�e�8��bTH�<�>��#^	D��4=�t��O��+e	7o�N�R43S�Z��Ix���%5��!�+���0s�)hY 7@%+k�i-Ӂ�H�U��Yt>Ȇ����d��@�����t��@GGGǮ�m"P�X��kM��h�L\,�I�56O��#��-��Hj�Bz��9K1�u>Me�V,"L/�}-�)T�R��"c��씔HKY2��R�f�B��NA�F�R�txH��]h��"є׽F��V	�V��%C���	��0��h�wD����TH��o��	+c�.+gq�
�.5����:�R�TGQyL�^e��2�;m�2|d�͌���cZ��mI�Ө
�k�IA���3
LY3 �$dp�F�o�#��,��-{E[�YR�+��R�й���$2���fHs���
̣e���Hܐ��� _-��MA�I��u�#�&F�)�%����oG����5��z~�4	\���^��[j$;R��״��f���R��T��p �@^�"@�B���-D���Z���ݶ�M�'����h�l�K`٨�=Z�x���9�)�l7��YF"�/�"K��l e�ȥ j����uW8�8@�JD� D,�)��rL^�����WkZ�� 8d)��)��T�Vy�H���w��0~y"���%<N�B�T��B���$��p�_�S�Z�����h�~7Is6$�4)0��j�ec����Mв��[���|�ј	��ف �׷^��$��Y5F���c2��K�������cA(F����i{zT� ˾1n~��n�jg_�d�a�	޼�+�\��t��T������(}�b%�-�TL|�J-���[���@����nI���g���B! �vx_ V�A�Xs
�@����C	N�Y�_����G �<Bd
�"��;�)oL8r��̊�X� �#�sn���2�)�ʛ��HS��$`K��㴋/EM_^cz��ys�����f���u3���@LY��|R����C�C@,�E$N�/��P,`���i�S�9�R�=Ԃgd:�p��l)�mY�+��w4�
���A�͆o��8d�ޟTHGSF���#������t8�������/�]�i��6��N�p�̞=R|8x���o����>���ٟ�<���vt��<�Ag�/�{|����'���_�ܞ��m�ㅡ�~��/�]�~���t<]X���w�� ��A��������~'�qw��yk�>5������'����7������"�yi�������t��u�,��r������/>?=���^�wwxqs���{�}uw�U��o��>��E���� �2��zW����$�a�RŖ�.�A�{�ll}E�Y��7o��"v!B�������G}d��-A��&�$D���3[�/�f�{��jg�T��*���%K9�6.OMG�i+�jB#{oʋE`�q\ޯP�-zcXz�D��p���Q�;x)�ŝ^���SSn��y�^�<��d1�1 ��r�pj!�
����g��,�.J J\lNc;���ӻC�*4�R�!��R؝ �fZ:|���r���/%�]bo�y���0�u�I�FP aR��C��-͒a⭎,�VG�@Z�� �J�|�tb�a��;C���m�1�nH������r�C��J����w�4�����!u�6^*D�8]��"0�6�0"�BLxR�@��aY�
U�����8
̹�p:;���x�[E/�_���&��^����8~o�썴�<���<� nMfr�H�f��U�&]H���&��3Y�B���}j��lӷYG�+L
�i���eb���t4d���t�8ƈ7IY"b�2f��+/�S0�w��5���O��_~��߮��tQ�öj�ʗ���x�|���s2F�CD'L���Gs�4>Z��{w��7C�u��h���ܕ��tt���O	oɷ5�v�{��I콱i���迏s,ƫ/\� ������J.�`��lxKxUb) dKv��Ʈ�B{GF��Ĥ"���q訂8�-�Y� Y#���0R#wz84�)���r�JhVeYS~������IŷĄ��-�i~��� f�k�+��)�T�ֲ.���l�
�rV�S �k] ��j0HY|:��j�T��E�]l*�uSU�	A�:Z6̶����[�d�h�!զ��"b/HU����M%&�P�l��Sm�uA�t# �ԓXw��ү
����д�
� ����ic;�E͏����FRrO0�h���	��*���sF�G�`�����~uv3WE�s�O�����LKӲ SIç`SYSy�0|[�(3��!pK|ޒ́�����������I�*��E�CJy1r��˶G����e�e'�a�C�w���f�)�o"��o\:��d����8p�Aj��j�I1�3A#2��UI��V����7j���3�ZKY)R��H1�TM^�Jy~*B*D#�L�L���L8�A�Z'ߖ)C� ۔�e
���a.B#��D`���ʲrL�r)}���A*�T%�D� ̦�0 ��7�`��m��i؈`�X->)�vb	�K��(֫Z%��^�8Mb�.%bY��W�ֺM5'L��1_�b>溏�/%%�3�4�lU�!���Ѳ��e#��W�j�v�>)L���L�7F"���T�ڥ�F q�(�0R��x��	My�P|�eӤ�����q���,>~`%�u�e�KY�3/ƤY�c,N$f
��D������j�!�j�A���&,;>B��Dp5={gS��q�Y�qH)��|��9��~RJĲ�y1����#RU!^-d�Dd��R�]w%@H�Ul6 ��I	��"�;@xZR��,�$�;��^*2��RƏ�)�N٭�8���Ӏ[���Jc�;+`q8��2�斀�R��ey rM�b���cꅬ�u�R�Z[*��Z���R��Q,(���b��G�s(��&��s8+�|�&���'����)DJ\���l)e�b�HG|1�D"���À��E�%�ձF���e�-�V�~�R�5�*8��	�Cj�D ��e/��N23�o�m�f���Y�� �&s�3!� hp���T-�A,��<�f�CA-��u�K��w�ZqK:�� � �5
ᔽ�+LP��
 RK�����4#���Zfh����֖өJ,`�6B� �����8/��i� l��"�E+�J>k:�^>,�lM�
����b����!�b-ĝ^�B������sޠ�.��S�`iSJ,�8�F<�ZYR�ΡWNjV \�����.�!��җ�Z����~�kaG��T�,e��59&�؂�+f@�]��'�����!�_vā|
y������ ��|�����������a�b�!N�Еwu|��G�Nw�~Z�����p��Y߻�|�����Ǘ/n���/���5Ƀ��ӟ__��??._1�_��_-�|�y�Kew�ˣ�-��̽�U�|���+m��Y��x�t���RM��Ǟ�*�5�������ɏi^��>��Q�ϑ��r|���t~�s�g/t�S��Ë�?��0Ƨ����O��������Lo��g���_o������O>sZ�cq\�qV*s���$�����Q��Zt��b^j�ĝt��L���f��K3�,K�9�y8�v�Q��b��,}K��l~`
[_yç��r@�����k?����_v8)ة7�Ľ1ew�2%���8�hԦ�1�y��    IDAT�FB�_�Z�O{��5Mk7�B��w��&�,�r3�0�x7Ƌw�вq��O�x��S��n*�fN�� ���^�,B�Z"Ї�Rk�J�U��f�0K��)�$F�T���b�d���mP�\LǓ��"J���o��C�rӥ��%��8���x�6��r�lK��TE�5PV�eAN��N@�J͜�Yv�͵s���Ah�v�霻%�w�d;:���+��f:
d�,�@k��r�����v��kBL����Fp���0T��R��^b��7w����Iz#�Qx7�`}�B��7���|Gw�/�1H�:ot8iG�Ȩ�l�[�z�PS��ͧ���m@����~T��#�hڧX/�@��AX��핏�2���g�p�4]H3`�8y�l�`�c�kai��i ��+l dA�nT}����������S-5�����{(�*�r�r�������)`IP��k�G-}ӃL�k�.(� ��x���"�<.��K�ޢ��o~S��v�Vś$�V�Kg%�̀qA���Q��l`�Ro)�Ye����p� "���I�w��B�j¶0���Vk��J	B��j�j� ��SV(�M���-)44���6��B�x%q꨻S���tt�1�#�EL �^"pF'�-S��.h01SbY��Qۂ�jyx��<k��#��A�f�Y�#��Y�,��לR�hs ����!��W��2�*�d�Ԇ&кQ��Ī�V��K�׻�$�<����0�wY"�=��/����NG-��^	JQХr��fO<�Ų!=e=��z4QPH�cG�W&#y���=g|�C��?����󕈃�裏>��c|�k� �f��l6�朣#"�UIi!��jj����L����T����(�
hJa6!�6�m�8���)4F��/"(�+Q+���42!o����rЦi�D÷�G�i��.�%�)@V��aX"�R:J��� 
��\!+ȣ��lMՆk�B���������ע�-x:y�-��	���<yV��+L��3��b6@
#+�3-&U�Ϥ���bN��o)p?(� 0@)H;M��R���h.YK)k��tR�*K!8^ʲi���Nv�~����.qCv���)ʖL���BY�c*Hq3 e��G�F]2%��^yj�p�M�l-(t��v"� ��)fhd�I�Ra������å&�;XM�Ul�r��N!o��C��H��3i�p�F�<����<B�h��4/�%��:��a���Ԓ�����jַ�Sp�+'�Z
d�+�T�)�yj▕�lK�2܄b�t��<\�vJ�$�z)l0|H��t�L�mVR9~��<���h�ɇ1��-���0�psZ�Ddq0� q��vTj���OkA1��S���`���hB��'}D<2/%8`SQ~��u�hu�B��2`3��3�����ڶWq��H�P>�ȍd�;1�T��Y���X63_-fH)�ત�I��jA�2��V�|� -fA�R�r8_/A�uL!�,� k�}rq-�Ҭ��N7d�D�#��U�钦��Z��^���$�,��v�v��t�8����H��H��) �{%@����Re{��n�e;y-�MU	�@	��&�Ȋ��j��,�J��4 KGJ�Tk��㈙��A�,��ǟ*�p�u O�f��Z�3�v�&bN,@N��mk!u�l�),�`Rj�L�0|�#���t�`�GkZ�rx���q��MKY8K���8��K\-�����h���g`�"G &"IV�R�������7���~ ��O~�P�K���BYG�,ӜM�Z�v8b
����+O��XV퀤�<��A��!��%����1M�_�����h����T��|x%����q��W9)>CcJ(��QFV��3���֥���K��A�v�'�~�)�_?ܿ�r���~���������OT����I���7}����~~�f}��ɟ�y8�ޝ>{}���;�}�1?sy�p �����#�����+�ӥ���v,�|���4�'��Kk��#�����(�����K�C��7оxq�p}8/�|t�w�.O'U��ؽ��v��x���������Z�.�~7������xy��ݿ�����ţ?�yye�'?��c.�rA	:�N�I�ؐ�'��<�,��/��!!ż���K���ǻ�y`�ˉ��phpU�@�������X�jL��,�|K~���� Y�B]Sy-u�b�⚮�k��B*o)n<K4�8��3w ����~�G �~��-�{O�ީz[�I�J�ZF�$�d]#���J:綀�K����������B�ZG�4���t5d��P�aZ�틧i������!�[����tb�VaH��@(0 �������T��kkffjud�XG۱�a��� ~F8|�L��I,1ٚy��%��<���e�����dq�i�P (��b>�Y�8�<�}�*#4!�uC:�R�6"�F`:L^��O��wt����;��A-A��|�1!q�!@b[J��]zY�,�f �&�&�U[!MA�T�&A�NC�X֍�$@|
}���W������?"×{�b����;x����"s�ڸ�U�(0u����^�(ˆ�؏B̇dD��j_mUƀ��T"���
Y�v[U�[
AV�`�k��¢���j���b���4�x��� 2ܾL��N}��f���Y��+��L��	Bl��G�㨼*4�e7�G�v>�@6�K)�a׮*��%>%D���zQH�3�c⿪蟲>��M9oG���~3C�m\G`;�r�^�rd1�̀��*lI�AZ�#�DJ�eH�Ɋ�.�&����(@��YR�Q�R�%��:
j'�x�Q�T�ȭ�6�d����U���~�DP�,8��#�ƻ�ʻ��$qgeR�N��~Y���ZoJQV�T�)�.M1pR�UQ��6���M>
���
�M��Ȧ,�rM+F�]�p,Ŭ1��E �SP�"1�cv�~'/)(Q(�<0���yu�i��<�=��Uy�{!+1�gT�y�+ll�yhDB��l��*j��i��O�j?�/�o$ S�l��ܓ� ���߆�9�H��m�=�U�֘�7A%Z�������{5ˆ��.O����AS C�҄���&.k96RR�xRc;F�^{Ớ�N� `"��h,}{�c*SI]x�Ć7���0�8S������QM�����`�8O����ey�*:�@�S a���T���"l����o�rK�l.e
RjI!����.�S��*��+�����mN1V�kGL'<$ڐv-b҄�;�v���P`���!!"�$�]S��LP��Z#O��I���UH��'�/�6%�h�y�!@TQ#R��ɪ��^%<S.eIY6�4vj��DP۴��^�0#C0�����Jd���������c�)�UX̫�F��[���3��|Aw����2AF��)���p|1D �<���D�!4��Z���Ρ���+H:iN!Y ��b
�f�e�L����Tç9Y�����7d���ʷw��h�)v��������!���VkY���T��4C�d�^�{U�O�2}�f3�*^��&�ŪNd�3DW�IZ
��FK����!8�h�/��^��UV�t��9��U����x�@���`%IEn��N U!�����[6^"�֑���^�[N8�e�hix]"��uek!�ĳ,nY��xS	ƶ�pAMy�z)7��,���JJYf��Z#�)1YA%[\���
�-�X	~���tx'ٳE����+�S�f�%`� '�:Z��I5F�K�.�4S"51M�Jp�@��!b�I��T��*)�k����ٶ0�8�vD'LA3�1��Ui�j�|���(� �R�^�t�B�*�c�Ó�Dt����V����w�Rȕ��S.l4��yq`��H��`��ˆķ5%�2a�
� U��A���+��p�_��QKu����%������X"�R%%�a� ��ŕ�!��3�"��u�5�ޕ�>��zW���V�d!R�G�ٗ������23q:
�LV ShSq�*�S�_���m/ױ!-�v8�ّ�)�"5ޒ��0�3 M5�Ԑ�2�jp�tL2�N�BH�yuZ�E@�M�v�{V��w�of>���T~����_��?�������]����v����ڽ:^=�n���|�?a�.����W��7ח�����<\�����1�����?ӏXzh�H�ǎ~�ҫ��;?���5�e�ˏU������w���j�v>^=�
�ϫӅ��o`l���c</n__�E�����������=v�O7���^��������t�� vq�r����?�����?�o{��__o�..}lz�uj���Ȗ������й�;U���v�6���ɳ._����z���V ~����W[I�e9�^E �M"Х�!Mtpp�I�B���d���u��P���B��`j�lH/]�l����8~/7��J<"0�D�ח��T�`;� ;R�ڑ%>�r.���@������J�0���Rb��˄�dma�Lк"#(7�
��"E�H@f�@�@\� ��ށD �xqj)�4@��Q��.i�p�)A`�T3��*��[v<�B�7��>�𑊏*��կJ�=��PFY�*��3�2k�k�rg�Om��%��� $&�Y�ȏ,�T��?��mG��8�xֱ�I�F��$�"�� �ҍ����a_�A$�a<#��u�����Ws��X_|�E��w��dU�H8S6�e������of�<�N�.�d)�]|��o�>$�O/8��h�D�Iv�db4����i�&�,��侂4�.��]���Y:x���%nlY����n�~Ӭ[Hʽ���5ED�;j�FY<�Hb=�[�������*���ܚ:�*���)��+Tkb�J�oDH�8,I�[��Z�7}5�'M\�K���7�^�Y�)��P��Ƚ�,EM�l��.g����ć+q�tz����#w�ЀR8���dc���XL�(��Z#go0�P-sA{�����V�$]�>U�j"{X��T�����? ��A
GӮ�y�r�٨|#wJ�F(+Cp�ZX*�w�ᘺK���A��7y�j�,<q%��Y%��ISX�fn���+�0�IH�� k[f!�8�A�R���j�J�m�غ��9(j#"n�b���
�Ke���k)+e�,>)@`����,��=�vAg�`"�v1�I.MZ�P@ͽ:q%@�@�*A���p��4!ʙ�]{=B�I��j;CAq��th�IYVe)�d)���y�WV4^93���OG�Z�1��e�|
�L<��O����-��ӗ� k���A�)���@��߾p w\!�gUj���?&�:gl
&�1$�_��K��T&��<m�}�����<�����7��G��kSXj�S�'�v=N��L6q�j7�C���p.G���������ZG�$H�<ʕ0�Z 7���&�,ю��=�Um:hm-~٤x}{�Ⱥ��	?����IZ��0]b4)����;M�Jp�$�Z�8b^�:I�1�̖RC����LI-f�R�0�j�$���䶗A�j�,ŵN�0�הWk��>NLY
ui����r�dۈ �f�!\��xJ��If6�%)&�v�'���f	tg��Tp1Ӯ�x;��1,I���0��F���F���I����y Gi�D/����#Ĭ���	��u��pF*��] U�l�M�a�M��)�1����bv]�z�X�M�Q�Ɇɧ �FA����x�ҙ�p�tǑ�/���x�X&�C<e�gK�T%���;Z>�j/P�Ӱl��	�,)W��Tu�u��Pws�Y�)����k/�<�-���H	裍`
�^�N��@*L3A���/����YL�%r� ^mW!Y��ũ��3SI��$����M2�e�k-gr%�,D+K�5���uik�����c�����^D�4�XU{�#�v�N��iM�F�7C8��-ӗe�u	G�C�R���gDx�m�dՊ1M%HS@RSK1�W�z��#�!E_����|HF�v�B��-����Uё�!��X�*�+�P�7g���D����+�i�#��Zn�'؈�jŪ���֖�1|�Rb��� ����8����RN
�T:R&є�e"L��U5��,��h�X�Q�ڔ�V�F_"^I�b�J�*�W��ЯuAju���PUר\U�aYA�,�U%e)�����T�8��'<5xU<Pm�YSm��<�R]��6kSb&@����5R�6'L������Zҩ�.b�%��ND���Z�ڥ�i����xq>�����tl�M��Bx�&��>�X6N%b��&$�a뙆"k
t���
����+��|h'��	*6^��[Ҵ5m�vD�����$kɷ�:�O��4����4�(7-�6U����C�^5q���Z'(�&z�N�;{���.fb6���������_x��fܞ~Hs�	��U�0��7~6ҟ���{���;ܻ~$����K����������������#ů�����ݗ��{q�?���p���a/�������v�Z�M�?�y�'0}X����/Z�K�^#7�{���~��?�i`�~�_�����������x�ޫuM_^_���?���:�������[�4�����~���>]8�G�G����> }uu�����w_>~�_���9�������������i�,�tZ�t]t�2�,�؍q�]MH�����F�H喲t\8�yE�D 8D��򁓒_��W�lQA`ɚM��7��^
��&8%�*�T�М	"+�BH�_�R��(I�W�#睆�y�@�G��bo�to#X��hZ8)A�K9Cjp{��s�K!����p2]�����C*�KmN��2�B�d1!^h̜�Sk�det��L��Nyq�8L�@����JRk��d����Ԃ�A��;�R���C��IQ�����W�D�"R�kB�Y��)3My�c�|�`���e'Hd��y4�q,��X��y��2�����8��,f�	����IQ�q�4�3��R�O_Zw�9���$	�*e%�L �&��&H�N��C�i��.8�2�� � �F���0ޮL-q^��#�{�����(�1_w�*:^>hb���W�(��GӀ�PԸ�I���CJ��x�(PN�D"����^�&k�&Ȕ��@�p`��)&�Zfo��)�l 駠�H�v!�[�ũE�����m*�Y֛��Z3�����})L-�a-���E�:��3��^��G�Z�<8j��?���+�F������>o����5f�j��%���)h�c�����oR��6'��)Ѣ^�lA�d�m�R9����t��CqLxc�B�T�3K�V��ex>M ٤�,y'�(U
�Id3Y �Bh���O���MKv��7&�F�1l!|8��-f���bx[��:U:
S��D��߄�� t�:�|�X9�%�i-JBx�6�Pk���TU�B$�3!$���I��C���/V(�O�21C�<���xq��S9\�e����]�Y�$վj�&D�z�ۣ�-L8�
��T��<�ߺ=}����<@��f����k����_�����zy,x��U��d��֫؃��A�*4 ����z@v;���tڪ@�笞�h<Uz��;5���ϓ����)_۴`h
y��k���p��c�T� /6R�v�5
 ��1����%_@��D�G��"0�����v*�]�moF�� ��Ҵ�tz��S ���\����kl����ۿ��!UM�J �&�͜�v)�P�tW�+V�$]8�fV.4�d&��Y��[�u�,��8��"�!�B��%��"`�TX_��i �۸,\��bU��û�|]�)�˲��)��*5%Rn*Ub)�R
4�eQ"n�KU<�l6�8����T�|ʵ���3)��{�|�v-�Hْ��Դp����l�����f8��8�����Sд�Nvzi���K��H�G�4q�\�@��0�㋥�!�*�22~}�A`�@H{�5����,E��    IDAT��0ՎG��fI_y��0����Q,`�3S�f���I��y�iڝߥ��>[	��5-�6H�;�ad^����5�v|�X7>f�
�-5B��]���x�� 0&�QBN`d)�	��z)i$��/+���v �b~���uo/RSU�W8"�|�k$5��9�Χl޴�஀0Rp�<��0�	d�C�Iq"�P���m<����FӺ�����c#��%e�e�b"����f�$�Rն;���:�*qz�DSD�ӆ49�x��J���ڒ�'��L�R;1��R�;21]�O�C)tDb[kxc���iS㋥2K`��,G���ِk��T�S(�8�.P4U�v���;���V�+�Wj}3˘Ñ��R���M�	�oI�D`)H�%%p- R�{56�5�$�&�L*����Y�g��r��8-�w{ԗG�j� u�)�W�vD+�CH�\*N���ϐJ"�W�r�d������FY�=�R��,7�fh��M�T�1A�!HZұv�J%2���GI/��MGJ	5Kc�6�����o���*10�|�b:�J��C�Ǳ�t� �4!�aʪm���t 3m������m�,fcX��aZ{ht��qwi#Q��ъ�V�)F`Dt�-0��yY���G�-�+��G𝼪�r��u�k\��=�I!K�ll�o߅S!�&Œ�1j#%��[ۿ��⧃cY�\Ø
����ͮ�lq݄�\�������
�ϛ_�_�޹Y�#և������O`�_#{����}�x�s^\ݼz�b�os��vW?Iy}s�.��p�z���H�CX?��s���+��<ڭ_C��xܟ\�+�Ӧ�� ����4��?�q���p���K�j��I�A��o��{{�{�a����K��^�����q}��q�?��������p�����м|8�|�������߼�ӛ�/�A{y�Cf�������+{���1xר��t'8p4���c��Eq�Q��پ@�}�f���@�.�d����^��7~��|��'���,�A�@kK�Q37C��)
|AYY�����H)4��K���<|J �ػ��b�Ε��M��Y��	X����`�(ph��0�r'��'�^nR�{�8�ο�I�l�ˤ�!Ka*'��xɚM�XU�K����or:�٦"б;H��0e�dq�BA�<R5B ��d�8��)�SӖp�a�Ȩ�IAL�����f��O0�1�k�S���d�7#�T�RX<�	Z��gV��cU���H��l�
��B�Й����:���р�9L�y���ܕ���D� qT���	��!��$R:&�\��E��FRpW������ǁ3A���A0�Y1���d���𥼟�򶳟�q㹣d�̝������`/`log{ź�ĵQ϶vkb=܈��%H�1/ָ�ѧӲ�'ܡ�O��.8��8PܒZ"M³s�o(����^���e	�	�pT��EU��}Ǆ�,��r�I�r��.vS�t�cz����axU���wa���`Z[�Q�kd$K��B�ł7�^F"��Z�@G�P�k/Q�����g��y��NW�~�^*��;��PS_L�����ΜO 5K)}�̺�30��)����"��'/5��f�T��3�BK)U�%���_`��t����38�Ętd��Ȃ�4y&UU$���ڝ�x�N�xKdV�|������ۦ�o"��\
(5��j	t\��4�h�P*��S�;�\�F�M�:j>��U[!��%^�%�XIU���v���O��+����R��H�8�BAS���6ַ��%>��Jp�*���gH����dh�`��w������"�C�r�k-V��$�ǎ_��Th�x�
z� ����GPc��@��ݞ��"��&��(�/%��W���Z�Me�-����#0�XwY�)FY����IYb:
XjDS��Q�_D��:��G}��gNҖ5v�NO��r�rCc8b����J\	��D&�Rl��"0K���Dd���aʊ��i�킏��b˘�>q���A�l�i�H�r\���RG]<���rUL;)-�<)`U �>��gL�	�&2�:
��?�TY�
���*HNv�5�0�l�-Ӭ��e�T�����������t��N 5;�'�6jw�)E$Z��i*L��).ey�L��9y�k43��֝��rH8��<�<� ���)�AR������v�`�� %f�mEk������I�,uI-B�Bo�Rtx�UuhU%l~t�,�m�b`d��רes�vq�i ���e���G0~)��.@1���b8�Y�ϗ^�`:��	��)��emA�KM-2p�������L'���l�M��*G�h��̲��Ѵ�z��#S�ד����I�`�	d@ Bj1yY�;�e�^��׽��^R����<ʓ�̯l�LwK��j��Hʎ~H���(Y�L��.)�N�<<M��4����>Q�ΈO��SP�$|_Ȉ�x�x
 ��NP;`C+�7��BֲI,��x�YS��ˁ�����$b!� &/N_ܜр��)	 �|8?����R�+��/�gdS�Qj8f㣵�e�&>L�h�i�}�"��3�C�𦝗���_�y�8C�e���;�����X��+## kM$�ti{�Y��*��D IGp��v���1f��&+��Z�J����B��Aq )W9,�¡_ t-(����+�&�\<�TL��T]0!��̒H�i$���S��IM0c&���+�y��eh��S"��V�D��.��2��@,q0�����
��i�Q��)�Q2��Z-X{��L h�8mpc��{Ȋ�8���e]0뫊���V
b�]m"�7x�BA�,ӄD�)��&�/��Y�x�w�d�tOmM�Yq��S�� �.*�5@R(}
ż�8C�Pn�����+2�����r�7������C�_s�-�3_��/��j��b�<>�@3 y�J¥p� ̲B)S)��:�R6)K� �;at�#;���Ow��/d�q���������i{x��\\�pqxq���� ڿ�O><v��.����]��.�W7ׇ�����/onw����t�|X�M�j� �׾j�'��5�r��̣������/}��vq}ܟ|�;�����+�D�_����W�~d�pzqy���
�����]����䝄���{�f��������?��4���{���?~���Ë�ݭ�����;���O����������9%����M���\'���8��?���;G,;� G�=û|F� �f�|୒?��wq��u��87�*j�Y
|C*Tb����6�4�Xjq��,���t�!c2`>�g��v��`M��׻�|������J�%�*K�Z�)4Fo:�X�5��!�	�MGlk3��&,P"�)>��A4Y��@��fn��6��4�GSeږ8�\���tpLS��q褉�5�[K	�sH�ZR�-����3)�4"m�ZM�Yސ����;o٩j�a� �_;8�,��@d�')"UY�,��\��?�Mu]��T`�&F87�eC6@�BWWgf�9��.k�Q����Eq�]'_	�#?�S-P q����os��<ӂ�@�����He�ߕ��y
x�rF3��eCR����?��1of�~��pK���ש���?��O�����ֶ׳z$G���hC��I{sP�db/ �|#ʢ5q����D�0&q�D��HY��yY�Ύ�TB�u� 8��8��&��B�k��ҙb�����:�>C�W�7s��8P���r�}l��W/�:�q%\�&��d�6��U�_
.^�1�|]t���6��:'���d-e	z��wB�"�a��d-�Xf����/Yw�o]S�u-mp���Tٮ`ǌ�i�����x1YÈ�6��K�j�P6;���f�@y�����>%5E�K�b8���/F�I�
� .�'�2���;=Rќ�s U��+�/P�Y���H��i
0IɊ�@�)�7[jb|My]�R�1��mF���&���p�b)��5���B��F��d��W
�?� d)Ȫ�K�%0jm|���Rj�,B�-K�\;�@\�u��N�5���W�W�,����I��ȷ�N�^�~=%|�[_� <@ÿ>�����j�<,��܄}պ��m�4�HA6���hTW����	�,5���){ĕ�B��M{4�G2���~�~�|�2�I���3:|O�>��j������O?%kBR�ɉ��f���l�L��76�21fޱD0v�B���T([9%��pK:!��t���U�͠����G%2|@�������o8˺�̾���!;v��ix�r�\h�pua�̀��:�j�ۂx+ZUɶ�3�kYG`��$U\ ��@Ё��|���:���[M1#���i	'�w9h�!YK�K}��3��=�p0�V�μژS!��!�IA�2PL���W�7�@/�.��+�E����^�z�֐R�9�y
55�*K�0
�u��|~�������R��@�w�h���6�*8f3w�#���ך���E�� �&YjRh�@^92�,C8�^
�* NcX�%��~D(�+�M����$���,�l$K��&�]�n� ����)0Y��RU �0�������Ʃ5[T�)�l��|��N�q�@^,��9�Un�]$��D��i��i�y4a���4ҥ8C�*������ >dc���h��%�ٔy4���Y|�H)��
,���#������;/ORm�Q��bI�@�6h9��
T!�h6��wԲ͙����
"�ia���3�9k*�|~����,�r h1!LkK����)L)�pYD��¡Y����B
�͙N̔�3p�*��GA!C��#x�&�	C2��J�';
8~�L�rM;�=���
��j���Kˎ�,�@��6��^b�J�	:�D̃&�y*�bYn��*	�<��b��!|�PUq٘�ǯ����X�F$}8�!�����۩
'BUb��
����)���DV�FY
Xq� ��7UA���|��R)��p���3)�vt�|�e�24��yKYd�r�$����u\e�qd���y4��{�)o �p,�ل������K}eq ��. "T��#"�eA�0��Sτ#+��Bad��"� |L�^��U�7Qd�V�vd�]�(M���G� �W"���u��j1#Cj'�.�kd_)*��/2���U�UHВC�t�Q�yd��5'\��TSQ�j���`��GU
���"�g��j��Z�մZ�Ǉ��'⋫{��~�����=�����W(/D��<>���W/�n�v�}��{��+����a�#�ӵ�����c�`�n�m��yl�7�j��u�	����`��������0���a�wD����:��K?%z������@�r^�!Nߋ\^��o�`/|z|�w�7�⻯��*?�鏹^��Û����>���nޜ.�~U�_>��.���j�JٝЙw��g���q�|g��=�����w�:jmy����刬�z_�8�n!:����ݙ��N�F�z��0�_h��R��x%����J��T����I�[Y�`���ul$A��~��A:s%����&�7����_��W��no������:UK�#ՋH-��MLY
�F�X"��1��D0N")c�� y�tbY;�t�z�/)/a���O�o�bv�MA#�H�
���:�e' ����騩¤������4����Z(G��C�~J����"�R�l��f@A�AZ"�o�!l2kwS�
-���i�U����bY�r�@>CcZ�4���Evj�q�����F`���m���j�tt�)���ôıL�3�<}`w�����ƃG+%&Np��s��qL�PnKVl�N�]7�r#�D�T�L��*=��X?��.�{u�T��'��Kw����?�����B�l���������]!�{N\�9lu���h
�aJ����d��e	vX��*�ё�g5��X65i6%h�4�$��4�\���e�<�%|��~�E�0gx��Y��g��\wL��|-T���l��8.
�1���x����r�Cj�8� �Q'����t�Ȯ�K�����[�;�:�h��ߺ�[ξ����!��8Ȗ���R�S�Zj�p�Y��;��D ;qU�R��F��X�F�r�������&�\����&�q�=m�Q�!<�6M��T�xL�| }�/�ڕ�)eB)�Z��=}3Qg�yn!)��uER曧�hȚJ5	BV��F��c���u��N����v���ӥB���HUR�&o &N�=z)ǯ�8�X;��ņ�j��*�V��}4ax]x�^q�=�0���^z>���д�;��}�בf��o-��`�"�B��/��·��sU/"u�}Mq�^R���D-��3v�Dn;�����^<:��b�~y��4�H�f}�b�uS�š�k�ה��܇���(1'��oX!=��B,�0HӚ��b�@����p�R�b_���B6v-FĲB)���yx4��I�$Nʖ��814�O]�F���21))%,YM�^�<��O?��C�����ʉ ��M��Ɍ1|ݙ.��T�}q4�q3���r-y6����b��֢��F5�/K.�V��<A�0>0Z���R�� W�ԟ��*�T�Z���<j����xPI8_�D���r�[�j-�Č�{F�X9���X�^�D(PR�.n�
���W����BI�ՊCh��Dӷ�<ZL� b�f�B`dM22�#�#���n�y�ЎZ��b���m�1q��@(�*�N
�Z�$��)��3�(+̦�-t5��Vb������ò!��c��h8)C:L�IM���y�<��� 4�.NO���`K>Z��y�d�5*P�Q�C�I8¤"������+Ђ� ��|^���G��� YCl]�>в[ź|�nE�;����ϊyq�Rؒ�:j8��7����PT0>��1M�h'�|�O��Ћ�^dI��%h�ni��y��,�΋��i�JY�)�!R5�3p`��$eM���rǥ
�iY�)x/+���1yF3�BV_]�	j*k9�b �-�ӄ�f �շ!!�ő
�3jG!a��)� �E�u�zEC �,�XU�pHj�z�E�!���[jy�
ԦG�i�e��w�����^m|�-s��,���
�e�fkw@���ږ�d`w�d��*�r��0� u��`Ȉ��R��pU����$�A���p���Rت��e� �3[KL6��TY��5� ^��b�
�M%%�w��u3��ˎ�Y�x��Y*7۔'� Z���oT�]�����j�h�Ĵ�@�Ԁ�Hu'���Rs>R��q��5<$0��3�<h�H�X��_3��҅���&Os�f��:m�"F:�';w�v7jj�}/
�0-�
bf3���R
�)?|sV��	 4��pH�¬�2��o�jq�!��B���:J��cB,k�t�J��7�jdIP�~��8��;�e֕e!ک-FK�2Aa��_�7îa�Qn��d�i�w�O�>K����'0}��{�Iھ`���wW���8���W7~g�_G�V�Np?������uԥ�~<�	�����^(��K?�y���Kb�>"u�x���>d�~�������n�����W����|\�H_�/�W����W/���o��C��Ӆ��<\�<~����?޿����7w��f��W�?�y�å�8��x������M������M	w��r�<�d.� ��ִ�m钉YW�鸷{@,�]W���;�?�7 ��9j)PN\���n�R�kʹ֎��yS�����ANY,+�%db����U��&K��,e)�0:bH����xJ
�7ܜ���]`����A)a�g���e����|���r/jG����Rb�����q��@ߒZ}1�b�27��5�v
tq�T[��B^	�v��f	/�Ë5m#d��F����"K�R	o�R�#}�B���_9�f��Yڗ��Zyc�;UK;m�o�ȵ��!�Z���vJ��
�+�[�r^����� ��em��-3�nE�g)�ɓ�@�yz����~��qW�14KgHd�8.P
8�R>���    IDAT]�8\#�j�X	�����U�V�Zǂ�u�5I��b�����b���Bj�W��``wE�R
N�9�R��6C�S1������N?����젼ֻ�6���������u2�9�Y��d3�i	�����(4_o@����B����AIG�"����"TΛan�j1�x����9��1�Z��R/�^l��owf�"���	�C�\mCz|8�W"ޤ�!���q
5�q�*̤�$�n>W�	��oHcw	�����e���a4R�)� Y���'U���M������&�NF	���D���Z^wA�`��cJx���@(�o޲q ,Zc��A��lS�%Ϣ���.�P(��y���y4��o��%�*�N�-O� �ڤd��Ԓ�^5.�r8C.�&){Iٲ,��ҁ+Q�$5B�eeg<��⍸�#b�8�fH��Y �x��Z2[�e��
i��!�R��Cl�]Cj�fKnT�BfY�g4S�v�)��vV��K���U"`	�DI`%&���z���\}��G�ש�}�'Ό��0��u���Yѩ�@w/���ş���O<t���k-ƴ�756?������o3�F�<1�,��&�B�#�-�z�y�8
R�>Еjf��x�{�A<�|�e�ץ��׵��`��utbFߎ���x�dy��h��!��&��4�C�C��2��W��'�Bd�@~J)թ��Z�1wn�Ù�/�R�,3d�N�.j�D�۔g�o�=��}���Z+��	�����$k��b){o`���Fp�NӁ#ӧP�ZHU8 �H����0y�@Lː:� !�BqK~��� �j�s�m3ױ��PIYUR��t���84H'S��91"�sJ�u�Py#�H�$@1���vi(��'Y�C�Ñ�) ��Bdf���@KddqHM{� �s��1ŉ�K���OJ
S��'ei�<�lZq�h֒7j�p���%�T�rR
��Q�� L�f��&�6`4KA�$��r`"J9�FJ�/��d�"!�f�d�K�j��oY_|L ��ۂT��)����8<P�I�Gc�"b�v��B����J2 )q�DKw�Q�7������c���%k ~^bDꂬ�Ma)B)H\
G<^9��",����/ň����o�pA]ʦ�V���V!��bVȌ��F9��CH�lC&(�dRd�R�h��6[�`�r���S̷�����[�b�l B_�(�@|
�h�%3��l�6N��X����kd1tc��PS2�P�K�(ȪB��1ʆ�{Y)"S�lj)�v�56�R*��,\��"��Z�ZR��^|��<���*W([!d�e�'n)˔[6��-�PB���xFs�!4�R�����^J��F9f-�l�Y��ZLwj���2��2�qTY2�똔�T�l�5^���j'a��m�9`|R�|݉����DN���]z��9
�� �3C�,ۣ±�ч��I�-��3�d�(d�L��\*�R!�RF�FRd�l�-K�!���!����3� ؜�D�� ��񲋴����Ѷ��K��l�g��P���	O�/5Y˹��c
b�h�![��R�
��ǩ�r��/������s�Qd}
��ƫ��yL�]�^M������,�x��ZL��F�݄M�Hd-ӄ�� >�_R����ub8Z��Zw���nO��4��vڱT��[6$ZA�����?oH�t����K���'��G/_�����#����kO���du������?y:��J7��������p�����x�;����(���[?}y}�^�`_X��hw��rj�mv�^n�σr|��8��{7~�����❗~g��W���=J]���}�'GoAW>~�_T������׷7W�����7�?����a��̓�3�O_<\8tV��x�6x����p���:��X�g������}�ar�Ӧ�������`�������41�@CN��4�.~�j�LA�l���`L�8�f��	祘^��<$B:��٪�ηF�r%R��)C(�N�9X���������6?V��6�,����&z���C ��N���Jĩ#Z[�IܲZ%��,hl:�\3G�p�H����r�b|��l���^�����~�M���dŲ�e[�MU�3I� �ġ��j��JY2����7^�L���]R��6�����9��j�4���!-Y���K��#0�z����'3�sδ>W�\*�8oy���Ϊ.ʻ:R��4aC�Y��)�}����� uW����!8ag�A)gݓd}�q�N�!��z	���v���F���IA�N����X��C�D+a��+�K�Ԙ����ϳ���Hy^�4�;��{�����p��/����G������r�����~rH��w�%�!
�	4�6V��x35�BL�L1��B�J���,S�`o��rَC<] ����a(TM���Gh~�$%@�XC&�( �텗�l����,~S����A�n6K{�b"F����˓Wd�B� t�4)�$�9���69��B�t|�!�T>�V�mM���S����?�A���1��E�n���l�.�B�Jhb2�]���#ÛY�*�cBj���\kq���B{З�'��Y��j�&2�4�x��K�	d�lط�P	_-�/� ))�v�cʃ�b�]��B�J�)���9A��h"�)�f��ʶ�f�d
��[�����Y��+�i�w��55��& 2)��0fH�������vM>L�d-g�b�.� h 8��f��lpL1f���<?-��!"�t�{�~����>s�3� L����ߋ�7^�^龌�b����$�Ǆ^}�Q�`g�U��Y������Q�>�H�I�!�UhɗScRb`g�,n#N@��f�����B����NY`)�i�k�Z���Ԉ	���p��W��ܲQ)�Ŏ�r[V���o�VHh0]��0 �Z[�hLm�ǁ#��I\�I��	
H�[ҡ w�`;IwE��g�t2<�F�T�'��:p%�K�7�����w�Ф��J�3a����Jo��P�q{��w8�ĩu)�� ����^8�C�Č� ,nx>��%;�ݢM��"��d5�2�N�y0�<�9:�d1K��g�#��SlBfR��&>|Io[Ю�;Svt����!�~��!m$����4y��~hģm�O_"ј��*�`U�l�U�o��{�Q���
)+a��w�k��rۛ�2ڴnG�*"�d�-�
��r^�!#˒'�G�vp{G�A��8:�cj�����Ֆj~Y
u�d���.j�m�##ls��1��W���Z�:V�{�Ar&k�JV��r�4+�k$�Y���e����}�rf�d
���ҕ@R��v,���1@�Z2)K��³��\��,.HD�RG�$eɖ���a��]URtl��X�~㮝2��{Y��H���`���v�$��F)`�3Ph����%5��s Z�6|%�J�V�3%MU���v�4L2�&ţ5[��B:LUZ��k�P-�rd~�äxx3�*�2�%Xk�2?)AH�*g�����s�ͬ$��0⤈�R�)N�����Ȃ��H�C�)k�H�B&�䛄o�.�v���,�©��Ex4��F��U���RyqgUȖ�Z,#{��TC�aZ�h��ob���R��(����A�<r~&�|4�P	?��Z;��9!8L��nZx~�,��Z:Rb�Q�фC�B��t �R�����Z��`,q4H^���Ժg|3��Uۜ��YUhbY�Jhj�B���M�l�\�v�33�x�p�����Ԉ� qU�24��~7 ��%�N1/E�����I>K��8�z����UYN� '2NYK)K&finm�^�v�pdK��^(�7���o�b���i{��3��Z ��'�W1|�"��9��]A�-��M���қP�����|�"f����R���+�;+���	�q�*,�pf�2X8o���x�>f�Z�������||��~��a{ѽ�	�[?�[3�_��[�.٣�W^�~��ʉksy�''�������v�櫇��o�=~sw���!}�[`O��~���~�:���p�/܌^�tv���g+m�N�.��˯����]�W7G���pyq��]�}���{�v�����w��o�f�y��^���4�z��;��D��\C�<7�O/�<��Ǉ��������yћ���ִ�]?;<�'�F]�s�v�-�c�������Bs����h�(���,W���t�8����@���pل�u�Y� 3K����[�N4���pYj����x-�֫�v	��~�h,��ZU�S
�Q�1��|����	��E�3	����T��5�(d!��P�^��!�d�ϋ�Kf0�k��7�T�J֋�$��$�\SݕX�SYq��A;�ǂ�1��h������	e��)e���;8�^] B[��*A��Ӑޔ��ґ�Ԝ)�@k
�-�
����0��Y�%<2dj��-�XUq}��$�h�N����L�ڕrD;���W��/r\k�R:g�94�8b&�����qojt����e;ұs���u��Qv� �,��T���1� %�c
z�Q	)YK�&T��#�|+�p�������A�S���8>�tt��%ߙ�\��O?u��?�f?H�E4��=M�_�+��{WW�4��ӟ�)́�!w�q:)����*`$_̈����֡Ǘ�&Չ�D���@�ת�����!V��T���u�F�ۻ��#`
D�D9M�r���8�hd!&o�DVb�p��@�T7��k�)�
)�Q�r($�˒����|�Y���3�*_�\e��:@��)����b�*x�O;)F�T>�������z��!�(	��)�r�R*߮1���u�)7��ɛ
�7psZֺ�8�����
S㛳e((U0}1��U�4dJZ���A<���8���'kZ-��[ŷ�g`�/A����zMU�ͨh��G��Ԛ�I��F��Ƈq:�n���2�% uϏN�����-?��t)�d�bj�dR��k�<B8��1���,i�2�8��ݟL�˘��_��jУٝ�)�Q/����ۿ�[��9eH[�0O`�S_���S�r��w+���#e6ұ���c��p��O�6-��+1��#��r�|��E�_�̗��e4ŉ��>�T_qFY��7
�b3H�qJ��엩���<ap�z�(1!��*LDP/�LUd�Tː�(8�6e�[2d ��yg"�5PV�
����+%vb1�`>�&�����ߴ��,k�&�y�c&�]$B��k���ׅw��e;�hH�m���;�	7`! -I�w\8�	��/�<�F�Yq̺tVp��T��cc(V�*��Qq������2��XG��@�Z�c����Шu�\��T:)�VX�̲u!K�����x!�Z�)���5ɤ 	v��J��� ��y1���N�V���O#)|��/5qY�MX�w��pG���l�#�B1CfUM��yR,�/���#�7�'Wv����S8.q],)��H�0U���U�YϤ e=X
z.m�2�e%�Y�S�o���VE$�i=H8L��2�`��aʻ�����Q.�*Dpbp�������p%,) f#�Lȳ��*��8|��	5��<~K������KK
��R� 8�RpR��J�gR�Y7?-��|;��S�<�B�i���T[k<���M��9X
��[֥*1ӫv���ͬ])����)�!L�Q�il)�W^
B��Y�SI��XR͖�hVN*�#T� N
ӨM+��������u�l!�p^yjp&�+�"(@��-��A0#(/U	~�,N�B�{:݇��R	Cc�j�XʼSE�/)���BL*�e10�b��g��K�R�R��Y��e��v��9�s����Ф�#�3��Z%�T��7	����t!+���2�>2Bg�г=�f��,��v�-�H4���M�T@�M^I��G�5�F���E�L�� �2���b�k�F>Ř��IuV�'� ���4 vW��Ӝ[��)T�����Q��p��8>MY1k�@#u�{�&��Q@-��"W˻|�񚢵<��ǟ.bdx`�|˺��Ҩ��V\�������%N8����ֲ�.��)�S��/��J�)geNU|�J�J�7�X4�J 
����]߆�7��ѻpf ڝ gͷ�)�f�	�p�����ԅ��i�Y
��+�6�����8i�^��Х��3�b�sA}}|�]�������L?�y�[�v}���.�^Y�,?"������o�A��7�������u~��t؟׏Rn7���t�?\_����T^PO���}l��ǒk|���a����|Ly}u�Y�[��[1�/��ߙ�[�~�e���? ����@�����W�ĸ���Ս����l�_�w�ޟ}8�.o��~���p���q�*Z�A�S넏O?��N���9j�]��ǲ+U(�!s�Mazm�ٺ߬\q��������t#y��?���^�n$
�b��\�w�3�h�-3?D9���X��5�*����h4ɦ��63��h��o�#k�=��f��M6w,RjUiA�I��P���`����Ɋ�@͠ߙ'�Fj�����M������3��۲rj���)#7eaI����.��U�� ekRZ`Bh��	)��{�F���)[	)-(0�?�w�l�'>��|T���l�B6�%��dِ'B'��5����Y�W�x7�T�8ţlɤ2�.�e^� �VL�]��gvt
q���u�]&%L D���N�̓��mB�ox�F��v}�W�3��7��mNI�x��pA���W�+ԗNGd��з/�>��
,% B���l���ej��O��������M�j\��uwaC���G��ڞ�W\衽@�T���Q��ԂG	�c*�;\C��$eI_vN��v���������Y9٥���I��	֫�k�EU4�
-�r�ښ�6����0�Վo��h^�~-֫'���ͬDWN��6�S��6�eѧ�ZWH� ��YSK�U�����,)[R�d�nJ{QU!5�.k)�ᛄ��5��xl	 <ӥ�
-�b��FV*���3�8���w`c� �ZD�i^�ٝ� a��p����y X�=�Wz?D\a}'o��Rd�J<��L��h�62��E�ǡoiBse1����@����U5�����a��Y8_�tꢰ��NGIA���r4KUti
T����l<Y#�-;�&���B������۸�B�%�V��	Og� ̫�W�#N�,���sI,`U���>��w�}G��
���������?���������6���y|���0�������vک�Jt�N���5qKALRsS��c
���{j��֨�!���с����@;�R|�|��[
<�茂�*4%�qL��x�ha~�pd�TS:b�4U�t�D�5K}y���yY4���-�� n;�,��
OVL�27X�%S�� Y:R�!0-
���;%N�e��^�H�7���v��<&�V�tnt�q[2�h�	���%ߴ@��Y�IMa��q�U�lE����I62D��\UdUӥ�R���ZU�+����ز��)�$%�G�k��62��.�����OS���u����$�J_�(�#����)L�\\;q�d�b*�Ϸ��]`xʼ�&I_�8��&�r4��e���!<�,%XVŧ?&)�*�^e�vb�szb��#�s8�.Df�j�F��j�h�l�@�L\Ӧ�!���4n�N-BV��#��g'} �_,�EP�-t��d��-�UAf$)�#.�!1-�rL���Q�y�C�*�|:*)���'�T\��U����r|��74A�3㝫)�<�P	8[���Xjģ�@���#��� �e�X��`:���15ʖ� sD
f�`�T�V��즴��pK�ic�i-���n�'�J�o�Z���8R�-)�޲i�3��I
,kh���Q�lj�Q�X��,�mM����i6|'9���&�W��R�*�q�
�n�eg�O�*�$    IDAT lڙ��6�TY��d��<L��)�,&S؄8ȲS"�V6������T�+q���A����ml $����@4F���&,�IG;eߴ`�A0�	研e{(DH�R�NW��Qf FG
Ry�D:�"��{��T�j8d�y)}-1�Ĳ*Y��f1����^
�I�T@|&hy���!����W��p��0	"�[U�(��?�S_h���T���
DS����.MK��"(�I�n�O/�:�L�N{�E) Ԏ��ZALd�@��,0�Z_�d�&�|p��*��9���6#�F*58�%��@�a���kW*�XG~J���@_��Hu�i��,�7��+�?��mJU
�w2��Ԙ�׿��bRS�V���7O"q����dZ�'B
3D_�n��Ñ=����߿��)��s�4����%"HܙTΫ�B�ܴ<���[�0�A��j�e��~����<�_�zܟ�~$�}��}�������7���{�P�������K����t�W��]�Z>�zx��|��/��_��ϗ~�����z������~���埽�s����7��7_�yHE�¯xR�3�X�k���#}�y}ح;�/�����?-|���Ⱥ�ˮ"���VU.����A.�F�.�xA�s�����H����16��Ƹ쪼�����.��A�#FĜk흕{93��<7v�~��ՍK�7���<_���=�ڿ��K������7� �ﻐ�G9��N=8����7�O��^>����������S\�����ԏ~��<��=��������ū���0],�-�&pu�qn_CI9�pe�����H	��o������w���H-�|�����|��+�J��o�gQ\�J�K����٢�w3 �U>K�:�͊K�)�K&^@�qS�wL񌊃������&�Ћ����kR�4xǅ�O�Ջw�p�*w	��6P�ajT���G"��	+o64�F����Uo��Z��*��C�{�RHSk`�Y�����|�������̩��;LLK�J�h��%%i��Yw�8�[�5�p�nKL処|�Gv�;[��6��,��XP�c�ڀ�,�P�/�͊� �B�Rw���JF�01�5|�<��'Z:<��:�n'�s�;����t�;�^�@���!�$�<��~�8p�Ha�<%p�D;H��֮x�
C���7���M�d]SY]t���ȞmA0qs�'8��0��AVe�)7L�yL��yC�/M懅������f,H������b�^M��2�X
�1�ed��Y#��΅g]4�%2ob%�d#��������[��%5�7R�4�l��b�N�BcT�_^�@��F��ӎ���AP�Xܸ��W��;O������+A��|��CV��˺d@:Z{�h#b%R��Ć����j�^'��=1��Qk
���i�ހ�eIDS!� t:RR�$ck��!���� ��Z�!�����d ���G������At��b3�%�D��-#���~'� P�y05'���43[���:�pZ%z)�ˤ0��G�M�1�M�MX�c�r��J��cl�i�T�˦#A�Ԍhb)�cY#^l�U��$����i}�Ȕć ���l��L�N���*��p���R������5�.�"��f �픤�˲!��/�.�>���=�m�U�#�0�0	�W�B�7��M_:=�p^
B�a��MM9�7Hv�C����Y�R����d�%�3Sբ]W��Dh�P˧iT����#1K/j˾zi��C�f���Ԗm�������!
6�<~�տ��+�i��%��}Rd��k���}�C\k4f�Owd�t��#t�p y٪x��^mӒ�E`"�F�)8M)�����ΐ0r�)Qޱԗ��Bdw �����}�Na������zP5�F���ם
����ڶ	�]K1��fn$qK>B~�����Ԇ 7vG�����1�S�m�A
l��̒�F��/�v��D#���![�0A��^m�1�᳐<Y����%S+���?%|)�p><�5߾�^S!h�j#�U��<D\#%R�N�$~W�͙T�vsD�H	��wJ��C�YF��i<�P9B֫���v�BIV��hT��b8�x-r�Z��Ad��9y~6Rm1��!k����y���&�Q�DPU\a���hR�*tt@3X���8}�e�m����F3��l�D�Pe9#�+k�{�Ď޴�\aA'��<�����v�N����������VmYk|��n���U��pđ�C�IU8)4`�C�3)d6�ӫ�iJ0#��`}���>�M����B7��`�iJz�:+�|
�VKy4;�y��@3���Y��5a�[����+D0�������n`ML/� ��B���v��˦
�d��l$�aj�R<N�� ����&l�h��21~d�x���?$�[��,#S`�֒Gc�j�C�[�:��OGࡈ�p��R@3*<dD,��E�A�m �D*G� �&@������ǲ�"4�7q�S5��b^���`1�j�0��lN�U����
"�H�x���Z[K��N#���@!Aͭ���T��>��+YR�R,��R�Ɋ���#�,�,�<J��`����şQn*���J���/�[�Ш1K"<&M+E�Y��>k��jU����th	�K5�l8>�@�3Ljm')L�����IɪbR8}��jY�>�#��9��P Ͳf���*�Z� �\
�xK)���}]��x4�@�����Jի � �{u7�O5*e)MS���.�Z���B�b�Z���L"՜pA�b��
v�E����g_�җ���wqu{�I������]�1N����㓧ǻ��O�#�;h%=ִ��Nw���㋗�w��O.�v���%?�y��Յ��tT~�Ǘ�Ϗ}v�N��K#mǸ�d�#�5<H�X���#��RW���������������O�c>1��:�{��x����٣+Ew7_z����=�o�N]�^<�=��ۦ	�uY��3��߅{we!^���er�,;vKGх���C��Ƨ��Q�BqY�����,}��xL4�.Y_j}�OЧ1>�5��*� 4����#�$R
�1�8���d�j6�ԈӁCR+�N�D���N�p_R��:��D������W_uJo�������.�c�#�f����u!e�S��#8��c�
� ���h>��T"�aba6U�@�rM�tMթΜR�a|R$�#���x�t�%���� �V�8���M"����ss_!S�-�ۯ0=4ፊ懸z�9��Z���e�Rw2����-D��E��-GV�����!<�)��v��PV� �#�P\;�Dp�J|咝�8(�%�����D�J�sdq�?P�|D*�2B�$0|��N�"P.ۄ�[��zD�q�b�-�*q�(OM���p%@Kû� ��,�,��C@hT�+W	�>��KM|���}��W���s=����O����F�PL�ː.D'�����E� DS+�r'UL?Y�!3�iNG�>/VnHFY��ITE�D{a6R�,P5�+��@J�������#,~�����M���WwY

�~:@�z��!t�	(;��#�� �79�޶��`������I���B�!4������v�����,ܲi�a�!oLXh�F��feu1 }
��@m���~#�F�̵�����_���N�W_u�l��?4Y���b3�ep-�-�����R�)�Z%,)�Ո,&�f"b��TM��"���%��B�Rb�R�WAH`
D0u��ђ�d�*I�y��X�#7I�je!�q�e{9ď�c�+�҉AX"p�ZW�TR@��S(�$f�
�Z��P;K����P��LCc��u�Z�YA%R��@��D��p7��{Ս���mB1л(P�;ߋ�[6M�QS���R��H���+0<�qe~Vk�����xY�	�w�y��%��H�	���Y��:Iގ�jLX���I1`�$I
h�
�́HAh�F�#k����5���@h�����T��0��+��b�p�Ԑi@J�L�A�0�@&`Rb�����e�Z^�8�*���$S��l�S(�Q�f	�q��2"F�E�hYJ����8�n?'�?qҎ ?@��u�U��SVe0��_�t�����/�VL�G wiҙa�h-y�d!�KU���Y��� O'%��ئ,��H��O��ħ�{/�Q�TU)@c�Vn)KM`���APUW��"���(U��y��C��Ҩ���:O���*	���RH�&�7�0O_I
!�,Y����'[�׷��X�̮��8��d�V>�p�H�U�(�-erq����e�f;�,f�Ȯ�����h|��X�#H0��Y9��T5�W/Ks�t��$Bٵ��3}û��J��p�&���S ��U����q��.���.Ē���++�� I5���#��[�.|:�L�CD9$\���֍�����;�ǹ���b�@��1��vMY�Q��2#U�qc4p�dc�k���]�	c���7�F�h�0'+`RM�m����d	�Ԩ���������!����/���\1�!��g�q �̐�X�XG7�0�ʐ��Mf#��CS�6��}IA�h嘳�C�$�-��O��PP�e��p^ܒ#��24UYH�v�l�pv�9%p��9,�]���F�Da4��	��cxU�%�ȆW�]ۉ�KH�K �O�֔�!L�Z ��-Ka�,�Z���K��@GA�
�f��gp����5f�3�Ԇcb
�#X"X6R��,N��1+OS� )��쾒����ܽ^�����_#%Z�}
����p��-�2"Jء�,o�
�i�@����X��Ys21q�g�o�yL����x��*��r�LU˶��m��l�6+5YUJ1GӴ@K^�S� S^��څ��+4�TY�er7��?��a��D����W�D�Y<��'d]ʊ{W��x�?]��t����}4��%,`h�++�o�r��� yY�uV��a�z_�7vj|�����B����F�6+�\�I�,ud���8���=��w���uo�6��t��� �7ΎQ�
����*ɮ.����T�z}�������g�n��ܫ{.oO���鹿Cys�Į'�������s� o/����Ώ_6�͕������~&���������iϮ/�{[�m�������&1�N�O�o�B�����~6��������u�!��t{�ÚWW�_�G=�o�7g�=�=�H��U ��:�k������}��x���n��������裏���K7��gW�ϏΎ�7W�>�߬�t2>x�m�cd��R.��e����N�.7�� ���&AxW�K�a]�p���6ߏ+���C�)�v.�ec��(��连�,�IY�F�w�� 1!B�@���Dn��k@�ć8��Ɇh�
��#P#@��%��ʜɷ��mW�'����{�s�{��J��
|���\kׅ8>���[/�*��Au�k���6$�Ft|����j���@cz�#�lY,P�3@����m���q�LޒB�l����uq�h���C��6� �r�|�������)�+f���?A)��Yj�?��ǉ0偘pGa�H#�,��D�y&%�9>)%�jq����A�)�G<}2��HdOX�EN̩Z�9]G�뺔�1�>c�$eSG����˶tuX}e�3�4q�
��˓�ݒC�*��YB��R���u3S�/����9�@Ɖi�,�۸*g��ý�-�g<{Q��r�n�'O�(���|�������n��쌮ҙ�@�%]l�:��t��<_���%���@J#d/9�Z'�fK�������$��r���A�-��7#�%B"�b����B)�f�l��0�}���Մ�h��ȅ��:��T�g4'�K˺��D�ʁj�p!�{h��l<L�Y���� ���S��w��@U�U��t�@
����k��i�!����	���^u��N��Ef��,�7�xëō�K�֞���'?Q���M%���o�+_Q��$���%����)�)�	LH32H�,�`���W^li�e+Wa�����[��K�vp>��bA�4�#�I60B �p�!�T#� )4���2Age����IR�7����r[�7'�<���r�)Gn~����#ņ#��"dI��ׅoZ`͂CHY���[h�Fr˅�t8�O�4b����F��^�)��X��ΤF\��$�^�z_(���&��;���^���E�����jG��0l�K�{�Mɢ��۷}�}GDI�Bhk��L�6^�pLf*��W%B�^������ ؾ1�)��s��!�f�,�����QH���ek��T�@&�-WS��r���+1��諘e�I!th5Yj�mʕ�K�$���qcD�e�^��J_ !�BZ֔7��R<��G��
�_`��vG'��IIavRI!o�5b@�� ��6t��X���h���@CQL�y�N��0�ئB���g)+fx�FZj�ỉR���ַ��4$2&H��X�A���r&���kg����!d��-��D�!^��U1H;꙳.t���i���
tJ�ٌQ9�����<�R28�,d1ľ��OV	NFx�Z�k�H}�q�� b䘫�~�D�ֲ����q�S(�v�&t���Zv�/)�deŽ�R��� �p)[�Ɏ%eI�2s�����<ZCZ�;�R1�1�j�@>$?�6�c������
,)S�Qd�4`�je�*�T�.p5��x�� f1�'B�N^@�
T�L՘7:ct��\���NM,P�����:� g�@���pk�@��<q���
[���$\���7�8���0�DL�-`�*�E����[�k�7@|
ђ���Z�$�i��Qᥚ���UŧDhY���h��`�Op����Sa�A2B3X�5-P;�BAy-�Y-
�3�Y�^i����
�y�,�Ɇ��e���!������!5�Tm�	���]0���hk6�6�:���B� QG,hLqS��o�b�-�]���͐B�k�<g�� ï$M��O�.)�Cؔ��B:ᚊP���r
8��Z�Q�X���9!�p�D�ө�T����A����OD!�a����d�!���'���L�* ���,��:�Q��^���y�Վ��I�%UI}c�A��_ U���l���t�-��+1�k�� ����GKV���zɊ�,S(�Y5��)յ�l��KYS�[2"|rCV%ei��vV��Q0���9���j{��CPմ�1��/�4�� a��QG1)�PĄ3�xLRb�#�[�yq�<MAf	�m���R���j�h��LGx}�ͪ�A��:�h<5�J�n	_Ǩ�?|yrs{}��߼}}�~��ߢ\?wy�ʞܜ�������}�s_��3���7�9���Ks�=�|��+����O?���D�i������ӋK���ͥ�"/�N���vc��]?��5�g@��N��ֳ��kr�O��E��s�b���������o�U��;g~���������~�����?���>�<����v�����_��'g<��.�:���+�1;����.��� }"�s�5�v�8ԁ0W����w���בn�p�"��.d��z��T�i]��i'����SLS%��[xC�6���cm�v��u�j�K5�8CVE���^*?�@�Wz�cA"4�"���/[�8��X��h�)H�T*���i�ϋ }����<Щ�p�:���&���/�Bv���֒�XV`H��H��y�ߟ����j�R����9&k/���q4�h@�N�g�u�*���Qh��y�3�X0��-8F��;��݄���@�I6��Ӯ*�i���3ₘ�;���	�C�u���6%k���G.F�C>L%ި�LӂQdpL%b ��R>Y��۸� ��=i�J�x��/HS؝	w��0IQ��.�^�b�	ǲ9��ޖ��M�%�p|�K�&��+nl�hJ4e�R��0�����`I񚪕kaZ��Vwjj�?�����/����S9K����@����k    IDAT�p=���k���w^}�U�j�L3�X����xr�T����~���Ӡd������� 5UY����t����I�M�Q�~��S�Ѧb�R:~j�;�_��h�yh�y_0܈���q�@�?�q���D�����H]��B�H�q���3L�h�7>5׮�!�}�E�R��P	�%����e5�& k��h�Ų$뿹P՝Mց�(i<̕�ŧ�t���A��cL����{?��!L9~��� ݣ~p�{�����_yѝ�	q}�"�# �hAh�l�1�*�l�p 2$�D��c�,`pK���C,yj�%����f���gH���t�TU`Z){�Ȓ�׺C��"�lYjē���QI�� `�Y��ƃ4B_���)��Y�I*�x����⪤�5-�	c�w��/�C杚�6תj �΄�lj��@��|�
���b^�za�c�r�}Q��
�[�W~�%L�ҁx�o�-� WA��HQ���ɋ�]x���曾����Q��B�F��b:��7��F�O����N�n����D�����/۵�[`c�����3:y3I�u$.��K��=�ř	m�&N'��O��*j�� �8RAR`)^_`ӚDv�9Y�vѩ#hI�MV��J_&���`e���DV
�c�j+�GK�0R��+W�*@�a�&US��z�lW�vT���i� �Z4���<T�&���Qg�0Y?��G�kQ��{1���
����#����`N�
��U�W��¥�dK
��YK�8)��Om�N։��I��	��u�bU�y��B�2Nh��R�+����\VIY���%�K��B%#՜��݉��������t/f�zu�B�$�����`��W�<�E|X���Z�vH�7���B�wG�t�}� ���e�2�b^
����6�ub|���:���4�J�k�� f�_6�� ?�00�e^@���.RC�!G�KIC&�6"e1�0q�hb6�`ۏ?��t�XU�y �x˯��|�����ć��Lat�c��!uOP�JI1N#A&N�BqKY���{=�a�F �a�*V�cY�.�I	���Z4^#�*S�#�"-yS�G��vA��8e��:dc`NI���v:ʚa�(�VU6uW��Zt� ���E��#�c���i`�ʑ�L6+楺C��,2+�U��#�
T�G`f1�Kn��k��� ���,3픋� �I�� -���/�L���(�=}�Ad����]�zU+fh�)��1>'^��9)�Ue�ΰ�x�H��WD<3����]�G@��ʆ�y)�l^���B�&[�*�5���S������-AA�m���FPJ�Nq/�R�'��g�H��!
t�᫢9"��BUSh)۲ M�SΛ3�@
�Xm�ډ;�t��)�e�
ᝧ�&�	��'"����^UP�XJ/)�ų���M��i$EA� T՚�i��C��6��
׮��UwxSE��IeԜ?��M����X 5��I.Bǐ�/���Jj�#�T�����q/v�#��NLH��,HS)d��+D�$��L�~�-�=��F���(d�3d�6���O'Ρ�W|8�*�@B�#%n�<d�Q~us����숞yv�r����T&�ų�'��{���?���O����ٛ�<�<��]_\��P�x�_؟}�vq���G>��Ó��>y�������׻S�Q֣J��ɺ�~!���zD�/i�8��s���S�v��	���A�/���[�ӳc?�s�a���ͱ������7���[9�NN�����{�g�<μ��������_������6��ݼ�������������~����:�����33�3tAe�U ��ġ����=�����A�.�zH��_�˴U�L�����G�>��k?��կ�֍��R����O|��C$ˆ�KlVǮ{�t,Cjʳ�&�-�Ov3�ŋ[6|:K1�hC>�G��n,�#�N
�^iL- ���SA�幦Ө
���Z�e��u8}�$�$HͲ1L����S���%��@�9���Hj@w����RL���K�Z��Aӝ�%�Z Y[���x8D���&�L�S�h��m�0Nғ��Z�O���������� k'�F�ݯ���h/�!|�?�[����W-?�U��l-��p��@��:5�ªF�v���� ^ୠw哷~ƚ�Ǚ �(Ջ�w��#u�.�K�B��Me��N�x���*� �	nE��<�I�������1-��(�E��B�Өa�5��K)نQ.k٨=�����c �� �Q$�l�>x�y�.b)/����K���?�)����N٧�y���X�CnV*N֬}
B(L�\�`2��.��.�R�X5����۪8�,r'N\�+�e3��R�2�dq1����%{���7�B��{��EEܭ���u�o��YG��S���jW�9}^���m�l�gtJI���<ߕ§c�e�e�:ܬ	��H��+Ү;R�M_|�v��Ѩ�*
��I�2�%�9؎B�k��\��G?���T��Шu�^�Ⱦ��
�h�׾�5�p�zu��=׈>�Pw8�<Rmʲ��-+�+�,\8"����N�V�-+	O�r��#���Ay)#	Z�D���\�C��I?�M)dJ,e��Qc��ż� ���X�&�B`�)�f|�(�*l6�xƨD��7���dnŤ��t?��_-��L�n�vk�_9����Z28ro�^kb��*_�h��y�40/�jե;�kؐ� �$B��~��_�X^<A� /o<&~3�[zk���~�����?�1g�3� �Y` �̗R|}i�,�n*>���k���e_,*��Ŝv��\YB�o�l��K�%Uy�4��;v��v� �K	P�䶗�e����@��XGYL^���X2K^U4�WŔW� �6�av�n��QC.�\A�/��k��P��]Є����(����ϲ�@d%���L;-p��c
��.k��Խ��sÈ����L�ٴ��e#H�%^��B��)����%�.��B�4���qU-܆Z� �nB��y�,����e�y���,v�U2��)�B�O���He-m���A�Z���}��g�	�nM<��8O�{���*��e���vLL��������2�eG�@V`β
-kg5B��16��-G�d� q�Ȳ^b�9��Ng���H���p�3
�L�6U#)�@W_�Yʪ��x�ȧ�l�Tm�	*�7���	�m�Q�T�H
�1��R1mȋ�Hi�<�Uy�eYd6�BJ��r��������U�M�G*<Y-��j��R݁�KcY�ej�v|d�D�7���v1���P͛L{��8�:�CRn��Z�B�t���J
���p\��JY24��yK�_KU^U�*�Ld�@1��!���r�0�u��CVb$`�R�L�3��
0�e��:X1á�W��)pR���}?���z	4j<L��L�H��1��l>B�	g���5MJ/"U4�HY�w|j!�8<��� �m;1+ᙒ^�o�;4V
�U.�U�c&�W���m�Y%����h@���h�QW���l��+!��
�y&�B"J���hi��qb�#������.�v����Y�z� 2� ��)A�f����4�b���� +�MI�;P�4��X	�z5Uq�H���lKC6'_	/Fc8������-��͓T#�	����_!D*�¡U�O��%~d ��MR�aIV����rԊ��~�N+��g!��j�xA��۬@y;U�\�)��N���?A�����B��ۦԽ��F��	���H��*���B��P�l�� 8����Xm��Fb)��!}��{�(Kp.Y
z�s�d XӔB��W��3��_��>�������� duߝ��̣��嵿����;^��/��ٛ���w7#�ۧϞ^���~w�og'��n^�=�l�ڛc�,���~wy{�^��W�[󃙷�~i�����Z��ezʸ;�;�������<���?���l���-���X�u�����������;�g�v�J�������ӏO�}|���]>���>x���?��9���E�+oWO����G.Frt>��5¥�Y�.�uV�7bN��F.;X�Z�n�[��B�QC��v����'ҕ����3?�ߔ���8�8�^|&���^��\A�pf�� .H��T9��T喂Z�#��ď<U-����K��e�.���(�8��A�O�� Rb�\S�H�l��۔,K���i�ut��5�� �}Ҩ����u�("���%����%\#����Ztg�U��v��(�6  1�6���bS!3�6�q�;��������,����WN�H�V��8M�R��"`SU�e�R�ǜ�i!N�aR�Ř�BN��a!8�ޕr�����^� 8[/p�s�l��O�=�P�C�>d���q�J�"w�,)�j�������0�LǇ���1���D���.[��vݽQ��� ��w�!��1���X�e��p1�L��|�n	$��|<��۝}�7
���k*���?�'snDF��z��Y��N��lC;��;/���Zć[6��ei&�������\��ҝ��b���t�^/<K��f����&4[3c��~�d� C`p�]w��4N�<7�/�K
�Z����^�Iy�Ғ 2B̮���r-Ty��o�R�"X_;�'�F�P����:jg�)E�l�M����Pe_=fK9"�l���Ą@�ݐ!���7��u��L�k�N"v ���l�bfdU�YM5����oqsRX��q��/����R@��-�:S�P.V8�p��ϐ���)G�P��DV>�S4U`j����vf*�uW��l�Zlw��T+��L�[�2�f��j�
����)��d���l�Rb`�U�m�.�4B�[v�n9�l�,�ɽ�ܨu�C�����A��80��]{�u�y�x�eL4��N��4e��0�����R�(�.�~��{-0-�����b���=�˳��P�
|�����5�����Z�%fx�FH�S�^�ͯV�H�ҁxGb�O�<��0����Q1;�@��l��d���,��4d��|L"@ۧ�_-�!t��Ȗ
��ݴUA,Ia�,)�*��r�aZ�1s|-f�Zx��SJG�^f��<�@V	��l�5sR8�-y�˻O���l�dU͜�#ؚ!���t�Mg�64���7� Z�/Pac��n)F.��ܿ�K�.�*<qY�/)#ёm/�hf�-����Ȃ�N�aj�[
�����ڡͲyZ����Rb�Zv� g�YkdA�
A��[2�5�Lxj�^�b�X�S�VwA�A���I��
j�6#5o�����^e!����w&���f��L�����*1��p �i)�ߨZ��7t�K)K��dK��e]d#Xve-�4�-�KV�	y �r�!��W�@�p1�k*`��@�)������
-+;�
ᕫj��Ԑ�Ȋ#��G�����K�$�l�Dj�!+��BY���4���F����^J#����EK�$^a%b�@^�*�����c6��Z������ߒ�L�`��M	&$��"�N<H�TY%M�x:��zReyD�Դ��z�C��4f���Z�jLU*�(O�Q1�QƑ��� @�?���!3��-'�@I	�SV�JI���0�����;.Y�Ht��ӱC������3�mS��T�n�w7�;��fp�m?)�
�j
�jY i�f�Й'�cB���	S���i��J,���A�i��,$eH_��OI:�]K� ���-U5<��nE�Q�]8"+�ë�����ő8fM�Ju�	��I����D4�;N%�ê�Ub�T���l̖8���j�C�ﴀD��*�ÍQy�8+U��߽��C�;<�r8�UM*st�-�)�.@���żs^Zhx)��H�ReU�^<�W�QnY/�e�R���W��T�u�&3;姝��r|��Y���P�l8�Έ��+�ӷ�Z�!��j����Ʀ0-�L(N���m޻O~eGVL�r�-�&��֋�,Sֺ�����E�?5q
|/ae)�YH�<<p�l)���.��V?Y��2Ҿ���Vu�~��c����n�1��ե���G��W���I^]_�)ʽ�I<�t����,}��֗��]_�/=h<�?>;���������C�q�����v�?�u�O'm����5p�۟\�e�
���O=ݼ��ң[�v������dN�FڳsO/�z��w���!S_6>;:�x���=<=��������O������oG���t{d��`}}����V�q,�:ؙ���C�(��Oo,����9g&�H9���r��"+V��� >��aD\�ٔ�δZ�0ǧ:�Z6ƨ��@�Kf�q�@�5���owlH�4`!����b�GL����!/ �awO!d	0gY6^IU|qL8�� �,��\>n�utp����,1}� t	 d�0O��r��KYA�F�V��41P�eUb�,+4� 5�r:U��,�-��XGS8k<ø�� uG�-D�ɺ7��h�b��2Y�1z�XV�0m����△����z	�f(Ng<\����UU�,�Ἢ
臧9���J1%[��dŖi�n6WǇ���ЇuȮ�҇�~>���?�����M�k�ϒw5��OJ���]��&��@�34~������t+�7X%R�O�T7�X��ą�]-�P���N�Y�V�αY�'���-�h�>�ٸ�j��]�����J����j41����v��B!^��Y�-^�ΈsdN��@��e){�z��� �\JlW���6,GD��u�M��C��Z3�z��K�Ҕ��p4��|F�T��%��G�v���/;U�[RV�J5��t�J9@)d4�{��R�㉴�А�B�.����rް��(ff�,)�Ď]�#��,{�F�ѱ3�eͩ��iS�P�U��2�,O����vQ�����l7������[�T"��ā����
2<}A�:��R�F�lZ�22O" �E�l�"S��}�68�!�n$)�8�ZK�g<Y����G�	lJ�0	�eK$�i�t
��%��6R�q���Ӈ���I5��gd�6���Ku�
0g���';�� �m�-��aIG�MI1o
4{})g��~�^M���l�Z��ZB���׭�rԮ����� ��e�����vc�e)����CL������x5��� ��4��%��6*�)l/:{Ԣ7����/�����h�G�S��;JV��믿nB��������S9�:ڔl��Z|>�$hu����XGͨjq"kW%% &�!3:|S	d�Z�F�d�J�������6A)1�l[NI��XSd8�*K_�)W�ٲ]$b#�b�Ӟ<y��Sg4s�oB��n����o �$�̀'�� �ڔ��d-�c�� ~`�����+�%|�{?���<��.V-$~��+���2]Ф��N2����b�~���"�5|�&�C�DP�Ҝ*GCH����L���i��%Y1��b^���P��D�7&��Ah�8@�`8��!�T��������S�r:� ��r��@)ִ�f��S��8��@6��3H�8K�a�[�bF����vi�p�����8.rxb$�8ն�97���^����x}y����<��U5vU�!|%R�:��lAd^�7�Z�d���f��໋"V�j$���Ԏ�T����f�⚦���K�͉5O��p:�Q�mGR5���4;.��DK��Ӯ@U����b��5'Ϻ=R���G�J4b�R8$��@۔�S�G6����<B�j�l)N���}��_\��Y@<c�ᣏ�Y	�Q����'�_��⑝�AL�#7r#Z�.k)0M)�mƻ�cée-e-;.q��\ �D�	L,5�d�p&h��ښ%���)Om�$%��y"�7r�FUĉ��l�4�Ec�!M2�ff��:~"��f)Kj���A�,���37�Q���    IDAT.�-��0>�z�.Y���(��M-ZM�Ք�,�8π<�N��	+��E(��h_h�"��p �pA`��Ԩ�f
���R,A��fU�&���o��ݽ^ZV+f
#h#�D��,Sn�-K%�i߽^�N�/Y˶�`�����NCx����~�ܿe%n�V�Ko�%9q�?��]#80Z��m�!hJ&%`8�R͓�eWX9�`�� ��?A%�ad���eV���mRК���D�~�<�9|q�b�t�X�;<�X��+Ȅ�Mo��1q̀�����C`�jq�J��J�K�o�����t�*��o$c�k)n��+�Ƀ� �$n_�ƟX��j�h*�０=��ΰ�p�����>W�ŏV�nn>{��l����S��<�4ަ��~�ǃ�k��S��k�vt������gWן\����T�+�g~d�ٮǙ�h�_�!����pr�ʹ�U�i�t���~y�3�X�_���%�g�����ã�G���O���h�O/���Շ��>���o�~�?�ǟ>�o�`�����kS��׮����ߒ�r�_�2O�T���!rX֕긜�B��0���).�s�w9��7�Ȍl"�y���}�����8� }&��w�{нG��ŏ���ݧI�Ϻ�yL&�@L�Tf[G�m��&�B�&i��9�����3��F
-N]�M81�C)K�fZ� 3�������K	/8RF��e��	������9�s���F8�FO3}>��7$$K'Z
p��ͪ�50P�3:�/��J-��b^lk@۱5���k'ǯ����g�zٸOS����(d-i�@�u�`��YNy�%��!ҙ�
�"$��l�:��.����B�������ٛ���>�������Z��~��~�qI��� .�@�T���E���w�-�0ϺX�LK%ʑ-۔�ep|�e)�S�0{�K�T���ɜ|o�͖'n4�����'�����BP�3��������'O<TsL~�7Y�k2C�`MLQ���mX���MYc�ͤD�_��U�ڤ�H��T�-�����x�����6�u��=�P%ū��i	�Y����`�Mc�I@���p�`j�bj�� fS�Q��"k��"1d'���# ���&�ط��-��j�Ec6Xw4�4_�QϷ,�PIY�h͌`Ɇ�Ɉx�����rf��;�,)�P�#k�˳	�`){��d��Pk<
n0��Z�x1���N��9�.N��fŲ�:��D|����+��� ��uTXvUn��Fٲ����b��|;"�*D��/���B�3������Iͻ����6"�f� ��JiQܱ����K)���$�M�Bٮ�Z�*��FA�p�R
�=
��&M���N�����
i
L���!��Z�zۻ�f����۝Ó�ٚ�����]�W��S���W�Cʿ��j(�U����!x�x��� )F�K�ۯAR�a��#�0Z������݋E��������o�A��z@��ȨZ4���M��R�f���6ҡyr�,=.ű��5�xC�q,�TË�MK�.h�(qz�A��tVIE��<p��y���@ch����R�:F8$C���p4d`�����≳�Mb�0��<2���_�Nq�J��c7�tGO;�h���Mu}yr�.��F�Kei2j|
���v�Djm�`hU�����0'Pmg�HK 1+�0R�1lPy8�+�.ŪR@:�R�p)Bt�޹Q�t	j��P�j��&h9U��2ͪf��Qd)ԔT<T��l%|�[j-�`�ֲiSK��9�Z�8�8��}��%�M�%��,�:X�4�8��X���)
�&���qg�.Y�IU޴
;����&�c2Vl��m_V�<Z�!�]�Q���{��ݥ�g4-k����L/8�pA��!�(�y
�!����jcB����P�]'i�b�Y�)�a4b-��[��D)G�#P (i*KY�L�`�Ъ��d�!�.'n$�V�4���<f"u�P,��.� ��j�)c6� ï�a_��p��"�lSA�mv���r�L��K��"ƑM��\�LMG �,�w�-�R� MN��Z���A<Y�BHy�I5YHY��I�#˦B��g��۹�(�H1%�
R�#�4�z?|�*��o�6�'�mG5R h�V,��M����ራ�G�RU:����R�&�'��%����)�~S�c�X^��đ�
�Rk�Ixd�FiV��^�T�B���l)�:���}1c#�)����0�*��i
g���1�z�Oa��%���^J�j˪U� �,N����+'5{�<Y^B��y�!|-��ۦx۱��I�T�Ua�FHn��x�3^����+��UD �5�.��*7����^� '�`hL��R�dզ|(gqxq�J�S���k*��;�k�6�rp��`R˫����^,��{�RX-��$?�(�Jp����'( 5��6�Z�3R�
���>D���M�%ʧrjv$KAJA�JDV��7�l`���h���%�v�?�x�UL��A_FM��]S}єH��<&\	\�5��o6���"YYH�v@���<�f�o�/��y+IY����}pI�V���g�(�'�~��߹��Ѽ�����.{��'8�쮞_y,y"�w�>�=�r�/d�\��n��ޏί^y��/�<}��h��N�߼�����,�����h�A�cf������:]�'GϮ/NnO.4�i���><�����o�����O���W?����~�����ߟ��O��l������h)�_:t;��h�=�=������\J{w:+�U�a���G���ȿ1��ǿ���~���o`���M�}"�9I��vqx��%�G7
I��cR�uc�> �t��5��eWS����d�@dA>d.=��t�� #�DG�I1K��L�*�#VT�3�|����'�����VkL�y<����������,YY���o��`�T�µY�U	�,P���G�#l<>��4�`�0��6����S� �yTn�jM����׾����l��ѱ�܄J�<���	ڋl�jݮnH?��%��g� ���Nմ���x��M� k�m�e��� p8@1<��R��?�NiR���F�1,��jT�W.��r����A��Qm�e�O>}��[o�!���%fO�<���t���*t�"�^�׾��e���G��ʾ�넾�8��g���Z7��T�;���]���Ww�lV���?Ĝ�y }��}Y1�%����Gz�P`b��vg��a��M�1�)y4w����׻�ۑ)�@%�R3�)S;hZ�lx��+�r�w@<)
���8�MJжۉl���#���?�B݁�V�a%����۹��A�𰜚��^��!���=�Uk;����Cp&��w���X-�O�q�����.�*^�&�\�'
@�uҺCF��+������;＃����)qY���Ԕ�Yj���!�<K&S������&�/e�6�K9���Y2)L�1�P�F�T����U�I�L�b��\G��1�f{��� �`q����D�� N�~�R�h8L���6 D�V�)g��%�4��a�@%���f��w�k�T/��BǞx 6��5���l��Am���7e#7[YLA�Q-) �P�i�P��b�|�vD���-p}�2��52�%3 ����b%!��6^jpU�Դ0�8)UJ�N������Rk��nw���▶�~�"�"���L���M��y���Z�D��y�gl��>�W���>��cS���/�r ����]@2��uHkK30���T��i�L.���+�T����t���2Ĵ�\S����̄z�Goe8�ͤ"�D��	�=CU%Eʐ�12�"X��o��
�-N��z�`��!GUR�����$D�& ^�@�S2*�9��(!�,ɶ#ji"0q�BF84��c�BбH)�ml��n�(d!��J_�0R�.z�-�C#�R�i��f���4����dז���R�l ��N"�0yUYA���v)+I��TA��
�p���L"��
,���<Ն秵T�!Rth��%�B1��cF6O��<y%d�-�֨R�ʒ��8^)�YfWA-&���U��C���
����S�SUʕ뫊5C�怦bp��TMP-5�F|(�Ӳ��LA�Y��� -@ҿ�?f�&6�v8��AL˶�.:�C+@��dm�e������"��l�cˤF��?���D�5\�O�%e�,p��#Z���e�Zor�Cc��F���H��3�e:j�(th�3-���X/y������`�Z�"�Ϩ���c9;t�@̖::����R��u�*V��E�ڐd�h�^���#p�)�� d�pg�֒�߹��Q�!��K�0��*1i4e��"��<_c#uOƑ��D�	D���;R41ߙ�{�pb�&4!2�I������S�&Ls�'q�b�C����R6�d�X�n�N�sNCܡũ�H����iw��k�;� �Ü^3ɚo;|HA1M��C,8��>�e�S ?TS�*���j�.�v�1q�aiZ�m d���W"hf���U^[ILِ6�T-���@a.%P@Da��L	P�P/%�A��@�4z�Vk�*�r���yM��r�
��H����׋ Z%����#�9|���t��eW���3ScbҀЀh�CcV�u����ߵ�.J5�b*4g"!4��C��;��:��r�-�˗/��Ͼ'"����O!Zj�GJ����W�0~;0��D�v 3��%qL�J��8N_M8,�rg��D �:`d���UM���Q��oʗ�&~���&=e�m�E}5��h��U��_��`�4>�i
���r�喵���Q�Uc9B&C ���]1�!`
eM��c�i��-~�I� ���@�!�OW���	��s��=�R}[�G���6*�o���c̗+˶�i�8�Oj�v�k�!���Ƨ���dj�*�A馽�x��f��>:�e��E���Bܻ�����<��������Ş?���I鼝����?|p���{7w�x�gIo>����>�y|�������{����P.];v^�˯�5�)O����Ao쟝�M�<�|*�̼|�GO}��g�����~�?�yxt��;�y��w�y��n������f�?̹|�sݫ��u.k��k�ƽ��wў���(Іt��8�|ي��(����R�1�k͜o����j�i���������DS:�8=�p�=u1uQz�ͥ���UO����:��T()"����@L�j�Ki	|NcՍ����q"��-�(o�JG<e��L��KIa����j'Z`���`��i�C��W���^M�sͮ�4�����"�
m�im��
 �H:�vCDY@#)���s̀�@�qY�z�Eh�x�R�N���@%p,�����p0E�3ƁP���U��'���:O���!��靋��.ZVj-��z(
���5��\�-"4�I�s��G|�ɝ6Ɖ&gr��aκ L�^Ȇ�=R��(ꡨt6M�sT��_�GOV�o�����^l�v����������q�����I��N�����I��KՈˇp����|������+���u����"Do��ِ�O�uk��1�3���ȵ|:4E�C�� ��8E:E�(ҁt����P�>ј����"1�t.��S����n����._�nՃ�\�f�}���oD3�VU��Y~�8��.�1�C��X�19����O	�:�F^���Y|4~����ҥ���R��%�HOЎs40}�BFP]Y�\)@�6:�RpT����U��>���0(�ӈ�&�&MH?8@���7F����ե�+�<Տ������2���
��,����c�}���Qҹ�'����^2�-mֵԾ��g��!H�~���K��Q��H�>��2��ش+"�r)�b�&��'(�%#��Kgu�ԉ�"8������>�+ad]`x���#�W�.�S
�{K�kۅ����(ݵ��"���Ȅ��]PNu�g��IC�@g��q�Pk��S������m��s�z�Zh���5
_3z���L:|7IS�A�L$�Y!�)���"ʾP�ݹs�7��1�H�hǦU�؞�"U�FW�%L��/���"����F�F�6���g
r�ru.ŨU�bj���D=�w@����*j4E����T!#AQ����b$��Ǌ��d[�Vo����r�B�C��(��IA�(��,���z3&��8��K��V!7�et�&�?YhF[�a���Ρ��N��rQ����,b�r��#�.U���(�ѶW���b��J��P+���w}�9��8V�W���BB%�,��o4�P �#1f
|6�c:I���B�F�V�mR[5��Qg������F|�q �Bբ�N�a*dD��*���R��Xj�����)T���'�)Z"p�3x���@��\��Z�� i:�����H#��a�Y\
�!�L�(&�Dn��#+͢�mZ��р�D��BU���89p~�Z�ϡF�S��F��L.� 0N��5f����eb�/}Ѻ>�hr�#�X9uX��Zx���b���f�P"΀�s ��W�#!�)[��OQ��r��gF��Һ�ƚ�-Ę���eB�R-�(QLH�� �de�Y�ixE�LE)�V��CvU��Ѧ9�-!'Y�k�3
S]�B����T�V
:�R]�b���S"K_"�N)� $)��!r��@铈6��N�תK�[]
��?m�9^W-$�)�L�T�I��oo���45���E�9�r�k���鶁鳥�B�j�3",��	Ԟ���b*�C�hH� �����U#3&e����1%�O-�`*��J�3~c��d���Z5��iɮNu�j!��d�^ō�l�#�$nd��J�A,ǔ9��L�R0�B�t �ٴ�L���\c�R����낦j��%!�X�p�##�a:B)mW㼎��W%~�H0!Ζ\t�X	�Pj���!-�T	�q��W���Ж��ڢ
�r�O-�h�-�M��+=x�f�l�EM0�����Z5�Hu�Bt�'�L��7�e������QN��vJ�r�M��RK�#��J�FB���K�p���-!��1��%*ͯy#0|���dU��F
O���S�@!����I�,"�0����R�N��3�>)�f����yF�,$_:�r�F`��:,���Ƨ	A�D���>�R�\�&�dB	v5���-��X�FRB	6�F��M�^h>��6S���Zwy��^z�q�ay�p��a\03���<�s�{��D�ʭÛxBҗ_� ��v��oi<Vb�R���υR8�Z�\�8"ࣛ�Y�瞻�㞛|�g^���������+O?�����{g_�;�����������8�=���~�U�~���l��:�QQ�88�z�lq����ֆ�L���~}����t��t�~����1�X���S1ߓ�ɯK����׵�|�=�'�08�x��#~���K�	�ZRK�F��%���+j4e��)���j��c��������'2�pb�0�e�r��D�/���}�Q��-�oӦ��U0��+�4�yM�75��S	!�C�QX%h�B��1G��\V"h:O�����	� �`TS�3��0=����Z؈s|�ʤ{H(T�zUE�yv��>�����<>2��W_�xkS!)j�!���Ը���ظ�~ݧ�up��t�2�5Go�W�t�AJ���� 5-�=�UuQxd;���������7O��_r������z��w����~yH�>�>�u���7���z�	�m�������)G���er�4�����8��/��t$��^�cF���g	D��m��v��8B9h�Bڐ�ll7��LC� rx�e��3�lS/��]9/�������/�� z��MU�P7� �M7���&u&+��R��Y�PK�� ������I��-d����(T�ٲ9�Q'���{yS0��u���+\���ۊĔK���1�L��ޓw8��h8�F�y�u*    IDAT��n�6���l#�Z�
�f����.��U��s���7]��,�g���K"dtp�M r�r�*�D����"#�-���1/����kO Z�r��7Es.m�h��.)�t2_E�P��(eΛ}��r\���:�=�WK��y���lMF��\��꫈K	�GОNDSn���?E[��pЀk�e@ShmaY8�H�	���VQ|V3�ӑ��JT9�\GK�͌�V%�8F`��rk^T�frD��Z^�^��8|-�&��[�Zt�-�ϐ�p��r�tA�oK��h�j��8�W��D�}_�.��,dUb: �N�`7M!�G_�D�2�L�V$��t'V�yd��*�C��2�[�:��:�N�˒��l�Y�-�����Si9��y�6���c�E��4��_`�����E���PEQ�Kз�o��fk�j�A$đ(�=T�o�ZK���Ffr�@�$���q��W�5ZWm-J�ڀ�L"��lM"Pkzcpd�q��x��/1�(�8J5�FTT��'8�/C�*���[�t��!L�0��+�~�74��"�LS��(�хc�%�%U9)6�v��F&��NJ�_��X��Hp�ᘖe5V^���6�h�a�焸@U1B�U������O�P�|!�Q�M[Ѷ�Ҵ�e�@��}F�	��*����O~�FV�R�K��In�,�F��8DY=Xf"��tRb%�%�!SV S��̆���d�mZ4�� �zv�&e�	�Y����:�k�Aѩ�A`��
qL9qf
��D.j�Q���԰����1L>&�|�J��2�e5e1�lt�����J:�||
z�� WE4r 8!�U\ʬ6�H��/����(o�!S����*&MN=�	��9q�[B"| ��Ҧ�ݔ8�^c-�P��i�@��'eB�8�:��B�\�ßS��h����G�0>��z3��t�1����'����|��r�O	�TIЈVo#aC�j��A��HMå��b�Y�64%�T�h"�09B��he���ߴ]����V�n�H�H��`T4�%`�/���(��w��a���� �j�$M�hl��@N㺬%�&G�L�SK!1I1�@���A6݊�{���M�,�SK�4�,��*m�H���io/]�#Ѹr�~�1
�L	���[H�e�Y�����%U4B��G��1��������
%>�Ae�8�R갔.(�fZ�t�H?M��A����i�Hn��8�)�)�(j�9RZ�ס�k
�O�|�^�6��v��F��r�5��<M�C��B[]"����b�1Ѵ���tV���'�J�*%���4Suc���4��IДՉ�FP�N���CHU�Iatړ��j��+�Z��`-їb�
aB�p��L�Z��R�)�f�_���D��GK��R~��W��ƘF�,�s���~�������"$>"9�(�Gj�E�ۦi7y�r�p��P?|F�����9� �l*"���Meu���vJ1M�D�7��3$����s��%�/yտ���w�;�:Y�TRe���i�AM���8=�s���d�w�AJ�+f�Ζ�{�[t��^|v���ڹ�0Iڑ��eQK�^ �P������N�.�w��<�8:��}}�o�z�G�>�����Ǟ���{�O?��O?��?��/o��W���ѽ'��<�_�1��*�������f��+�|�����pV+d�;pݚ��p��n�+�%�)�gPF̶�,c,d�`:�t8�A۷��������=�񘂦��s��;8tpL�$)�Lc�|�Ł 0~N�hu8l]�Ww?4���UA�q���HTH	���l+Tz����
qD��gZ�>M]��[�-�F��-��ٟ6Ы���ZפB4��\�,֫��5���\�(���P����_�j�k���"�1%�Z���dL�׿��S3�O��t`z�d�&n��3f!���-L!"���cpLE��(�0�/TF~&=p�9��R
��ÙP�D��k��-�M��-f�������e&�g�]r8�w5�]}},l��G|��7D�b��/���֒��(���)D��z��_9�X�����V�����F���	�7���O~�̭çl\hL���l"O������F�T�R_�ڟ��u�uR���v�8F`�C]GK����у��%�ѥ�!e�9��r�[!���vK<�n��"��ӱ[wdy�I�����MS�5���2k�}�&L۩�����l�����r�C����ʲ���R.���]l�u�±}JD+��)����bv�#��G�{�r!]��	\��b}�U	�vY��ņe��NT�$��[��!��d��8��m�Dq��aS��x��3BիK_�Q�u�G�B������zA�pY�q�y2}N����B��/ѕb8@�ӑ�ajޫW�D�Y- ��-���� �,L(�ݳ"S�p>A���}��j�i�)G��6j��n�MB�4��A��E[8��q�!��i�A�Z�sd��C�r)I�5)�~ |��4閉 ��t�\_"��R"#����bum�6*dJ���kKe��6��겤�� JT]9����Թ22 �q�QQ�z��<�>E-
8^n8jJJ�ֆ���՞D
z�(���B�aK��(��;w�rM���f$�)}�4}�ju4����PF65b�ReY�z��*�[�\#R�r�Q�5�`�Fk�ɗ(d�/W
')w!M|���ג�l�Z8D((GV
�>�S�nU�Y�4[�hF��8�R�R�2*�q��RKp�-�M�©[>��8@�#��N�)��p�4Y�B��=���Ek���S#�ÖV��܈򁕣��o�e?(��R�������5̌�}@�jR��e�g�"�3fE1�8%$�w�
�ܔC�� ���p:h��+��!�F�1�c�մ�Pn*�*Z(�č��pJteeU��_i�R�"DN�����(`���l�PK��Ő!�O���)����>r]q�e���Q��2!u+���^S�Z@!ԉ�_9���5�O!~Ս���<��V�nd�uR��j#g�DFX$�w�T]_~Sc{����:�/dl-Z�pf!�E0?�x~Y@K6VE:�tc`:RD�z�LW�h���Y��J_��%��B�L����S�t�I��J���U��`V�hB8��
	��*���**���p��W�M��d�%�ռ�95�O�t�b�j�ҥ�rm�@�A�b����%Ri�!�V�F&�ӎ<Q|"��j�&�V�J+��ޕf
𘕈�Q�8�lՀJLzi�܊��UpO�ݫՊ��tŁ�9��ֹ~ �1�Ϛ�lL�6Έ�B:
�B8@Ȩ�+�E���ґK������pg�R��H�_��5e��+�38^�h�p��b������3>�� |W�(r�����2��ǔ�2��:�h,q>sM�BF���I���1�b�S��
A����=�a��R��jq$�S��.4Hd �`H�Ls��oq)�F�F��
Q�MY�]�����'��JS�.��X��؊��LN�߽Z9M%LY����Gz�I�l*��W��A����F�#�t�IѪ������/%�f�w�S��E�j�t�@!�֩�h���5V.~�ٴ/g8@Y��i�Ȋ���e��@�p�m�u�t�&�ϊ�kh��z���ϡl?cv6�zC�k!�bV�� �e�(�A�t��0N
�i�L��d�hD�BX�8!DCD#x�˙g���3rݢ��t�~!��
B�O� ��$Ί��$�4�sZ�0+J�����P��VhC��b�[ _H�*���Y}�H�j�_�\���U�ʇ�1J�C�몬Rj�k��Kaה�����|��IGj�j�W��ޅ������`֢���#��o�5?�����������ݓ�>�������U�؁w}`sǻ�]>����<����:�������w㎽r�=�<<8�y��7o=���������˯={�w��o�������w�����G_���<���r����O�~��_tk�,i���M��;�*�U�%z}���Q��:�DI��w�N�+�q�7 =>��8F��$".݃J�hz����s�y�BKjQc������wr<^c��Ѥ,Q�v�Ki
��5�S��A-|���Z;�PLj���8Q>>�h�^��Y$�E���.�)��)���W_���֋ɑe�W�.�,�7Zo��V�n=xA�ҏ6�ߔ�'Uc^�6���إ���f]�F��ɯ���rBpS!:nt��*DNN{� :R�'����U�	�p�U�e	dk�T�uY��D�rz���Ul�>���t'\"��������8M1�?~�G�r��44�"|!�l�,�!��>�ش�o����|Y��X��
B6�ۓ6�aq����_��>{�||���^��w���?����{�G�{D�\f���[��/�칺����woܺ��_�z}����g_�!>�����/��RoQy@��?�Iu7"*j�������U��54����w���j�'[(��]9Tj!觢��e���P�5� Q��LY��2z�
@u�
Ӈ��
Ԑ-S�R���?xk�F��?�D�*m
��˥ 1*g,�ϙ%�Af�$�P�VD��IV9kL�Y��n�LiV��=��rq�7�)�eo~��9hNǅ�H��9zCh�|���V�j�%#+ԅtu�l-~�S�t�4�Y�+����bw�N|y3��h����\��HIܨ�D0ьnR�q�ږb�:6�H�^Q����1���`@L�b`��j>}!�pT�ƛ����L��D�)� �Mq���k�sM�6$JQ���ͱ]ֈI����1��Ug.���妳~O��A��PӘ���*!�z���&���tFG��3��,�qR��ui�_�Y�����ĈXYS��C��mB��_ngO�)ҕWSK?��k:�{V�n�ʵ��Y�e[T���:>A��C({�X5Y�C��u�+�۷o��+o����5t����"ކ�.w'�)J͏=-�A|�zVNG�U\4G�ۙʡiFi�R3J7}��EK4ڟ� ʱ���Ct(].�hb
	Ѭ�DNQ!S���OfuD ���|�^��#D��>��O����)�X{ħ�8�R�r�UA�RbS8Z"Z�ZWΑ%?���MM�)S��iN���@�S�]V���|驅d�8@>���N����h#�(%p��zh�r�����
>yD�# Í�A��U��r�@�+H��98�K����DM�*z!(ᴋnki �h�J�RN"�'�zӚv��l�����%#��g#��Ίr!ӃТ���!DV]ش��]8��[ �0d�1>���>f������0��`B!j�ȟ~J0B)J[���J�noW'�PcK�P;>m�/���f��>�W�X!�R�H�>�U4<D(S�%�P34x}9���r�V͡Y"B���]S:��9hCJ��#S�&�1��T���&�bf5�ϡV3ڨC�Ъ¡Ä����6�@� �n�!r�Ǆ �`�)��C�
��h�����T%"��ԛ��WqM].V��F
�6a&�K5S-! _.���1֘t�gф�O�D���/׈�NE�||82�!~�Z��8*�]����q�-Zk�I�FӢ��BE÷�L1��c��)�����/w
�<x)����q�憎R�t"FHR����6�8ri�m9L�A���,>�Id�Msp�h8��J�q��Lz
p�Z���e+�(ڤ�I� |x'�xLc�ǩ"�������)�f
vR-6)!u�Lz��W
�Ҝ(�o��7ѐ@ʜlJlE0��2�Zm�U P?�@�NW�~פ�7�đ�Z��.�Bj1M�Nl����	��Xzʣ3�p�5Sf�Z~�J��_^!�E�������¶���rN�A���d�^�
ɪ���`,�(+p�%%e9��tN�����>x���ܴ�L�h�h�F�r-X�8E9����SN�(7\���!�t�
A��h�r-ǈRE#��R&���8�T8�A�#D6.B������~uHDˊL$eSd�m�q*3\
NN� �C�7�>M����-H�8�#�9+�&�ʺZl� �'<;P	��V[�B�>�V�T���l�	���Xh���$�*��@�8r��h�o�Y��W�B�Mcv� b�Ә >D�.
�)?�k�_?1S�$GN��I����Z2��g�|�Ɨ�Y~��Oe�_����3+⃕����K�%��/����̋=�v~�Kٟ�����8ޒ�<�����/n��=�y��{pF�`�������Ɓ?��7��.Yӻ�����o��M�ӇT�w�G��w=�9<|�������w<�z��\�����������=/����s;z��Z�<<^~���72�ﾖ��`+Fp	����?|!6�8��#d{m���#��p확G��Ms{tH��f�zy�ғ(R�I��d��(�r��q��
�������j����)��pѪ�ۓR���#1eNU��G_��)�_��RPWԴ��YR[� ��[����xЃʟ��g�&�?.�.��m&���W\�FS�")�h9�~I�%:F�A)��8Y� �Ę��".��Z+���͓�|Q�D���!Fsh�ЌL�*�:��`C����x��+e��E��.
a ���F�Q��Ar�L9#�:�j�a8!�\���Twh_I_oZ���C��2H�6w�66})�L�H�&�´���ى������?r����t����䁿������=�����?������&"�q!�����r<���/M~��]~��g�?����x���;O˟|r��f���Us3Y.���xS�7"ωU����1�D��3S��%qL��5#�eq� p�X�z,�8xnz�����������aT��*���M�1E���{��[�%EӖM����7�brHI�f	U���E��]K�F�	sH��D6|~��Ɩ �=�3�Z�RӃwVu������o�|υ�롊{�-�o�{/��\��WK��&E� M+��ԛm4j�e���7��x��24_ހ�v�!v&�W��3�S]L�\�V�c=IG��p���`q�P�Fk5ҁҞ�"kZi�� ME[�&;���D b5��m��#�%WcM���ԲR��z�#��;ؘ�Z�,*�w6N��x[�}��~����#X}�6s�b��mճ�Ɣض׮
ѧ`�Jb5��rt�L�F�.�Q�e�	�#w�(�@%pl5�h�>P];�^f7�`J'EY��n�t�>�՞"xY�J`RӤQ"��,�� K�c{U�."j�c]�K��2D�r�Ʃ���e�thQ����?ꄓ�#�%�N��$*d[��OM�i�luz��	qX��#|G �'�UY�Կ)G��6�6�W�E9��#K�/j�D�%��[ێ��YfQ���1��n8������88_����j@��_�����_�EM��sQ��]Djh	M��
�C����r�\z���G�g�(Y(Ј�ֹZ�N�]�Q�	���8��CS&�T:MӔ����iQ)�Pc�ߑ��r�z�J1V�O���}�k���D�#H#2�r_�F�jš����,=���d���$X|
��
�t�-d�('�(S�8Y��F3�GPw��]�L�X
&�6���pc� 
ń�"�-R3�V�{B%��A0MوPݶ����2mT�ؔZ��@A�߱�O!�q��|
��A� N���p ��@1����4>��[?d�j:���,E4���j�n�e!���!�&��O!S~��0e�y��r�V��k�*�-M9Y5&ʧ���ֈIY9>fj)�+Tu���L��THb f��eR�Z᭑&_VdcL��S{����V�r�9�p�N �3��K���R:q�M9i"pL˚��	�䇧S��l�
����c/�=�Q+e48�\8)6�z�����MQ�ȕ��H�&d*�S�hr��I|c��RJYJm,�:S�)�?��P�o5�8��0�҆<�	�FÇ�Y)���4f�c�&����T���Z�X���M����p�DT�4�UO���M�v@Q Zǵ���&QUI�*���2�    IDAT�b@~�B�+�geEk�g�FH�� |
��4�K��S�b�I�9��B|7����*_��>��J'�V=�d%��Wݸ��W���YJ
���j#f:)��$�x~��HY���d[�&Eь�L�ғ2��J�ZR����RFMtˬJ��S�[��˂c6��Z�*1���<������O�$���d*�A���r�۞�<��ۙ�J	�Y�Q����d� ��p���]�YQ�!�ˉC�3�i����p!Q�(P�T]cd`����C�0��0�[&���d���"ck�_�J���I�(MLjF�@�����at8p �M��I�G�/�7O*�������ޚ��C�m"���E{ ���S��Bj��骙2Q)�Z�,���t�6e��'��g��81�$��dL-J�m���qj��J���č�''��0!�8ub�Qh�|Zw�a�6��z��/�.�׸�)��_B{��=�=�S�_���o�t��|��ǥ�q|oy�R�]vN|��q���`�}���>�t�l.ojjϻ0G7n^�/�s9;�;�7�vn��=yc��Ǽ�y|���_�߽�����Û��w���}�Ň����қH'�I�8�nO�O�I;���q�|�b��"�ɲ�mQ�ٞ��6��4E�
�K��1خ:	=P�8�����$?wC�v�?�O
������(�QV�M�Q���ڶ
��ɑ�!��Q�y��������Țr�Q�S(�i ZdN"�^����2"0�D��?aM9��e-��7��22��h����ҷUB|���3d�v���	�\��*�y��������p�H� �L)���#�S!��L�Ǒ����	�
տ�B:�D�u˧��rK��hd�D��S'���r���Nk�����O���\�I��G�P���E�����%yc�pd�_||�&�Qm�VW�#�В0ճ�|��6����D�`c#���t�z�?x��g�g���~p��sqxc߻�.��x~�����W��#G�<��/ ^/��ͧCE٫�@�F�����|��Ǟx�ۣ�|���?�d�p��������G�X��Ф��g�ӟ��7����Jwt�Pt��(���Z;9��1��5u����mkǀ8%�+� �2jw��M����~��u�h'�K�jy���-]�e0O��ё��c>G#���*f�@��u��F"Q
����a���$c)`fJG��S���K�q
���QC3R���V�>�1&"��p\��"������F��{m���:>>e���vJ��U�U��Q�r������^4j��K��*���z���Ш+/;ϑ��TcpU�
zP�Z�������_'�vl�tYNk4m3Mk��Q9��--���ҡQ.���tp��]A���= f�`]�U�7ꍣ��]G�~h*�k��-�|���O!м��c?i2��h�]�m$E�8�׿�Ԓ�xM�[Qo^��z�g/Ʈ�wq(�S�B�E!�M�v�q��Ar��t)��7G$���վ��$�%�5�l!#�Y�~��!�1��X)�vC�����䭷ޢ�sf��+]JՁ��H)Dӊ�$�"�כ�T��.�u<�Ԁf�+c.E�ҁ|:j�du�2%e�G�QV�4�8R���Cӭ���( �������5��&�IVH
Adc�d{٦i��Hi��H��D���7�(E9�fĬtS)m�i�q�� $���ı���0�tQ!���jK��'0'������.���B9�V��i;�*L]e���,)���H�a]ɚ��4��Y�̙��ZV
H/%�-'M~M�1Eփ]r�'��� ѭ\����8I��V����n�7ِ�he���Mq��x_�2�
���!�����WH
��рR�"�ƥ��v����C\
�G��j!��� t���h��Yò8ј�)���#G4ʪJ)u-T9R95P(����PKS� ����z��o+j����U���e*e�,W�B��M�*��N"� D�׌����9F��e�b�O���aS�oC�ed��V:_瓵��6MWE[o������� ��NTJ�T�1�16�O@�m��!_��p�PS��M��!5�$ۺ�6�b��I����u�8ت�p7�cK���B����C�B9�� �0YB/L�&�Z������Q�,��|�,N��j,�5Y!�I����t;�H�-3�Q����C8��H!���!,&��H�+��J��雦)��O]�,�Z�sR���x#H���L��J�L� �\����!kz���eu��Hu���rܞ���U�4��CL�@��M�D���-���+ĩ�#���k$����l��H�6�>�'8�vEH�;���4�I�r�h��>��R��<�h��hjͫI�-_��8hC��Muc�D0�� f��3�cJ5�$�`�!Rn����jZ"��G5���BY遦8XLQ}���/��D�,��S:�7��?[�~;C�S�SN
�)?A%��ݲ'+�c,Z��^-�RR���+Q
�^���rj�Sc1M����B��%�r@#5#0:�����đ�IMz)
����ĔR�B�Rp�Zr%L��O�tz��N�u8�8B^b6g�@��n[jZ
?�,N�ޘB����)�D!��]-
�T:2C�	ԛb,�3�Pxˤf�_T�[�
���\&0�o{�i�isJT�C��(8�r��V�|�:���s!L# ��U�zL ��Y?�^8XK�h�3�����Q��i!Y�+"K�ƀ�������EP�B����+=cFD��D�pj��Ili��eQ�����k�W�E�h��5�{�G��7�gM� &���=�	$�?�����H���'�u���9�_R|��p����*y�5��v9�����a��M_:��ؿ8Z~��������季��n-o�<�8��p���w�|t�˻��>�9{����;�g�g~�����T�V�_]�y�������S��OB��o�ej3�%>k78J�XN;i��6��-_���}c�J~5i�,�x�i�7с8��3��M��Ka�JKD�P��<�3�_n�S^�U��9�&�V���.��)�|"��Ʀ�F��!���H'��
��0$��Z���=N�9��7�L������d=��.�K��yH���������+>�Ap�|"�R궄�k�#(H$B� tq!7�6D"~W\9�p��VǑ�$>r#�a��d|+m�t�r�����6�&��ȅp�նqվ�����SPy�"'�_��hd�,8|+�?Y��O
��Hs�}Y����������ѧ�1';���[x���|�M���n��~�;O�|�ý'��y��O�ν������?�Pp=S`.O�\,�����G�����g���?����t�{�;{/����v�ܖ;O]=W�'M�P�RHW.���I�� ��MJiS>C��T�
L-D�:�I�O*ݛh�4E���[M�����+���!xm��U�\��jWmH/�i%�49�^x�-Cs�DH[�z�:���Ѵv���^p�.�ur�42��q 4�9@RVn�%8��N��4)��B
�Y�����H���/l��C�W8�ݾ}���-M���QȦ�*����������|G���HQ�q�4��1cYoIB�:�8��l��ŕ�.eG�?�!��Y��P[ݺ�@�r_��Hd~��\Aʲ���32ߨ��~�·��t�h�rcr�1-�Q��,Q�v��5)�njT��:F��[85Y���l�n�u�$M��e��&�Z��1	��hކ��r�Z�F�Q 
)��&��Z�ZB�,��G��@��&������(��4��,�i�0וui�*�]8u�Go�4�����R�^6hJ�9�S0�Hi�U!ދ��їkW���1)�!4�L9��D �f?���(_T���c�%��J�K��W�\����
��:�zQ�:� �4��v:���f��lԒDQ|`k�ӏS!�
U�>~8�T�I_�īh4���0E���`���K48Z=�R�|��h:���Y{��R%&ā�©%����*��!�h��Mcr�W��{�C:�,U����д�l�(ZS���\"#ȟ�Bj������N�ҽBL�X����A�'Ғ��41�=�QdYL]K�ĬB8��[��|Y�qL���8�sX`� 8@ǿ!C8
q�Ahp>��c��:Njt�Rb�1R�ʡ�l4�6)#ǏV���dr_����&��5� ���B�*GE���J��FK��kQuc�#�2�@-�f�RB�PK�+]�Rr�S3rqڍɒ��4�!�.W'��fچ����h�E�� ���F�ea�I�+!:` ��TtN��� �v�0��h|�DէV�MS0f�ZV8�R�|���A�r�jihmI"��#X�F�ҧ%4Ӑ�N|��w�8DD�hʡ����1�wӘ�A�i�C�瓒5�k��p�P�����1����d	�����FK�r��hڎ�¡���f%�l$����oRu!)��1g��]��1ۥh��N�<� �Ԍ!F��@ui�D��6���E.d��P{SBc%�	��
"}���Y/NK�L
0�&�(�iE;�JYm��j�%v`�j�ZZ�� 4n+�"@��!i�\L��-
�Q��۱�m�VKh-j��"�C@k�$�O�ZM�	��ɦL>r�E��j
I4���1��et��i4�S��\��k���i�	����:���ւ6	��)1)y�b�NM-��ڨ��qZ|�H��)�)1�R�($¶��r���I�B�� qX ��&�4N4���#-�X'Ʋ�HV(_Vˬz��)��%ވ#=�iӔL�2q&�f7ضQbU҉�_QR�M�4NVN4���qD}����p�B5�g%�8[�B4��.0��0�('�Ʀt�4�d��Ȗ[u̢F)@Qf�����^;xdQ}"sRK��5�r *�Cg��|��>�@�8Ց9B6S��K.1��B��i��KG�� ���8$��fY��ك>�R��H�F0��TMR��)�6D��!�1M??�����c��L�?��8يV���To8�6A��h��%��/���ǥ���%zxD��zg��G���}�z��REo@��������΍��ǎ�8{p��?��C��<�5��s���lO|��a�=�����ࡍ�=������˽}Rӧ�.o����������"����߽��O.?�뗢�?�I�[O����}�'��=o[�=8�ҭY%Ш�tqz�=ӝ��.����$X�[�M�c��ĴQԶtYvf������RO�<����3C���0�4*����)wE�s�a.�P�����hy�ybgw<i� ky��T�'RH��VWK�k�]�)��&�4�>!��%gC+ME�M�sr��R�ǜ��-�&˩�h����J9�n�h�B�z����21�~=׍�+!�k������D��br�8Ԉ��Hv� ��">A�7�5ʲ'vFæ�^|+U��(��#0�w �'e9]���@����,w;�9д%�����ܾ}ӍWȿ�����h��3eN�x7�"�-�1p��8!�0�h��]B���=�f�gK �X-S�*&oK�L9c� �m5pQ8�`�3W�������[~���{�'�~��8�<{|�[��>�y������w ���������ޤ�˽�;���}�>}�v������@|�ӏ����_���o���;�\���S�<��������z�o<�ܠ�������)��ܦ\�;w�W�M���� -���s�� Xc)�ڥ�4M�
hN,?A��e!3�i���#�%�N�=t��B3d������_��W:t��)��Ty�L婰fJBuIH%LZF� K+F�t4�,o�/%
Y��-�
IO�`
z�n=��I�(XcVQ�1)j�G)F=�H�!��VK(�gB�D�P� �]�'@�� R�k YiH
n%�tB
��a�9�fZ �So�֛����4�WN���ѼO)�^�����g����\��s��u7դcPc�ۇ6��Z��������%jI?R�6)d@Ǯ��.q��)��J =�כ*!�hVm�����Z4iDctj��B��k��n�r����k�uՃk�!�&��n��q��� "�E�q,sM�Կ�L��	f���*�A�#��uE�/�/�@L�}��[�B��ꍎ���Hي����1SZEY,fB����S�~���Q�H�)�s��m)�)K�ы�2��M3u- ҧ+>M���Y��3@YTV�|��)��y��Ӂiǌh��Q��$A-�w2E	Bp�꼖LɊB�����E� �϶L~����bM�8S(Ԕ� )Qf�*�9��񁯽��7w}���R�2��W8"B�N<������nM�d�6�M�@�V�Z���u��c	�ZEM<��,Дi�����cKs{t�� ��)�94��#b�V��h�w�d	���L�~��h8B�9|�1
�Ⱥ�{�H�Ѥ�~g[@d��RD}����n�ZK�O4)B��):h�fL�8�J�W�r��`��e�߶�R��M©�X|)m4� ���B��tjQ�O
�f7M>!�pV9x�����IK��ث��DӚ,7e��ĩN�Z2Vzib�@˟�.����R־�sȁ[�K���@:]��Jo	I�,8�km�&KJL�_Q���ô�3g�\�FS�!9|��q,����͕��;�8�#O�F*�%���
+'�� '�J6����RP�˰6�Ӏ(�P���i�
D�\�!W�-2)݁e�X��8B�!����3��Μ�ڈ��δ�S�X�����Ӱ�A�cl9�|���N��[]L����5< B:ۺ��_�� �Bd>Ӄ��FS�z�㗨�����1C88,�6�t*�I\��0��U�åp��*q�J��łBȔB6f��.��H͠�pBL[�)�����l��Έg��b8I'� oQ+ky]p��V�ACq��9KO�W�*�%}� F:�
�N U�bS!Yj5~��[Q`��[�%��#5��+�\)@�}�ѝ�D4����Z`c�)�#�M'�B�I�i
�f�V.��6!S%K2�p�+늉Sb�QKhR"��c*GzH�bE���FkʙZ)w9ZE!�}'�d�u���b#�L�~X�!�*�h���W��q��@&�&!,�vs�t�Ô�jF��v�U{�ms0˥������2��P��Ǉh�t�9p`NuI?&B���&�i��B(������5�K�K75ʪc���Z��W�f��$.��/sD����H��lQ��($e��,��Z� �S�%~��Uc��b�©p���N�|�q��}�_�rF�?S�4Su�`�S`L�ׅQt�	D#��FO�������d�[��3%Tq� �ߒ���wъ�E�>'5���1'��4�A��)DJۉ�9p�ƖÇ�͔��HE��T���0�@V����ԭ�*,2f�ՕiY	�1���Of�Wf�@�'g~��?[�'WS��/y]�.�*����̓=�W�O�g���o�إwE}�b�T��������{�i�����7�SHsOM��vǯ_���98��쳏�����O~��7������o������ݴ�]x������N�<����{;��7�*�����bw�w��Z���G����!��׍m��UQ�|QN�8�e�E���A��#wf��8ԺQ�d2q})��%btJ?�������7���ӛG��;��gop`��zNht���d�U(�72�G�F������O�Dck��S" �JFm�R:��(
�dq�r �󕠙���AΤ�F�W4�6{�驗O����;6\VOc�,�}��R�`�6A4�[��
���q�ֶ�@#�������(!�qݍtL�t����Y��YL��5�p��cL�ZZ��Y����~ �LL��^?_KDNJ��,Y]�f�p�Cҙ\S~߸��p���7�`L�rR�I���:�lQ���4�䎸�Δ�lDvE쒍9~p��^����}��?y�/�}~�=.��p    IDATF���r��{|��@9gȧ��.N�w�No8�ݺ���Zݠv�пj8��C;�{����������������v.O�w������7��­�����;o�������'���N�3�O�ѹe�|��тwZZ�l�c-a�S��M�H7��)� �i*ˁ��å��;V���5`:��a�x��y���(���(�E��:������Q u�[��� ¡����Z֫�(ʊ.��>�2u�86A�pΌ�*�cLG!d!S�p r��] 4>G!#<$�h�
R����픔ZF�H9R<�k�l�����ɨ�0���ߑ�#���MMQ�J�*r�+���Kq�<����T2� �`�r#��d��q���9MW�3;�/] ��5����5z\ΜZ���78�NK%V��B��%��QY)��������p���i�@�I�tn!L���#p�1>�hK�\3�.�3��s�z�Vujl��`� j�8�Z��%i2VW5l��J^���3RVg�S�t��+!�G�t�p�,eQ4F!�.���r$"XKɡ����K�,S�)�gVg[4C�aZNK�����T�t/[�`�h��2M)�h��QE�^R��P�����<S����DS���p��g-/%
���x]	���J�Ɉp��ƌ�284"p�@#}�q8���*��"�#ܔ�a��~�gRp�|����_z���0#b�U_�~�n
e��#�!`�%��|4<���	Y!F͈Pۺeȵ�D1����/�r�ο��/~��i��w��+�Ȓ������k��}�U�tR�F�:�L_C)���N�,���HYe:q8ҙ�p]�±LT�p��������Gֽ�Hz]g��sֹx�DI�d�:X���1`�؀/�@���?�����f ��c [�x�jɲH�*�y�sUV�)������������������#2�Hjhg�:t�ѐ�yG�O��ڱȊV�/A
-�_"�UG6M�NM
�#�L��4��U˭��(|;1_!8�f$1�ʲcфLë;����S�G:���J�q!~:C�T�T���V�l���R@�������oF2�J��T��"�CV���D�)��U�7�+!��O���P4SdVM�e%F��R+-�t�u]�J`�k;f�>q�d����� 
�QӲ���HO�43�IM�8UL�5�I���dѮ�[K�4�Z��V4e�p��r����9�p=����y���I�h*E�(|:��t2��Is�!)�q�L�&+���7
�t���Ԍ�G#^�|�)un��oE��-���C.��B�Y�$](M
���B�#"T����\��+�ѽ��5�2Wg�����z�Cz��M�O�źB���pD9����9�5�i)��+�f
U�A�ReAZd�b����oD0�n��T��H��r9�zD�c*�N��nT�>W(��K$߶'>j�!���%B8dg'�-p��5��L?�@L���V�4S�5i����u�K)���!�'�D:����2�ZHN匓�ZL9���H��8��o�FJb5�F[3�5�VY=�u}[�0s�2�I-�T�	ܮ���U��RX���W����+a:��K��Q��F8�(�h%z}��q��g��QJ
!�G��(Ω[��)�.�Y�R"(��7k���᜶"��i���@c�"����jh��6K�ٔ�ꐓ�_b=����^�T���M())����j&�TI�����&�~�6R0n#|F��p��,�V���%�ՁL|��VT���&�]{�3��z� ��B��6
���L�vF�6��E۱�1���;��x�L�huRn)�ުq�V?�-�ߪ�fV�x�F!GbSˌO�_�B�F]��K�%�B��r?5�(� hB����i	p�,����Os���B��_-'H;B/6>c��5�/^��@��f��������������m�� �r��޽��G��g><	����_��xx��jn�eM�E<�P�V��T�������޼�����w�������������l���ውmܿ8=���Ko|�n�^����n������]�V��km��}��Y�n��v���1#뢬����l,����������WuJ��������
M>�5�h���+`%�]hQ��1�ã�k��?Ȇ_����ϷP>󞓛n�w���3ug��Bt��=�:l-Z�	Sh��C9�Fdc��
YB�_
��B-d[!�飙���i��`��a�_Q��4[��R0�G���c�t���m��).��v}�S��,�+���F����ԥ��C4��Y��1�����@�5B:Zht(�u�_�k���H_�Q�]�K��4F���鎜Q�)�~��ΒwF�(C�R���T�R	��&��sц�W�5'+BL>?S3��A���ij�K��B�+wYQ
��ۉ�Ԅ�mZ�>!����E�rs����/N^�s��o���[�_쭯�N��<y�b�7	����>�~r�+��;;����5�͸��q|�糟���{�l���r`N��<�m��0�>������7o?}r����t�������|������}�������7�q������&�6�7��oO4�\�v��Z[�)*��E1%
5]�����󌌃���Pn�#�������|~Z!����U$��g6�,ϐ��y�?I �!d�Y���QQ��Np��#u~V߭�/7�ȝ��]�t�\S8���%���#5�L'ޔ_9�8�T�Fk��E<Nu[ ���1���Z�)'�9)w�L�7=3�(#Kǘ�*8@|=�.�V��h��I=��»�~�u.]`
=I��0�\~E�fd��I1���	1���zvB���!:�˦���m�r�V�@4A	1"X#�TE�%Br��r�p�D� �
H��Ƒ���M����Z�@�e"LH��_"���X>rQx�	�jƇc�0��4%��#�[��k�X�Ȧu^ȵ��,����� _���� �Ti���:��[lS��09p�ǎ!�5C?@EM+mħ�Uޮ��J� �s�ˑe�p�Ҭ�����<��
�LnL%p:�@S��R�3>�(���@o	��*�ʃ©�A�]�T�Psrd��6��^
�Vјr� g]����8R�J�z<�+ԣ;Acֵ(S���4*D�1u�;���3,�M�W�@_�!��e��@��N��օ̯�VM�z �E�L�(+P�~t���U��sǈV�Q�R4 �"����8'��s�G?����������ϑ]�{��y_SR4L�͡L����h	��Yu�9�Cߩ��(��BVz#����>��F
h���U]-4�BR4`Q�5CM�Z@j�U�Ι4�(J*f�J )�)Q�Q�hj+p��a�@SY��(*}��J�H� �A:�8|8�����&j,2|,Bdࢲ�VH�Zp�0�)=R��r�Y��m����KM���RW�D1!]>��s�!٦�#�1E`eq"�Ҳ0�Oj�p#��L�H$P��Rr�
!���!E늏�N
|�h:�)|x��h��z�7�j��K�X��`:]&Y�qত(z����AZ`j8�l�"��X��9���wQ�<p���L��7���K,+|8��g�p�l�����rp�d��
ᰲZN�,�ʑ*��ib�R�i#Bk������#�B��!�N���Rr�ҾQ�d��F�1v��gM]�]����N.�iF�r��'}ϐYJ�*��!
m�Rb��t&�K�jE�����zfB�94������(F���^��2"'�XJ��#�B�br$"���BjcR0k�QB�K�m��A��N��g���H��QT-#늓��a�G���LJ"M�<%��v50~̢����8�/ڥ2��"�'RJ���AԔ�%���T���')�d!U�"B|Ƒ�4�Q����Ri�2PnVc�r���Z�n�p����q�ȶU��˟��!��('Dd�K�*-��1����X���MD֤ko**�`����Y������1duM� 24S�(��8A�zXr^]bQ�oQ�
B[��1g4�	�b�R3�(/��.AuM�u-��YB~��τ褿�-�)[�������D��H)t��r��Z"�E������5�*�+�G���%}�A��\3�J$�Z�ghJ����J����Y�B����-��\zd#kZW�9�e�j�V]�|dS�P��@���=���݌8�����UHV"�v8D���8�\c���r�~r�I�'��@��=
�8�8�hMZ��1EF�������DO�(��B�� �M�P&b��S����5����1�Lқ�&k�r᏷�{{���Z�R�ÝS�<t�����b�ly�ғ��b^,������N�/�ݜ��쪿��Kb����h�¼}���t�pǧ�.v},����:x��}������_�������Ӎ�}��������f����F����ƾ��~YG��X�b��
^=B��Ʉ��mT���@D���	��q#�����\8Y��m���<�[���9�����S�8�=�"cb|t��s�c,��ٖ8+.�����s�&�����/�C�]H˒�E�E`!ۣ2 ��R8�|�@N
�hʇ�� ��2Zl��g�IE���!?�� R��_��*a�4���\J�X�]�����oQ{Ǆ��.��Zz4�27�T���y�WB���19]eL!H|�(c�L4k&N���O�CK����D�7u��}�Mn�n�+�I�S-#��P(]cpg�'?�	�9��7*jڭ��Q��2��)'.4��h���ʕi�h!�D���O!Όj�T�q����4f��q ��Gc���s���h���]�Ev����-��`�����Yn���Կ��U�����av߷}�ؓ�_J�������ٞ�u��ͅ��=O��z�h�����sl�2���ɓ��������k��*<��$���/?��_>����7�Op�󮭾���|�;��I$�S��8؝y����-ͯ;��uq�:�J�͙Sd
��S�3����[!H�ﳊ��Y6j}��#Bc�FM����@jX�������vC��4<�ַ��]��jZ�Ό���b0�����p#��O��
y !�ąi�bZ�Є$B����q�c:�����d��3#�hr�����p��iҩ+�D�߈�ՒA�P�#�'˔��2˪�y�.9)�@!�>z��-�Ɨ���T��χ�DH����N��k�S�'S%0I٪�\>��A�Q�o�ɑe!�@��1����7E�e-�.
� �ȤpR���P�%�9`�Ͷ�&q#���r�<�jɴ�Z�)#��Rf���Y�Z�)��!JRK�JOV��Qk�'*w-��q��b4��,BL!�L��Is�A
�S{FQ�tLsp��.\��[�l��!�XFS��i�*-P	Q�k�i����!ϒ�~~�	]!L�h&}4Sj�t�����dvCH�.��7�c(#)���g��»e^�'�8�O��S�*:]�-G�J�s֤e8�����s��[ �o;�0D�n�q*a��"�B��1z����;����B�B� RL[`=C�
!����1S��~D<T����Z�X�f
$�b�
��K)�is**�=q�|"Sŷ�~�������S�뵬��>��g���SW��dA���B6j��]B��I���r1�s(d��M�Ȣ�4`��@�dt�~p$�����TKrm)Y���I�o!��A��#U]|�|1I�%��[u��d��MP4g���k�$��"J��<�m�]�K�,��Ӂ+G�g�����B��R���1ʂ�����rRnu@S>ِFL�R@��($-f�JYt� 8
����Z0�+颉Գ)���Ʀ���	�Vˊ�PkQ�BE5E(��ߔr�D���h"|�KW����� :���p���~KHH)����Ԁ�98�)��i>~�5�Y��GK
��2R8����"#Ј�TJ�G�s*/˔ID��=|b"Ԓ,~M��*R{�C�j�F���s����0kC-8���F�Ɖ�f��9���A(*�ߞt~L�Ǵ�Q�D�>�@�-s��u��hS8#�ቔA�T�h74`\ʯ���Yn"�8�U��(�%v�W���3\JGE��PH�DH=S��7Ł �ⴺ:�'����*ǯs�.M)-Dt�e�b�ʂ�^�-a[*���G�t}ӑr�#p�2��qj ��=)W�=�8؅d�������J��s[
XV=��y)tZ��f��)L��ŏ�v�(�6!aDR�qV'�R�CN�t�V�Q���ɇg�H��4+���	ԳW Vד�iKlEʙ�<-	.�A(j�,%5>�^?}LYt zC1͏�K�/�����9���,ʜ�1'*Dߔ��ejg����[�1S�7V7>��݋F�*�ᥴ.��:O��N8���f��c�^�2>��Q�H`��^V�����,d8����H)T�)+����Nˏ ����/g�̄�YQ̤��ϘJT�,�,���E#��p$�ۙ��Ł���h$E���#�)����!d�����Y�)���s���'�џ)
�HA0�"u�WQ;��D%B�e�D��ꇏ�e|#ZH�N>g~�!�V"��0KD�ql�PE[H�P���4f��Nʔ��q�����V��J̗�5�4X!��4���R�(ݹN|����R���n���	�|_~)���^����Rc�]��q�{���������m�/�M���뾄��7/}Zҽ1�?_\�3O����@��q}�ig�p����������k77�{7�q�;?z��������?~����S�^���ؽS�޾/���:��5M��]��<?wr�v7�'5}ǭ����e٨��WO�Kӯ6�3�)�Uu�z�خh��J9HB�n�pL{�e���%�K�G����+gt�����o�n��"����Ư�?��_�.������i��t��#���,�Z�P��D3)Y��pu�d1d�tE���7*�q̧Y4����t����� �c#����͏`�O�J�Zv��%v�����z��ա�r3��~��_�U� ��v�m4Ŕ.�Zu8~��T����t����@}R����c�^N= �q��r9rIiX
���P����K����[�|4� ����t������t����p`K_)W�&RDp��1C4��"T`x͗R��q;��b��M�>SN�-Wcӛ���G �C8ʞz=�=;=}v�㇞�<�������?��7�ӓ˃��c�3���ή72/w��?�s�����K�����ӗ�_<x�*�x�ŗ�w������'�6��S�?x��Mo�|��G���W�>��y~y�������~�w�u6�dq�<9X�3��!N��Ď
��u������i7��'�Y�,6dL4�2���M�1s,=���^g�lGQ{ޅ����>��s~�Z�1ݴ�9h%�/�����:Pr.D���0! C6�N���n%@���@#Z��e6�oB*�e=�i���7��-s�l�cۊ(H15ҙ%�U��1ZT>����KS��8�J7
�|a��)c��2%���q4���E���sdiF�Tb�YWJ�*�mK�A�\`�U�\V+5���I
R��BV�Ț�iuB�p�88ɦP�����7�MqD9Ek�_E>M�hrƏ)�,�,�i��gy���J��[M�'�ǹ��f��v(J��K� j�ol�z��tZK���f���� �c*D���!�5o��`lu�tp�,<|R�E�A!~_�۴m�zM�OJ
@���Z�B@>$gV����\��UL�~ko��$��B׆+�:
A&n�NW�����S�~���^iO�|���"E4d�B{��2UBEo�1|8�)ԎU�ȶl��V�̄�8�1B�ߔ�յ��hҙ�1�Ƅ�!D����
�m!(J�*,�o��oE�~d��r2�(�*T��-��(e��I1���U����bU�d����cD�B����eNu!�LE�]q�Z��h��%�{ݐ@��c�:��?�����������$@ī=
á槧BD�Z���Ǻ8���-j�FFM�����G�X��    IDAT�_��(���NZ�F�Q�v�+Ec�iR�H����j��jˁ��gEӴ�pc�Dј��	�&�O4'P�H	���un�M�� �������ˊ�g�8Q�|��R�� í=�8��eI1.���D+R�1���x��V�W��mQqg-j%N��&��2%"�U������Xc�����^�љD���e�$e�D*hZu`�ɒr� )�^��է(?�>Z��vFz��N�*?�T+�~���ʖBd�$b���fp
��M�sI{�C?�E�F�\|��*f:-j�M�9J�LѐJ 0xӤ�%� rpj�O�/eh�Bk,T�Zib�B~�\>r4>�Q��t��,�_�iE�֕,�|�� rk� �Wu-�9�� J��S-k4�\%�ٶ G�âU�Z�1������̶Bu�T���j��ƶN�f�U��J
X��M(Z�Ĭ�:��]�8F�Bt�(���NќQV�壕>Y%S�#S�i@��]��{V:gV'*7#��1�khL��0-�,��RcݱVQ��0B�`�G:�F)l8�	�!�th�tY��<`!�mKQ�
qt�#�M4�$��F�&d�5L����vϸj\鴖�hj�|�]�q��х�^��TB�	���	͚4B���@�� ��4�.6q#3|MZv�n�L͸f/:%"ϳ����nHDN�#�,"k��ьcJG���Ƨ���t���1Rnc����ь|��L���!�S� ���ׄ|4Y�Ӕ��U�P�)7�K���_.Д�OKB����VZ�tY&�"SNL��"�U+$��p8ቄ� �_	c�5� ���:�fL��҉9(�Q�r��#qr9��*�Z�W�B���0��1u�,��D=@�rBL�MǙrq�9�X�^"��)�uଗ�9�3N��Qb�~'{ϧ�)-��.�*u��V���ʊ�c|�*�4m��8Ƥ&d�|��Nr��rJ�	��ӛuɢ�\3��s�՘�Q��A��8����M�B�:㍏����J���D�?�yy�-P}���/wv�.��&G��[.
;�1v�(;�2�R~Ix��_���|�����=�=�ux���ᝣ�������׮�zx�7�><<q_B�;{��/�ͽ���V��۹y�����>I��8􎀏2.k[��ɪ٫����l�����'�v����5'2	�s,mԿ�ۿ��W��_�k~���h�/�
a��K�3�L�ap�dq[�'U �G�߸~|��]������6�8yv���)d,�kD\3s�MC�-Y-��|c6k��;jB�W�`9ަ�M!h|c`S`%R�b����Ù��ub��l��(O�oo���H��,���a�:��=q;H!Y��Vq��E��O����F�n+���>��I�ˍ_�G�B=69N_:�µv�əV]�q[S� �s����z�;r�S����#NP�V�M\R�.�<DW�n��5 t�����q� j�	Ł��(��;�%%��늯%�\Ƒ���,}J�3��rÇ&��4�Rr��#��e��z��ݮ�����/|�O����ˏ����|��;;��v��g��<�8|N������K���l����O���������O��.��>�p����>���/�����U���?�XZ8<�x�Ƚw��s����o^޾s�{yz�3���7�ܼs��ϒ|��r��Թ˭U�[��Cckl��KS�¥� B[vj�+��E���g�CA-f�w2K�]���z���i�w����\9�~�!�C���r�{�eu�i��\	$���!�CT5�@nZ+���"H�0���ں^!���)'A�<n*=~��ч34MV�s�fE*2˔Ai�tF����h-�9r���a�(#M`QQ�pF3��X�|M"��̇CX��[��m�"W�'������bJa�o9��Ww�hi5)��V�ܪ��^d� �DM9霦9ԒmZ0��uH�HA�������ᘲD��p�|�����t�!��C�b�S~���J@RC��Y��p���"$`=��L��)'�V�_ᘖ;��� m�M�ɯ=���j��dvRVWV#5��T���@Su9l�!eH[*+r����q��R�B�BD#sZ��j*
���y���y�#HGcFV{�&��۫�0={xM൩PYjy.��쵂� ���R�o�nd4�ט�&�J�g�	iMYL
@SL�� ޺t���Dە_
A(�č􍬵p��:�#�qHRF
t���4�@H�ρx�r~n�G��WZp��^�<R��z 6��ѷ���nJ�)�@�~z�vipH���?_�tY9|&׏F`ꁹ���П��v�}���<��2�w�}�;��X��
1d�/��*ǆk�;�j��(�7�6�f�t�0����:�����������I	�{	k�p:�Dt���0�ć�Jg�L��8) �P'F`�rQ>G	R_Yc��BtL�M�:7��
�O�\`�z�"�X�!�pX��i!3��7�7�����di�P���JkݦE�JL��P`V��*�f)NNͷ�
هM�d��)�3�K���!�Ƥ3`�Ygja���\.q��崮[6?&2�4�hΧ��E�UR!���T��8�*��@�\
���"^bE�dK��,s���4S���@>>&�w�9��T!H��B�r�Y�  K�"��Z�B�L)���p�Ħ9��N��+WFfg��U�j�)�SiѦ��Ĳ�_Q0m�����q5ѕS�_ֶ�Y�F�r'
�|�{9FW���GS�H
S>�!�T�9��1��L)�eM'"*��2��i����D�h�USf�s�d�N�ܪP��SS7B���Z}&]Ԕc�c��e�Ē�.\c�-D��$Rb���K��#�g�s�F�5c�s�,:�;�l�ԝ�����1����8�E���Z�Q��X��U4��/��k�ZD%��2d����U�ǁ�U]S�����C�B8��v�I�~�xԌp`�T1�z4>C�{�jM(r�J��B|�8��j⠙NW
Y�Q�����q����W�NL96�q����hD���ɐ�E���M��@�B�KP7�/:jڀ�q�ā�v�K�Im ��V��[c-M9 �r�fVu`�b�!>%Z�(5��E)ԕ'�)H��˵.��T�uā�t��{y\��:ǩ�8�j�\~=����%�XQH]U��zF��'_nHu)@X���j������PU8E�:��)����Y�O�6h�N"�+Q�3�U��\r=��u������#�.������p��TP�_"bʑޒ�7�ߴ�a�����PѴ�>S�8��!�J��&'�V�Ռ���r8EgQ)�ؔ� K�U���5�8����0�����oR�����,��Ҽ������+}!���ő�`�������������������/�XJ�,��\��%=k8���e��}�'��n�:�λ�ܹ�t���;����������g'��[F��F�7Au�W����nܽ}�����3�긪��[y���m���ͫ��E�a|;��0�������@��.��x�����G��w�p���IA:��nw!0	b~���B�巯�<ܻ�ڝk�o�<8�}�����WE�6/��ݷ�_�q�|�vYAG����fjp�d]��1��;'Z�Ws>�D��Ȧ����`AƷ?Ff*� �0�mH���7�
�(�-�z��i�lEqD�h)���]S�Z�۷V��ti�̥�g� ��\57���B���W�����n��pF��)D�MEUj[�^�5�emE�A�%����>�G�O4���7�Sj�ҿ��o;�
�u�%�a�kc!�1nG��ٞb��}�*�e�1#��脦.�Ʌp���6p �鏿]eB�|V�!O!����D h�t�q���G�?�ࣽ�_���[w�~x��w~��;����[�.�/�>���������ų��'�?yx��{p�u���w絻��|r�p�G��ᣋ�O_<y���#��ɽy���˳����������ypt˛wo8��������"�_|�K[_<?�CJo���9d`��U��-��9O��x []�,���QG�(jls�U]n)��b"�w�yG���o����4� DcWO�αU�T��Q�*a[�L�T�T8&�)���_��2¥0Q)mG4#��V�϶q���|p�(��LYTV�1��G�-�A6��"U������-�=�W�>�8ʣ�&�b�X&f-�3ܴ�ɀ�3�g��0+��S�& 5@ʿ*]G��h�/*�B�ch#s�+�Z�B�"��1���#j�g�PJ �h���3gMZ.w`R�cj�0'��LJ��E�P�8�	y��:V�d�
!�)Z�Mc6%�1� ���ۓ���-?��ڨ%c;\��=�J�C\J%&�>ј,�L�Bn,��p��WȈYz:r���f/�e�ZH)S=3~�.�A0K���*7Z#A:����sD�����&������ 7�X�M�!.�'n�Ky7�N!mw�(0Rp��h�^� S �D�����������?��k� ����O4�F�����=?�<��"E9L#Qms�	�(����Ln��V��j����j���������\^^#�G-&Ŕ�����qH
n�������-��#܋'�^�{������!خ��CO�	�!�B)��2�x��2��g�gv�׿�5��ǺD�2::ђ%h��y���G}���R��?�����j?;~��i���ƑH����N�c\��b}í�,m��Ȥ�p �9�Q���e&j	p�cQ�T���o��v�Eק��^;�&�H
�B�52;LY�2�T�K`���*�M?�/��k�VWɫ�<d�8)�E�V:�kd!jU4��%ʂ�9�|Ʃ2?N��A�F��@�%�rf:�R.hs�rY���ƌo9h�Ʀ۴z�A`.MH"��K�#K3�)��z`
I��ʽ��/E��1�f���]����B�jڙ)W:���vuH
�B��Ó��h�4QkMm�X��rBl4媕P9)�8i&E�������MKlJك�Z!4jB3BXYp>~�R�2�����f�� �����&�Y��`u�qڴ
1"eg+�*��*#%��3�p~�rud�@��(��1eBU�EY�Fѐ٨�F!
t��z|~ju��1�9R*Q������q�X��!B�!J4%���I�@f���g�� %ℛF32���Lg���*4� d�S3�-
�m�_�'�غ8�Ƒ��ɧ� �γc�4�y����(J�e�!dUZ�କ��_"Dh�b�M(����O�pQ���ү�%V}*Z�}�^��ꡥ�+g�����H
|ʌ#����o,�����@�P���k�����RƉ�H� 0dS|���/
d|"�C�,L���Ȳ�����6�ϊV��C6�I٫���b1��d"eZT-ߘ_T(gFp�*�l4:mu�B��քT��&��m�(�0uk�c����رB�7�A8��,Ĕ�0NU�ͧ�bW�N��X'eE6����D�K7m1Y?
1�� ���פP:����:��tc=G�@.7r|�ąRFK�T�_'���M�]�D���F�"N���8�V��	��'B}�,dL��!������qZ�*�h����y�O�q>B)FS���fcMS�`v��B�����tl��]_�,M)���Lh���.e~�FQ����_:?����*U!��tS8�1�Su�>�3�_
GhDf�H�K!6
Ԥ�`��ҁZc%Ж��O�D\Qc;nd-G�_E��hB�T��}۬�Ç{�ӳ�Ã�_B���Τ�/,��{��\��az^���x��]�0�w2�+��[k}����Io�کec�v��o�9~����{�9��|�Ń�����~����G�/7{�>����پϐ.���Я��ƧG����������WGn�|uk�rf��I{ȱ]Θ� V�	g�˲k�c��U�n�G������,�P�Ū���I��M��RS��Ӂ`��Y.�Ņ�n&�w�kB��O��g2�.��^�]������'�nd�-��|lsytp��p��.��������(}�UF&�U�]? 'S+�)�DN��!L#�tJ��1���zx�7-�B�N��$�~��	,9<�/��$�:4ݖ2E�pLI���G���ApMK�s�Qh�
�}p���,;߿n����%OV)W�3��H�����p���q�ei�/�~3QF��.�hޛ�@$�G�BJ�����ݤ>��c_Q�ID�8|R�J@X�g�q����N��
j�猙��t�;	�`Z�� �������ĉ�x��~E�yd���g3������#(��鳳��}j����8���?���O��;o}߁�~���䥯־<y~���G����O����ݾyry|t����k�ǟ�m����ɧ����O.��|������S�����鳽�>�g��{��k�|i��7_lN����ט����ɗ��_��<�֦����&ɽG�Ɂ���8�;�v̲ �*�� "@hv���z��
9~#���B��Dk�z�t�M%�R�>=Cjr9ܞO=ݢ�O@����;��V��eS��E��B0	vM�Ua@#��hf
��6(��(��g�6�U��t�LA�v���Vʄ0�JN��@ ~R�xU�6�2>q� �!�[Gn�,RƦrqd!,��9ueL�6���m�n��M
��mB�*�Ώi�pj#02D��Q9���L:�&�,����G(5
RL��c:�P�6>���ԡ�4-�/eF�/�c	���߶8�t�U���ɛY�=)8c�����g5�?WG��{���z�_!�t����4E`98|��D�5��_���&*˔��Ff�J�P"�N�)�k s:Y���ld��9PzH:]�J��-"�V�k2�#����H!��5ռļ�h���EG�pO�V'��8���K�O��pZK���t��:� ����*�-��f!
�ZJ��GE�K��'��)�gO�>;�U��"tM�(���B�2��L��_��_��_Z���D)p?E��[!�jɈ �߿���@�Z��I�j5=x-������y��~�,Ej�(}vے��u���1	���?��?�#�W���w煾���3
��>��8�������Nz��}M+�&���wM��D�QNk�����SӤNLUl�Z�D���s�s,P� �N��������H�KF.�t�(���.�UX��G5����O]8?qV�%�b�/�2�4ρ�'A�1GP
3��m�9>Q��V�Vc�!�4� ���V���:�4ű
ά%2�huo�FQ])��04V�| B���e]U
��F�5��X�����-R�E[z�� �Z�᳢5��hL��1
��B���|���kO:?Y|F�h�Cd��קnC"�0j�e�"Y;P���r}� �B8��'}#}�����2�R���J��H�:�4QVo�����+k��h��)Ӕ顮 p����B"�B���q������ђjǄ�:T�,^�NW���+D�%���13ʜF�*�k/B�p�:HZ��ʯ(�)��@S�j[!H�`=�FS4�S�� 0��o]� c&+Z.�I���r�ZV4��۱��������Y8@�������qШ�hh��FS&d,�~bBp���4�H���z���_.e6���W��¯��i)�j,NY#�0~��2��^�`	:d�d%��H�d�Χ(�t,Z�� )N�U��L�T=��\.�ҳ}��d9��I(��8~�m)!&�#W9%�p � C0��g��>>��\���u;&1Y��,�U�K)���2��OAb�)�,~�B�@� d�t��J�"�p�ƜBF���|RR6�)LK�z�duq98Sq�IA�#:�� L�$�j��G����32-�|�}�������t�)�&$<ܴ��0�N!�HU"�2xLH]�o�_��C)	
�0[���N� �J�F��S����J�5 4R@�Rq��Ϣ�^�h�oU���5NV��N��U)L�8�1S�T�Ǆ�;��(�X�� >�i���i	1kAt��^��c��j�I�sQ�[qޯo�s^��q�8Lb����E@fjm����8s    IDAT�L�B��=*��֛��-�y��6���]!�R�+>�i��S�D j� d��&n�c�nU�����T�Dc��{ˇ2���p�U��R����d��~y��=L��>�ytp{s��ry�m�|��}_�7-w���y��/������Ã�so�R�8?;�~��bsm������u�g�Q�{?�>�������?�����Wϼ�w�9�Ƌ�}�m:�\�?\���9O�>}p��޵�͡��yz��`w�۟�̧7g������������-V�u�Ff��lB'�?������\� �~1�.��!�������q���;	�M���J��>�����O�}q�K��o������/n���y��OμAb�7{�>�{xc�`�C��G7�ervyx����ϟ>|���T|��[��Y�V�����.��hQ�uy.t0]vH�Zr�M�0\��v�H�4�g�!���l%a�JL_�D`�L9�T4�h����lg�a�aF�v�p᭎˄�BZ��ݽ��W�Wn%�
��܈3�����c�$e��F�D�=cT�Q�9)Q
���4\�Fӹŧ�{�pdO��_���I�R�����NDoh˦���e��JE��m�5�&H�G�޽h���9!��+:Y����U����)[G�6�pX�r�@MtD���v9��.��ZpQ_dv���ã��ӣc���/w��ᣛO�%����ً��Ƀ�G��� ��OO_|y������э�'��=x������͝=�9X>`�����oܾ�����>~�������Ӌ���Ow�߸}��5G����g_<8:����^{���G�7'����>���}���=?=;8:��On߽�I�!q�С�/3�T�-�Y�uY�:Q���L���,��)_��y6���r�@�Q���r��������0�Tf�xLQCX~v���0	>��-�҈�X��|�z�(T��6�X��0�[�D~��`��P��1�,ʟ�8���&}#){$Z.�n��O3��BF䶵�J�^?�򉫢N"�4!U�h~:|��v�S|�Z|>g�DM���G`��:�)G�ȍin��� k "��QV݊愈VѴ�r����mN���q��@#K��䳮 ���)T"Ĥ�0B�A�.ҫot�}���ސ���2
|�~IV�9IMJ͐�{�Ln	MtT�HV!S�G��jg	_�K ���L)�V:�����irp�re�JL��Q�u��=_@��iփ�)ksD9�Y[Q��׌���)�d~��Eˁg��$U��iM#h��i��j�Z���+�D{z�?-�D@+�b|"LE�~xR� ��X����v��W-h�F]A���4e��A����)H���r��B^�8���lJ�N��~�;��%R	!jhp�F��D��vh���8��l�!�������~`E])#�DH����(�DL�ӈ/�
����I{� ���ت��o5Ec����[�����c��8:�ʛ�~2�(W��Jc"Hט_W:����ZE0R��4`ĴE|!����D��&-�x�?��{�&K�h�(��v���SW$=��q�jL�͊������%D���:$B�45#�gU��U�J<��ϡ����-����P!:��h��d!K���Y���MkҔ�,�XE����h1�҄��h��"�cբZ5"�*�l�J��%#0r���zK9آ�J�6"�����K�g���1�K0�|���(�OGc���@Yl�g
���88�����Z~H�L&ߞc&%�C��`:e���9���zW�d�M�RC�� !:)� Du�3�\~j|N�q�h2����r�MѶK��XN��A`M����n��0���[��q�N��PUj���	◂��?�4Ɂ�T�t��B��b�Z���sT�c���iOBDo�ل��q��_��	4�)J��GF�S6B�H�Ӟ4BD�qX0e�I�%��j�S�k;W)Qֱ���4ܔ���tv����'��aQNp��g����1���o*k��Le�Q I�B���-���1�*8|��)AH��sD{�	����KI�N,g{��������b�Jo(Ϻ���J�	ʍ���|�:���I�����Ȅ 	���R�z�i6�I7�j A:S�m���Vh���N�_-;�?�|H!~N䖙>\
�$Ҫ�UQ
�ڈ�`:�p &�ն�4My��N�4QY�!��v(a�!H/��Z50�3�� �G-��
u �$E'Y8"Bh�qz��A0��h�4e|�YӪMDfړ�U3�a�hM�zk*�4�F-A�+�Z���l!�]I��4�5���?���xeዚ�D����d�YR'3�hx��ث���!1ժ�E}K8;�Y�բ�aM�:�hLԘG9�4��L'��\ G�t�h�uI>|�".Z]~j��Ï�f|����/}~â�Q���zK_"G
g�J�!wh��8�fR��(�ND��'M�(�)��'���å���j���FӲ��H���m�"�o,Z�v3�F���xc��meH�e1`r�"�>Ź|Lpwχ/v.���o0�=�쿸8ۿ�=��NZ/{�o���g�6{�*>ǵ��O�O6>��x�z_�5��wz���7�p���`���'?��o~��}t��7߽?�ߪW}ii�գr�w�^�ؽx��:���]V�_��\�ǬW�ؽ���[H;`\�ru[o#���	h�ܞ�α����Ѣ~5rJu��!���~w�#�v�x;$���O��FYǇ׬�p�����s��qx~�痧�i�؅y�y��v�wz���n�H�u���q���O������G���^�}}�W���rT�׋�3�f��U�;pu6f�B�U,Wu]��hr[�v�Ъ��X6`�e�!B�h�%̚��d�SH�T�q^�-��V4`"��8F3�=�p(����t�U!���w�y���\Y_	� �������I��\R@�,�rJG�����m�D9i�M)`�����{_�aRP����T�Q!����Q��ٶ��H4%
��ls�[�v���2�����Et�J
�>�N�X�!��ˊ؀M����7~%��pr��m&_.�֭;����u�޶��v�:��<{~v����=����������_�=�|�ؓٵ��g/���_^>�\������"����D��7�������o~��ݝk��ͽ׏w_���<~��Oq�~���_�ڛ�>���dgsv��񵣽󓇞��v������;o�u�gAo���W�OsY��u8Ξ�%��؞X��dg�Eh+\`>|Br�iOzΞ)߹U�u8��ʅ�vn��#������s*��|6ŝk�����4R�%'-��v!F9>P�#�u���1����5�j^"_[g�R�@4
���Z�Q'��Y�Ȧ:��R ���h��
q�X�sBj ��oʗ�h��+Q('��*��)e�p�I^z���Z˜P�2�FHQ�t�+�r�!|�eيt���o���*a妏)KK�����3mQ�,������E4�	��`�}|;/�H�q���4����d=������s.��?6gγD��
~�QF�3��!˥�>($��u%�B��P)�-pVJB͈����Bd�%e�4��bM��HRJ�e�G2��7��+�[���B��QJ�&��!LQ)������PC�&TRlf�8����EdՉ��R\2W0j���� �
���s��؊�<���^��1���hR-���r��2�1铢���W'����T�ޏtJ�֫o�9Z��PX嗫\������4��U��^VJP
�Si�3i�e�"�ǚ͔�eu��b���C�!2&P�^癶KF>SN]�M��.������*Y?�����J�#��~�3d�j@9R|;�	A�t �x�G��	׶�ju�������'F�R{��D?V���9<�����M�������{������>�I������1Հ�8��j!{k]k�'�׿B�J1ZE{�H;��[5�25�D"�.Z>��h@�� �e��GJ�
�04�4��I6�qj	I)+Z����h1'j�>'qH�)�/�c�f
g�䚁�b���5�D�)(+f�٫RZHkL�f 8�|�$�c�ܐrk^�,>pYث��	Ua%vɐM��D�B"5%�b�F~��ƪ����Jѕ�m'�J\dE�KB��G�B�Q
��ob���1E���J�k�S�F�:���A�4߈�� ���_�D����X��q䦣a��J�
��#�U�`Wq�X��]�D�^#���u�(�d'Kth	jl�P"p���'ĈPM2*ԛh�)\WR�
���i����F:F_�F�lD�3���?�@��ho[�Z�j�9�	��P{�Y/�E�̯4D���a���XW8���cd�m�r�k���^{�8��J�W�h'"���k�N�'%�/47�Y%0�I`M���@��:�鍯LV��dZ��fE8Ȥ���O���4�Y��9L�H��t����pXj��#%]��r��p�;*K���["#�Z)�U�d�V��$DK^�f:�8^��1"궽|-�8F"-GVS)4q8S�*вz�/��
�ȭ+8$�hF��	���^"�ҫ(E	!�UDb�FLS�����V�6��JJ�@QS��ϊZ��(�`6��H�檴HM!8&�� �zM9V'���|rQ�(���V��K�!�8�)4�(= �雊b2�NL��̢qf9�`LS���©P-�B�9p ������n��"�i���2�h��1Ǚ*h����T��t���M9��M.e�j`����a"�#ė��y��ʍ_	:53`<�v'*��R����W-����O�=�!���[�*�l��hƁ�%d�|�p4L&
7&��1b��]&]JQ &�HH�vۊVQ�տ\j��)%M4ζD��۹D�A+�xͷLQ�'-�����_=�����1/}r�{���]����;���ܜ�^����L�tA�{g>.����g�G{�G&��=R.��I�q��!N��C��v��:|��[�|��O��W���Ͽ���3_w������ιo��6�oe�v|����[g������8Y������������pzh�����v ���k��u�W���.��6�����?��_�Qw qd ���B�����)��[
����u�������vd��s�g�솽H�)�6,��9p�F�(�E=���O�s�*�p`�$�[[�b��e�Y����CQTՄ49�7��1�kE�Z;"���w�o�>=��w�{p}z���Vۿ�K=�.��{7�'.g'����=��S�G>����'ק;��Ҳuw�w6���u1�w��;�����+��14e���EE�jy�Mp�yh�Z��r�e3�"0����0d�[���e34!d���1D�������"�)�,4�8���`4�C�������n���-�-|[¦�	wcJ`��&��� �WT7�eE�+�	�	w?J^7�ⲯ�Lͭ!�Λ4�L_ P%�2�b�f4�R�ݢ1Z��"�ce���D�-d�/׀���p;Y�66#�ʋÎ9�)#$vQ�!{[RmZ�Xp�J�#r�^%�����7�=|��������n.�_>�ts��j϶99>:�<9��$����́�ܹ�d�������/=|��������������>�=�>8�������Nϟx�_�<�����ݝ�������ރ���o_�^<v��?�����G�_Q���O�/ߟg3�$�H4���ծ64��"���e��ps[��~��������M����P
�cC�"��A���O~��rlW:n�:w`�~��-����|���ޔ���2Z�&9=�y2W�j�"'7��UDl4���|f'*[s&+ft��d�Yx5�Sf�;H�%5�t�\E1���W�#ņЁ�,�B��d������Ȫ
d�jEe�窤ā���"Wm����s�1��b��S�x)�IQ.$0A^D,��\�G��!�����p�F3̫�ht٘U��߾a"���;���<@mX���lSq��B��E�K��ɻG�+G'����C�^�l3��f�)�^���Q���\z��Bؚ������&�=a6�2����|�����7��3"+r4�	��l"��P�A�5��dpYvF�Q��7^I,B=�W==Y [^"U%�=g:�V"j�"�"��%5#��;j��E�r4}=�������9�rQ{��:锚-�I��n�����.�le�K��Dޭ*O��
�(D�`�!��ք�hy�]��ۊ\R{~�yC,����Z.)p�d�ZF8�p^�!o�fj�ȅ&J�z���[�Ѥf��]N�����+�zV���k8�bѼT�e��S*Z:�/P�JL�z!�xx��\�#Y[¡�~�Pt*^j'��W��w鬧�|I/YˮW }���K�����!ġo��JA\3��R56�d�c�
t,,2�(;
��*��)Fjs�Ԑ��Ql�Y��E�NkK��	a#0*[xj�e��,ldW�]����zhv�!�#����bf�1٤��C���Ѐ�x���7�5�R�E�04j�\�B`����\[�z-��;�R!�l��V�s�\wo{b�d��x�UH!C"�Z�L��MR�B�Ţ��!�������+�V�7M�&[v��b�L
9e��,<�(`����W p�Rp���{����\І,<���h��+~��dŒ��\�;��ɋ�&��"X�t�ľ�b)bm�?Fyө�zy������+��T�B�C�����`�~�YL��%�ٱ;)�2R�(��D�AF�ՠ�+)���я��7A����AmK���Q����L�SO� ��T���luVU
S3/�- �Y�IX?�h!nGYdL��f�QIVv��4��iH`�����Z5�zR3k�M3�
����$�~�@�FP^A-C�CN_��-)����e�R@褉�0�ŀ�s�2���r�+ �fB�C�ó��Q�U�준���
)]�~@�	��иpZ�t �-�\�h�g;�E�H�k\@65!����q��T��հ����[�$mXaE���r�3��ˑ��VF�fas!��s���g�&������Ų��G��)ŅP,�kĭm. C?u�LR
\s��'$�����j6��	���[_`xC�(@jIeKG�f g}�4k��p��'��(�4���Y�5LQ:�a�$�`�nR�ٚ\%���*P_씊����(�2���`�7Y�41�yٹ�M�'
MT�X
��[����[6��� �$�B}46�t( ��{?������uD
g�>�-�F�Pch@jEE��C`��%!P�EbX (�H1 ���� �AlH�fw(��<:&Cá�N"jB��BB0�����BBxټ���+	BA/&׵'�;�1"�>~�<�fD-�ִl�g��x���rߟ��{���ž��v�<�����������HQ����{y�w:˪]_]�m<�\~���7#�|���|����_��b��"Y�Qݯ?��,���yN��g8:8�cw���oNϮ�kĥ���e�/��a�Vk�|�6SӌP/�Z��5Pj���;��f�wq�F�eZ���|nOR�Ew0��oӏ�P��/~����u������';�o<\���fs���ʻ8�\]��<��+y��r�h���v<y����������}���/��vx�xw���������ӳ;����ƣ�+OKֽ��ɍ��l����3��;�g}��Q�5|Y����/���͔[RC�bq2#"�&�˨EXr�	�av���5����+,�Թj��L,o�Uގ5�(��|j��]���#�M�x��+�л�cʎ��U���hzMF���})w��?�P�@G ����>�Z��o�a��w�HA�@ek����8�DcЩ�0�y/����6"��!�s}�8=��IjM���i��d@�\���'W5�5��5�(�2��3d)�>�%=�������<�Ŏ����Σ����s_��wt�r����W!^j\-.N���;��{/�,���>�����W^�y�g������&w�x    IDATgOoο���峋'���_<��y��ȗН?���������˯mn�:ߜ��纾���������o?�����������
v�ӍP��.j���U��Ms_����l���cǚ([ED� �zB,�F�li�^��QU�X7?e\�%���{�笐F �]� �HZ&1�j�"$%]�!6�@!��Nv3ԋ��
��PFυi>z�0����qF�:�)����g#Wv �3y2�M���R��3xx:\�@�[CY�>���ֶS�J'��(F�ʕ��\!���ͫQ��)p����� dۅY���R04����a+)D^!8�K)��nq�����m�M��6Q*L8B#4t<z���6>�#�5F��]�ly��zR�Ig��0������|1S./�^"�^�p���lW+�=i��TC8[U�r�+c��0��^Ũ��&����h\��ḻ!��跗��?��ZK���D0LYIY�A����ĄX��Rs�I�OAO�����ǑAH���5"��#^F/�L� ��?��� z
e� :�q!hC(e����y�^Uk��噡�YӴ�Y
����ѐ!���!-��$M���b�Kd��r��ThH��������f�КD
����x�e��7�~�����D
��+��mE.T$d��&�
V�X�b�6�!��%�b&�W8r[�T"jz�@slMw:���2̑�NLC����2��oh����#A��>0��N.�>��ƲT�%2�����}�۫/>�
Ճ�����as��@+�j���*Rm)���pL|L������%��_�ҮƟu�+��\�*!�"P�J� ��D٭[�C�bÑ�N��,rkkH�h\�T$�7�zd�׆υƕ�gk1��f��E�4�Ԇ���,�!eO$x�L!~=��ˈ�x�,8Cvǫ ���doW���%E���5T�!��8lR���~���BrMxI��m�A:vM
�4S��D�3�֏Ԅ�.�EK�@}d=\�VT}����ꕚ���M�P�1ve�둹f.��<G-o�	1,$W�B�[6<���Z!)�G*#~Ŕ=��h��e��jA2pحC�lH)L������0x���uf\�_[�Rn��4�zA:������Z!22��83dOk"8��w�dC��N�(��Va��
Hm�hä�]"D�ۮB����W��v�T/��l^��W�%�f� �����*����p�$H�MDs�s�r4�F�SmK�����$!C�k)�	dL�*�L�Fn�&/��VԤ� \@}"m*

 VFe���#Gk88&5Q��SyI*��!2o�}6Nâ05�f�U^��!i����۹0os��~���!P�*�,��	2�W%ˀ'�S
}��Ģ��M��h�\�Hx"i�S��͟t8ZY��}�&���`+ �hXy�2���
߾@�Gkʆ@��:��t��h��=����U&~���#�SC} y��l�)�Bӈg�y�6�B☹�®l!��B�0��K��Y�^�4������G�v�qRFЊJ��R�֥u�B�rR�7&�ƞt�@|��ȥ�GV��X Z����B�'2�!f��:��a����U^EXH�M�+.H5@���(�4�UB%S���p��>����'	ZL���h|��V�a�4L_�k���O6�)����׽a���+�!�p�]͉,k�u�c���C�TLIc�P.�\edi2�Z�����i�,�yM�pRg�(&��X(�r�����'֥�zTy�s�7>y�<9�z�!����в��G-��)�����;���}2:=;��l��-�n�zXz�p�U�&���~�՗�=�秗�7��˺�}?ڹ���²\�r�������g�G~r����oϖ'�~`��6=?��S�ˇ<������9X��D��-#�~	^�]IZ+dRom�d`P�-�����kI�]P��p���k��H��X�p8��\��{���y��˞5ݻ������������K�Hy������������h�����W�^��ӗ6v���(絏�^;dV�w�:Z��
,�`.�t��-���e��l8옆N��$B���נ�
LAl-��횣P%�0�!��G|[�k��N���f
��k�
@��hL���]&=č&�m���o~��B3����Ѷqǒ�=��]��[L>�fg�Y����֟���1��3��n%���:��J�h����h���j�ei�o���y��\p�p�ŷ�@�#���RČ3QF����=y�SKy�����ye� `e ��۫����٩u�V�V���_��\����ի/�����?=��\�v�}���Վ���_��x��=�8�{���77�����������W��1�_a�j���3�o��yc���{�|�~���>�w䷆]!<�y���o��9v�t��?��������O�0ދ)�u�M�V�����ʞ���֤)�1k.Q\I�!�76��zg�]
�O��86s�\$=z��M�4����z��t�tJ��8��\z�>�D�JV>�4SE�U��9t�K�Nd}����1$E92�-��\luJGjN�!G�K�&��y�� V?M.C�I�Q��
'%VC�в�Ր�I��ڈ��5.��eg34.F��DL|;
Ұ��dR%�)�*_+WC�4d�ڹ�
�4�qm�� ���~
`��xg���K�D1&K6f��F�*�o)��Wv/�U���;��w�_������*�����u�����-\���!�^-��+�ڟ@�l�+z��U���*a�U�)t�04R᭭@ÚDj3��uRS��h
"+ µJ.�T�gh8���g�˕B!��!�82/�������j��P�A3�r)
���A$UFŔ�g����(�DȪ�����;��h?���!�]�}�y��Հ����m 4͡�8Nd5G
G:V�k+�"�'.�Ԟ0���;��M����Zᮮ@dk(\/���x��FK]�!����l6|��dk����� -5L�X���}��7���?���\"e���[�;LtF����1-�z�%/#�\�:\,)d��O�Pc+����p�`*G�������Ƅ��5;yE��.#|KQ�ǎ >�\DO+�s!�`E��JW�E���w��*�"��F��i&����~����`^�4ٚ�٬�*�k�Y%6���Q��P`�R��Άh\bM�J�hjkF���MLk+�\�B��p��b�R�/qEb����3�S�z�p5�˲�tq�!���rA�j�[HI��\I!�jl��sA�G.�k;h��NF:�*a( W�e�M�t�t��/<>���dkyK!c�,8�I���೥r�y�M.C�^�2��tl<v) �a���+�f��Ao^B�'��$8:���ߜ�m�:����&W[[k�L�U%�Cȋ��~*oF��&ESx:��W".d� S	����e&{�,53�Y��FSk�BF�(x�Y��a�a,Zw����՚;�^H�!�!8�"�X6��
��D�M-Con("WC�jfL�����X׭���^%\�d�Ts�hp4 WR1���\B���G>
=�J�M�����TR���+ a�$YC:&�������*2;hX���*���GUh��1'Q^S`�e�n�����2W��Y,�1=
e���L��_:�.u+ǉ�>/W�b�b�&�kn�e�`��A�VzU%[:3m��}Ml�A`�����񢄏2�a�Rm�����N`�ۋVm�֤������z)�iRCj��E���� N�qxCұn�Sf50�ǐ����BE��iX���\�hU�����-�� �akV[�y�N�pB���;*8o�����F�F.{4.F���G���j�)\�W�h��B�]�
/v�
4ӦS"}Qy٢�bg��"�6Ӻ��);Y��tՌ�I?q�D�I�C�5�(V�3�R�}rMy�M3�@�I���2��elk�TZ��������6��75�!��LT6os,cs,~�������*A���&v�rEsD�w*�g�N6�
�#h�g�ǋV������_lI�b �5 �������ly뷙�N-;N����,#;r:ʵ��Ƭ���UD��h�]H�׶|�,��I�5�vψZ������E�7���x>�yu�|8�ҭ�>��wv} �j߳8�n./v������0�� M@���ϙ���7�G;�����|��cw�ה}��U�]w_�kU�vd��Ƚ}�-w�7g���/�Gگ�~��gO7{������_�\w�R�R�KqkU?�34�R��9�BY����!�?�-���������M C�
:|��L�_��h����{&��ϫg�ֻ�~*�`�����؂^]_?|���O���퓏~�Kf�c�˫�����˧�\��<�QM+q~r�����������9�/9.�o�������՝k��UQ���3����]{Ƕ��[��8���Dm�&�>���LY���	�q
��Q��_C�I�>�Ъ-�����#�DckCfBj���\h��n:��BSp��ihW�}l�7��E�E��Ř��vY8MW?��� 4�nd�g������&b�io���K�(Ȝ�lM��*O�<;��4�C�kp�@�vC C���M��V��g�QHM���+�N���G6Aj	�CB��Gv��m3���:.�'�O��ο��9������o�>\~)��ɽ��ÇgO��7�~�����M{�X��v��ڇ�/N�>��?�p����rx}��/뛯��Ҹ�ŗ��9={�ݯ�|����o����W�~���Ͼ�a��������������;�������~y��!W!�~P�}h33쟦3/���wek)�f�6sQ�抖8�IAS�ɐB.#����ڹ�j�z�-���vջ1���S�����]*$����e�F���.1��V���ZުIMAD�M�P58.-�Ԑ���@_FC5g�B�P�Bs0J*�Ja:�^v��*7-�lv����3�>����k��#�Ȯ1���LA���%��y�Qc�H!�ِ�RD�f��G���p^��CDA�&�G�H��@.��S����8�3Ąjp�(h%*#��c�Ve,ٵދ�ϖ-W��ߪ�+Co�{�飖v{�:��p5ۊ�mo���riE8���v��J��%�@�pF ����C�2����V�p0<P�h���	��AS	�4�l�Q�}nF&+�b�qᴪ�pR�L"%Q j"�J�Qұ>�0)M�F��a�k�5�U�dg���H�u�1�DRH��U��ʀ���Gf�QC��T	��	��Y
�2��/1qiF�
_m4��R�ޱ�H�005:�!5�i����%��w��ȖEU��s*���lk���j���u�\��ҵ�lj#V���b���G�%���_%�DpH��&4H��[����0O��P�c} �=�]=�r�ljK��f�-\��G���Q�(:f1�QF
DM��@C!4�-�O��O]
��B,&YH!�p���HQ��7K��%��'�B�y�I�*�jP�[�B�<A����G3�,����=�%�fqdĔ�D������5��e�`Ȧ@��jWD�h��Pl��$�;I���c�J�%/���6�r�A�����C��,��6�th1��գi#�ND�l�x�-�4��C��eQ3-~:�B��	l��3)�	!U��Q�h�E!����B��
a`r�ѻ�m@x�pC!�p��AŖEH?Z�RI���z��
��|6Mv�c����BH	'�ل��#�s	d�OS�4����*a��eՐw�ov8މB0���NU��������+�
�B\�zH��Ud����Զ5�8z��@�j��ԐhlH|He�U ��~{\�4 ;���g��U���Dl^�k��7k�*��&r��U�캁�� �*Yp��!W8�
�r��զ ����r`^4-A�*���4K�S1�2"hK�l�����k�����ckzeX��!�om��0��2J����b��O��ֱ��Jri��\D�~
������."*�Z����^U� ��+��t5C�#0f�&]�F@F�����\�p-x54�Gf4�������dDKȆ\� hc�X�ن�(;�L'Z{8�	7m��9�A�W�"����/dj.c�\��8����D�Dq��"��p�K'a`��S�"�W_ټU>C�!�I������1��@���Yа,�i} �ĈcB�p=5"8��C�+G�p��!IWեZ^:��G�3=�U"D+\*�ā�t>&�TQ͈-ֵ���������.�!xC�v �4y���S/�E������@�#�4��d�Z�TQ dl7H�14�B���#����)�P:M )Ql̔�鄤/А�F���d�	�I3|�d)��H�Aع�!���G(u����
�:�-�p!f�jS,P�3.C�p��E�K�?���%��p̐4��\�o� 6/��M��� N���qQ_���|�UUӶ�h�����h��A�bj)3FbX=��b٘;�)n?#�%�>%�\�����w`7��'�փ��w�����5����������hwg���m��́��s��}�t��b������\��XO�W�/��w�����ǟ������+��Sfo������j�K�Iv=�ݨ"k-?��w������ol�<��ч˯}������V�3s^k�}u�Y[�VfI���\V�%�7lC�q�0G���0��9�od��g\�ط!�)ݽ�S,��:F�|���p�<���ӯ~{�ɇ�O��ٹ���<8z��Co<#���ˍw��y��=��+����;<}~r������?X�>�-_,��nˋ�r�֏o.y}׸4����D��7��hw2��0Gc���6��\�8�`�!_#4P�6�j��ϕl�CƘ�!LҌm$y��&�7_��^��| ��B�:��5h�I��d.G_�;�����XR\�qb�=[�P�q��A��"ӑ��*oR���b��#d�1y5v�
3�>�¹��Gs['PRFv^���\�n�\�tK:�xŎ`"��o����R#`I˲���2��S�YV~}Xh�ȿ�8�8��{����`�_0,�{ǰ�s}�yt�{��ǻ�'���V_z��/���+?��tst���>��������O)ݞ�;��?��8=�;����_y���N��}����/��o�b���w����޺w����s?عd��@��,�c�f��<�f�4��3+`�2f׬]B#,ӽ{�!�Jؖӣڙ�[�|��sݖ�E����ٸ��R	g��j�_�j�8�D�	n듓[��J7����-_�ݫ�|D�ML�9~�e�*�l��d����D�5!%EM"�js��K���3ʈ�F�@R�ea�������E�\���/��jD���.��
���+VO$6��ɅΆh�d�04�"	L�2����"��ٹ��76>����BP��ƀ�n�/P����){|} ����̱J�~�m�`���*e!�O���?�я��H
��-��s��*���u���=�m!^:��pd��m�Q�{��1U��j�4/����EP���b
i�h�"�!)�)S#�/�(5���6�y�c�������[Rd".��H
�6�.RT /�At�D�k�D��U���]��>p�칗,��JAA �8.Rv�b[���S(�)�)@M��j�M�[�l��fa�Y����ɶ��ʪ��ye�"=���%k��g�/�L���1�ά+��@u7eH�#���*��j��#v�
͑l:[�#U'RU�����R�^jQ}��CJmj� ��\��w̪2kj\zQ�b�L\=�V�"�tfaDU�Qc�X��W�jM�jV��ч�m=R�n�D��3�N�c�0��+�tD4Ф�1�hMl3��p�U�9�q�5ʡDH�������e^��[Cň"�\=R���~f�ꢽ�k    IDAT��JԻ��q���������,�@6
�n���pCF^!��D"VL/�)�[�l��a )(؂h-&����co:��S[�ʅ���h����.#�X��)��63�$�h�5.�X|��&YH^�@d����ՠ�ǩ=�,��lRZ�ڶZ�V�05Sh�p�W92/�&[=x�l}��)�ΎV,^^��8l��h\����v�mBxK'o8�hH?f����Qz�����7Wx�
�_C�t��M��G�xCCRfwD������A�^��(CR���@�"dW��}�R.�j�B���dSЗT��-B�m���e��RKP_j�1��������S4Գ5dpM�tԔ_$V&/��kh�q5����8�s��Щ"�٘;�Q6��(E4x�UE��Q�d�0d4Ld��X�\pG6&$W�U���C�{�4CЀe���@W��7MC��KZl���)�ZL.d���E!�1[��t�-�@�Z˲�4�h�Y��W�2,5Pxu�\��`B҇S�Paz���2Zv��e�������^
���Y�x+������)=��h�꣭��KA�N�B:�=�p4�^m��'RF����vHQ�9^|Mx`�ЦxR��ȋ��B�vd5��.v;����&�*���-^�ʀ����as���yiB��`�,�J$o�qM�b�5���%r-&���Un8�(vU�8k�Ȟ /�Db��p�bjy�'Q�a:��6� ��h[�["��	jjN�#H�5Y�Ԍ�,�`�t8�p���A�1G�좨U[��!��!U�׸D)���a6�J�|����2�M�w����d�,\}�єa��kh@�!�R�]��V��6R"QpQM�*�l��3"pL.�z�d'��� ��#O��K��'��ebkC� Q���YL}�"����
c8jz��k4eR�SN�]�('+D�4��P�!M!\�����[��d���n@ad���]��2©U��VO�����\^�r��"����rUI�p^���j�����y�x[�r}q���˨o���K,��)ۡ'f>���p��T'���|�-t�z�`o����S߉��G�˧(�{ܤ>����W_���O~�_��_,�>�qt}��W:��/D�L{Vzw��qs|��w^��������ىo�=�^����^��5�Mx�ۄ���|;[�UfYp��yWC���էK&=��n떨 C���gvus����x�˯>wG��_Avy~r}u�S|;nQ�/�Ĳ�sY������w4|;��K������G�ވ-���襗_�Ν́u���MK�|����|)�z}�y���
�0��,��~8�C��r��B.�:�P?CF��c��
�޵=�&L=C�E�k%�����7�1��kl�jq�l�~�����5�����.��3d���ʦ�*.[h�`v?��e-�h
` 0Rc�J�z�*h���k�d��_|kK����ޤJW���#�jyG��#T!<cB MV�6R%�kہ��b
�0�v�(3�q^./7��_��Kۻ��잞����'��~蝃�*zx���h��G�]����tMu�>x�����q��k׿������+/+���7�Gz��x��I����-v�}������K�o������7�x�<P�΋�x��������Z����������.�nX�w�2��ځ6�L���wm\R�2���� x]� Z1FQ�����o~��]��l]H�m���;�R+�Q��{�\������ow��Q��!��%�}�ds5�&��*4>�a�w��@?%�"0/#5=���)��*/M�\E��g����`�ԗ7)�X�j��_ϋLn�l�e�kJ��g^۳��,N
���@vC� U�B�#>e$�PT�T@�����s5���{ʳ8�}��5`
����x��J��d$�K�����(CM�� 2��C)�;�n�{�唰�1q��o�����R��5��N�i���?k�A8)�x�!�D򴣏dy@�T��q�*ʃL���
.g�թZ��o�b�����y��-�
IA��@�3��d�5����(;�(縇.B��>8=��R����OU	��ǷjF��L�Pc�����*5��P�Q6q�U��'?�C_��^��""���\��(�Pv�h8@Y8/�j$h�~�_��<�2)4�4�E!+G��6t軀�Z��<��ш�sa:��1ԣH�ӲʳJ�����-�Y��B��OD1h��3f��R{뭷|1��ۿy�&#�T����)�F��)F�f�xA�-�����J�"��:[�,�&Y�M��E9}��z���j�U��A��E�	� r	�ԇ;��Y�"zw�� ��S�áw@���ubz�R +/�a
������ v��?��?����������W뜂���3[I�?��?��?�X�� Y�l=[.����PC+��������E�c}�^:b5�d��!����}�T�bGA�K_�DGj[���N
��D􅋵��>C�DC��R�P 2
D�ڞ�ᔄi��03�M���,��eQ$�N.���,�3돦Mm�QK�\�Dt�x#W|S,~�M���ZkR�hM
Φ9��չ�-s1_��#��j�xS˛`���ASj!U�e�®4���!B��C���5��@}:b��GHM_1��z�Jb��a׬m���#u��=+�Liݥ��9����d줈s�y��̋ �^ P���&����fpec���l�d�1Ӈ$8�M��[%��U�~�(�քQ%�+C/$ÐNQ�@5�f�$^��Paj(0f��[�8�+�>�t0�Z����z $��4�dl��5R.���d�G`# M�p̔��F�z��_��F���!�@vj�@
�����苪`}Yo
8��q�#,��4��!5�C�ΰ�:�b�ʮLR2$)Ø�:5 ىO��ې�aY��U��>=�P�I�T��W��y�))pp�l:���!lI��:˘�62�!đwr�m:����%��ry���#��� h��3�o�.��X�DV��)a�4�e4�x:3T���n����i:�:R�a��Mܐ-�!���O��<�-0�ѡ����fX8;Co��;B
��4î��k�p�0';W�q��h�$5�� 	)�-d��,M�M�X}k(�F�т���do�7�t(1e�MxkB\F.�h���֊-#d��p�:�e3d7��D�ŧ ��6ALF�0�GPp6P`.:�4K
�
�o�&<Z}�ֈ�-
�<Q���De`ͼ��y�5/�L�\���!��F�\U	r��1K��ڀ83,>��J�� �4��]����.�B�Z��א+��e�����_48���D�a}5d,K��6�#rY
A�-$�^%c
s��$WS��FhWS�7�R�3JA�:���p����A���ۤK��^��ňn�n��O���{�_������w�;o�e8���ͧ�;��O�s��ٝ��/����So} h�uN�'�:�_88|�����/?����_=������]�r]�/OA���_>E�F6�fw���Ue��3���~����o��=�w����ӫ3ON�K����z�I��¶��|�S��lY��#[4�сX.�c�'[�]�Ocw�4�c���T��׺�@���� ���]�M�斉��Ʒ<��yx�w��޽�~D��������OO.��xt�ʓ�]?��w~us|��koX�{/xt���ol^�n���<�=�;�~�o}���ڍ��]߮���5Aŷjk���Y�?k8!�a��4$X,��AV��#��Zā'�MX�����["!�m�ݞ5�n��"��g�_,XH"��jKaȁ�Ѐ��,�J��5RZC�2�B�_�����uՃS�Bn���
яB�1�0�ZH��1��f@�jޮv��R���5�U��\#Xvv�ȋ�Ns��H����E-u��L.�(���E��I���cwy�2�./�?����������w_H{�+���_�\>;��8R7W������������_����|N���=�0���b�GJ�]����^�;�9��ݼ�����~������?��{�ׯ�������Ϯ�?w��i�^�음���;����nE����=_�ցa���,��֫[�Ɔ���%xY��)��&C�D��=C��K�ެ�\^�=���nպ�R#뇷6��'WM ��[}Z�rL��"!�*I������%�)̎%��Z�@3��^�n/Fd�>���H��+��0MB�Dy#�yb�z9Q�e�lHM��F�!���Z�W��/���$�A|F.}"z
ڬڄ��e�L�p=\,���0d�%�B ����h�Zu�A�*9����-*w�&C^�i6���p�ى���o��[��B�jveQ�DU��_�ʉg��8�e�0��7��=��.8�锅r�⅛[s��|�$!e?X�֟�-z��1��l�=7����;������3�"z�����0Le0֤�NN�����dwb���@L�L]h��N5�6�x�����LG����4�d{��� "��G "�ҥNAR8�K":�p=���+@�t)� gH�0!`NPm��V��8�r�+�M\`�Q�i�~�9|�)z�tX]p�t�EO^�gC���[o��DbB�J��04O�̥%U$����ҙ�c����!�ٟY�w�y���6�
�#;��҂̲4���ۿ�������O�S�:�*��L�� ~����-#�>r�υlSP������t�z�g����;uQ�	Z���{ό�r�d��[��\��1��ąh�
�0�x�Q�ȅ,��U�(8(�b��(���9b�V��mj8���C��u�+I"Op�qܽR�V����N�ë*v�a!A)d��lF�uҷ�6oSV��o"D�ٹf��X�!�@Yp��jX���|����B!8�m�l^e�����-����r�i�����bA�+[��
D+j�X��0��K���!8&�N!���HV[��-�P<q�\I�'��VU ׶Tv�������e)dZ�y᪆�zؼd���ņ3Z�ɋ�&���	��
1�.��c�༐!�k�ټ�H�>�#/\
�z5�A�U0����L���0$��p��њ���-U�hbS>&�Q.vs�J�'e}k��R`�Hx��P��B�U`+0��;��Ļ�&8��Ӥ���_z?���΢�Ԁ7�R�5�p^��@b����u(NՖ1;��-i�Ͱ~��p���U�a�!hp��;�)>�z�^Sp�2ZIȀh�he�+ b%�h�Ȣ�����)@���3�(`�!c4��3J�N=��p���WM��6�=r�l}C8�^x��U����(���\�y��:'���M�F�%%�vR.�z��lüە𖨒l{�k
i��J:Lk���My�
�6��8�j�C���l�Sa�͚�U���Y^C8�����U��QKP"�
\j�[ $"��5� ��չ�]O�]����Om���L���G.\_K���Sr6�v���֒e3L?�2�,|K���b3�L�B!q��A&�]I���w�;�i
I����ΨUU��ˈ��"���X5�5�B�h}��F6W�zH.=D�Ui�Wk���b��ފ��dLFR�hpR���!q��\����1
4�oA���_��'�7�6�\�'5o6�l5 c��!Kֻw�iV6�Q%h
e,���񅷞j.;0�~m��
���IqM%�p���M%�����ʕ��,�*��B�掶&�M=���������p��v�kQ_�������D��4�U�+;��K/5��P/�IE0��%,���0(��e�(`�r�q�V,5��GI���M�X:��Ɛ%r��S(�cZB��
I_Z�t������Dv�g/���g�^��I���QM7�<Gs)�9��<�q�;~_no�w�v��%�{;/�r���O�|����y��K����|[���Byv���A�}h���cj>ɹ�w���_=��onwv���<[>4z�s��D��@l�6�S�­�64.��3�l�@5P���/��.t켢�Z�r��-��	NF)�/��
��O?g�{������v}���ݍ�!�Ǿ�w�����������W�{>��������L̛���y���ǵ��]��{�	�r�w_W~�o=�ftw�ݾn�D.M�����7S���Ah�·AH�r��n�&�@-A=�m��!�ީJ,�'<����y�Ԛ5���;>�bj8Z�����-0A�aRzᆶ_:�!�����m"�Z�II<W��/)���m�����9٢&6������&�̛]Ή5dˢG`$�=5���9µ�qŏY
}ƶ$�(4���M�kY�x#G�s��}<����<�<�\�;����cߴ����������������볇��]\������}���/����^����݃�������)>�����c��uk^��=�峋��g�����W�v?�諓��gO.?���������>x�x��f�U�b�RI�:�m��.�雅f�zL W��B�-��0<>��u�X��8�v�C��FsR��Zj��u�ՍV4�
�h�sxB���^-	Wd��݃��N���$4!zd'�4r�Ѻd�5s�c���ք�b����@j\�b����z�z�'c���
��l.֥�xRU�����dl�5 ��e���̀Wp���%2d�pj��D{	dC��@F�2I1�*G��!�J��CVO��bF�PT��
�%�px�\1�3W�zC���h
�yK���N�װ��V�'v���<�x��7=��Ϡ0�jͲ�y(؟�4o#*��Lg�X[�\��M.�����R����~���q��")2}�>h.Z�deԣ�L�W1ֺ ˗v��h�b:΋@����0/D"|�-��g�0g�\8\��hl�z�l��e �Z�˶��!U�/\
T��l�R�d��+�sGUHȫY0��`����l䦏�͟(P�\zC����zR%��_qz58�d[�$2�f��V����+tO"�S��������'|�C"dL����#6�G�O-:����C&������W�����v ��a�*C�5���<W�G�r���Л��r͚�Q�,&�
��hwI����Y8|�������/����#� �W	C�-���ǩAS�t�*�fv�\eAhRz�F`GΛY=�hi�����lR��!�3ѡ��)��Y We��Y1!^�&em����("f��9�dM�-*��+������x���ԬQ���w���2V�홨�B"[^�KIj���ee8�@��
SC�KT���L'Q��oА!\���"h�l�X
�\@Q����j�R��1�"6��!��n�l�N!tH�R��&E��mW� ��H��>P�,R3�!G�S�-{C�B-M��C�tB�h����F�T�2��\t��^a8�7l�0���XH�3/^`:S$-0o.x������B���2Q�IA?y#�4f��8����������c�̆�'���l����	Ǉhe1�@H:���T5�j hM!o�F�v�Q�Eeұ�[䪂��tEU$qC}��
��d�$�c�E��
h�6!��3q8#��ZB�zY��l �U2,�׹ 6A�	D B\�*C�=�:�]�2��VF��e�0�D�X�B6�B��l�AAm�r%�4gj+wI�V�6~
q ^#ؔK���M�fG!�V���1����,�>� �3�������j���y�C3j(V�EӤ�4�`C�i�zLF6e�W�[�p��Rl:Șe�I��K$C���HR�	q������p���'Rd+ ��-�"5�J6|Rj��j�w�%ҹ<�d�L�,�q�gLR4uF.Ky"�l��W��C����mr1�Ӂ�ь��R�+,�>�vN�p��,\co�*�&�N�TL=Z�)�њ���c��D�ġ�H9N�-c�b�H8Ψf"z��JJMks��    IDAT�HP/�7<�c\6})Ȁq��s��Ϙ�:�P��ࡵV3��0��ɛ!6�k^s���b�'�OG�ڄ�rIټ�3����ObGЊ�d�KpͿLت�m�k��/�a�%
QUd����dp�@Qi�p����g�'���f.�-)&A ��=����@���ri�h�� q��@� ����O���z�T�p�N�q65F!\���\�q�5��"�u�6�.X�Y �"�~�#Lv6/![K-'��a� V[jqx�E����?.�c5��`��I��	_��_�Z^L����|��/�=>:ܽ��o�1��4�s7�́�狠��\��m���{�/�tϣ����'�=�����??�l�-���K�Sa�b�-�m�b?�Ih��M��d�c3}�o|�ų�=�z~�|���j�bw�i�L|��2�t���k5��`G�oX���]@,�\ݤr�������A�P"� �mE2�
���nf|������㋯��,�������󳽝���=/��^���<{�t��z��ͽ��+���������~ds)��c]�I�����XS�
�Q]���\d.�zw��ݴjF`�	ꕊ��ہ�H�Hbjk�[8a8�(�������s�P��fNl�3dh�E�!�d�-����a��t��R���m�k�pA���T|ǂd��4%�`=�Ϟ!Pf�o۹§�@���v`�z c�ܦ ��q�6,*&�2�٩VO)
�?r��F�O�І3�riSR����R���WM�]��٩w0���?v��y4'w\�<���Л�3��g�w�]�,7ٮ��|����^��ol|G���o������>�g��>�}��o���ſ�ԧB]n6W��O��藟�7#ܜޜ>|������b��/���gg�_~�ܺt���BBo������fݔ��ޜ�����$\�m��J�%M8����2�2�ܰu��ZJ�Z1�I���fY\=z���8N��k6��I�?��Z�ŗ��	��m�c+��Wr��;	!K��!Ͷ���fk�p!�E#(#��;M^E�Kd&%�����ӗы��	�U�>P���(5�RKQ:d}s.dɷ�$JQ\��sɦ��;��p�zCjz5Lͩ�DKa2
�p��|�-����@+�S�L%�3�$�R�]�߾$SD��F�;�g����q�Yز�5+������}o<+���!����	�5��4�c"�t|(�CO��f�/-]�K(C�T�B8�z4�%aKa�֨I$�tzotp�!U82�`=0;Y^W$͎#DƎ��q�:���
��Z+5D��E��K�W
������_�Z�'B� x4��bV-)�Z���Ŗ�P^�*�b�Iy�F<ې�[S6q �cdYx�r�JG�@������Ó��f e�\�v�=`��$BJ.
���qt��Zjh���_�%��ԣG�<���'d�>_�Zu��qO��k}6q�0��������P3Ae��UTū0�5�.\@d"\�VI��(�M���0U"#0>�)F����v�'��&K��#���MAICMx�,WGӐ��E�K!�0�&B
fgL�z:R���֡1�'A��H��t��R�z(}
��<�va���R �&}ӷ�HIʖ�Pߌ ���քl�+
3��ˢ;VC0�/ЌZd���PV��yu��<���0&��Q@%bU;A��`@$šυY1�M�Q�f�6��C"PHK�����&Ԉ ��H�B"�m���m�!-���֝�X�%g~�}˵�.�"���@�E$@�C��H_��f�-LW�����ʪ��"c���Vw�� ii���sܯG�{��d߉R[���0��NU�9e�6����q��8usZk��?MB�Η>�TGZ�__3B���h�X�8F��
5%($��ֿ�QE�H
�G
�@�N��(����E.4���Rz5�rʵ��Ս��G�,x�ʪ"~ݢq�q0��8F(e|S����m-�!n�-��<f���!�:�Iﵙ�MgF��~��0�I0q��U>N�5��Vք�i�k��+�(��t(��`��r)��DVhɿ߇�Y�S�&��.Jh����+�<:ҀB@NM&��BU��NJ8+���h8������F���0G�0���._9E���!4�I1���Ҭ�P/��XN��"�C��JޝD��,�͉_HSj�1�15ͺ�u�SJ
�6E3�k�wg��#�N�d;���aQY�����Y�Y���"SX����7�#G3�7�ᴱ�&R
P�AjZ�k��G3eS�f>\����Q�)��=�|#���O�ds���B���ҩ�;�N�D�h��;�()Ь
2$��÷b�o�Q���$�_�8h:��!hᛚ�Y�-��l��`� di|Hk�į���qq�hQ��9P�IL�4eS����'~Q�C��;j�B:��8Y��V���/��?B��,�9A��4���E�B��ZE��i�D�%;d�1!C�$U���PYm�\Lx
Y��b&�� �N�%��D�'�0�U�I�X~��U
��d�!Yd���qЌ	�k`��D>fd�1Rh��U�vɹo#�~������iY#n
4M'4m�I�I�D3���"�O*}Vl�ځsNb��~�Z�66q��l�fj�Ś�$�5IMRo�5u1�����,gZ�����i�i���b{bj��Ų�~^��'e��Bj2G"G���C��3`mq�h�K��������ў{�>�G�.o�q��;2�G�����T����l��u�������α7�W[�պ�����O^|��ҭ7(mm/?�/5�1s]H[����uj˶��\���v�֧�=��?�ųo��������;��"������!}~�����dkl�9�FQH`�сk������$�	��ө�^�=��)�O��|��M��Ѻu�,�榧�hZz�ɇG�/v��n/��_ｽ�z}������?��f�|�d��'�ny�{x|��΃���Z�,�kx�E�3+=�p���Z��1��V���L��K�,g9��K����}�����,>)#�\p��(�B��5�o���i��wƶP�"$crK��&�P�;�t�7��HqL���i���}B6j>5~Y�A�������!@L�@>S�&y�Ș%rS�6RjZŘ|�Qz%���ɖ5����� �p���pUL��q��e�o`�i�	�av���n2�
���ѯ�0��늾���i|	b�A{���G̞��?��"ݺ���Y�y�"��O�=��������N�|�zg�v�/~��>z��?����\L�O�v�ݺ�����g�_>|����N�ۋ�>�vg������Ƿ�~��7Ͼyy����'?x����Ź���ѣ�?�胏<՛u�֒]����_�:"�1�����^#>f�#i�]m�P��v�\-Wc���t�6���n�pj	.�!I��D�4�ƨ�ஶ
j��6����Aj%G"͎z����_�YLx�!+dXF�*����|��J�"���(��N��*���(45f�B�J�RW�-���=�"5����(;�C���9��*
p�6"GЏkud�L �dq(��
�I���1M1���˂Lr���h�1�᤼�ġ�ǩDj�)�-0BR�F��F�AH����;E��:����]r|9�4���'����b��#�3����B� �����E�4�E�	��׮���Y�!�%Q�~Dၳ9%R�I��4�Q(f�pꁅ�	Bp%$�!bZ�h6�Y�Z�h�K�45�C\=�qL`|���Cz��ޝ�.;���LR�-J��D�|�����Y�D0𑅀�-Α�~�wWK��<��sY�.RL&��EB�. �:�X�vYQ]A�VV�h��S4"���'� {�&=ÔRu��t�g5�
�A�bݭ|�|K�����Y:_��ӭD��F����{Kb��>��c���i�Q��(:���Y	����:!��RQ��|�,�ڨOb��D���0~Rp�ڨ�Y�~온%�l��40w���u\\�x�,j�)���?��m�v����/����[Y���z-Q�$��a�M5�SQ8|�%81(��$�@{+�>��B9���
��<�t��ٵ~JT�SV��j�̡�A�MS��E����Z�
�`�)�j�T1�@H�sF
D
0����CBd�M��n�(~[�Nb"#���>g�gJ���h Gz>+�C d*�l=�!��C��ϦU�n:ӏ��&�O9v�բ��5��,�������>~SS�D>��Qu�\!Ӣ|x~����.��р�q�����8D9QS#8�8�^>v;�, D@��D��o� 81��5pR� i�BZNuˍ��,a3]�"�iP#�8$q�ͬi2�iL��ʂ�|#fY��s�p��ؐ�\�DJG��_�eNB]�m�,��v�tUڍNc)8���rМޭ��B��!%DĀ�C�))���h�!�V"E'�Q���(�Ӕ�)����BZ&+Q��\N,+�)'���B*��Ǵ�R6�kCȯVUL���cD�á��s&�/�S�r4鵔-��X��#���7 c�g��$hC�Zc���K��!Kt�6U�,���٢l� 7�L�>M�Rw�z>p�'"������ӹ�/��6QA�� ���#�2��m�'h�a������"0�0�[��&������V�~"�;��P��V1=�-� �B" P��5����}p���q��/e�}S(ٺ�+Z��D�ik��3�5I8C�Q����]��RW�F�OMa����r�89pV{��u�,+Z��,w��1��� ou�V����>r+>-A�1�H��)N'���O�c�� %��B0��Ʌ����Z5m���.��(� ��6J��X� ����B����I3�p�	�����9��g�=/�ILPo�
*�
Iሎ�P��q�UHY�4�Mn�P��qL��G$��8D�J��i�w�qf��@Ͱh~��Z[��P�J��~��B�ʇ���N�A����6*�)˧��G���gZ�3b�q���#[�hY��aE!�r-���M\�|�開���o�\I�_����o�\�g{��0�z�y{��ףּ�h�r;�~����5��9��9>,ѻ�n��/�<��F�'���۳ߝ��o{��K�;׻��,�6���Ҳ�:�k{�#�Wˆ�pow���GGϾ~�`����W۞�:�9��e9�����Bz��κ]
�p��
ަ��30�~􎢟���?�����|���n>n�Htʡ�r���`?}s�|�7-Y�n6.?¿|�����/����������n//���_��G��<����ã����s(���ԏO<~���ۿ�|���m�˛�.�O/��}׷�7����\���Rc��n��M��ivI�?�J�h>f4�+�P��ѵH��O��_����l�l=��q��sBւ�G��R���*�³ӿi�>���dt���5SQ~%�'q��:w�L���T
�[��l��r��I�(��i��ƙ�3�r2�At�T��M[�f� @Y
�ZD�Fj��T����p��
�&�%ֶ�Yk�NE���!7E��5��sM�"kQY��CĽ��'���[7W�����s�}{�|Es!uA9|�h�����{7g/���r����|�urqyLz����o���?8|��:����K�_�8?�xsz���o~���o�/��v����������ã/����G�Ͽ}��ͫ탽�ۛ�'��Z�ٷ�������_v�t����]zC���Y���7���U�nɖ6ߢ���@C�-b�n֯w�m��ûҺuis�w���(��U������ni
��[Lo���ȓO���۴+Y%�Ҋ����:Z�d�Y�+Į�r18�Zj�㴰��� ��m�u�)T�8RJ�I9K�#j�5�bw*����\b4)��+d��2dR�d��6��Y�,)����rB����RlE|������+�)�?̦8i
��o:x��4�o9����9��Lc�RV�� �
Mڞ�J����`����1~I���Ox��'|�F��t���R��P����ac�4�@ ��A�{�8��� s�U�3D��'����:��m�nZ�SY�%��4��(Q�5S9#qְ"��!=>5C�t�pS�#
�!G-��,�c��	�bT��/������jy3`��Iq�j�Y�r�PE�. ��Vi�p{�R��yIS�����ylj^J㨋&� �c��6B*�?��?��QƲ\�=��,ꪭ��c@�@dQ�gNKh7�BܓQ���,L�)4u�5lipq��M�4���U�����������+_f|!�P�|�����dR�ԪsULkA!(�H�oQC�_��,g��c�9�c�.�	4c4�o�:�\(X�-էZp�s	n�@:hz���\X����cg��mx/ۊʚ�-A
�E��#�*�I��팍J�)a �{��NJ��e��'�NZo���!^?D˗خ:<V�:
����]��^M��M�N'�r �D��B�m�qX�R�I��*��9�cpp�'�Z�rk���M'��P
<>234c����Y	~S��:4E�(2��T~�r�4�U~�D#@l��X4��R>)| 2��h�c��u45���pS�(�HY�i2 '�B���SXxk37[2mQ�U�ɕ� Kd|)���>YL��F���d�É�I8��!�z	B��Y#���@��*��l�2��z�o�ŏ-��}����!Z?�-��Eb5��ۦ��q�7�>N��GΉ�"�X8_:�Q!N����N�ٟr��zg�G��BL"��C-�cL��8�lv-ͤ �r�N���+�fQNSM{:l�C�g-�>ThL��ӔkR��ۋ:����c«HStվ;�W��7�T�M!&�T�>Yc�E;��s�ٜ�`�k�C_-:��(W��E� ؔ��N�@H��y�jO�2��5]�ᰪ�M�z� S��M7�c�[�7M
�r�/%e~��U��B�ԈXHm�ȩ���%�)�a�*�/���"��R��1�F�n���z�*����|82���J�}k�#�e�F���h,~+�
�Qu��WQ�uoK9�P%BH���Tm��i���ؘ�Q��8���yeI6�WK!�Qp"��V�hZ�����9Ʊv�3m�I!Y�B�LcsZ3}+T')�[r`�YuqںYXV���j�P�u�SnSL�a����h񓊟x�J�Ƥ�`N~��g)��K��tJ)4�ړ�ֶ�3"B��"#�/��X!>�TV)��D*T4�/� Q�	iZ�D֏-.&M[�;m(���"�S!:� H�=e?dՆ�Z>�6 tL��b��-�T�U���YQ�$�O���_�I��s��g�;��Xi�T�Md�1h�5����t�������g�=��?o5��51�W��Lo����N"�?�oGXvr{�{�����x�;�7�'��3xs�|�w��e_��������}>���v�Y̭����O�{��mD�����b���)��^�������7�п���W?~���l��>�c��ۭ}{']�m��6�T]�*�l2Ǐ�p����'���q��f͟���>I��'�_w����w�u&1����B�y�N�f��?���͛��_�ܺ�:���g�=|�hw�����CI��.g���
;���履<8<�x���o��Psy��`�u-�˷�[B� # !Vj���h�a����{�f�m?q(q88��ߜ.���-B�&��-M栍?
�n�����w�Yx��[&|�2|N ˯��M� D�t�6�A�:�v/�����X r�9���4����`��y5�'X?��3vB����F���9Y�M[N���>N-qR8V��Գ��$r�l"��h*w�o��o�\��!�/[f��?U_m���}��qp�������������?�������]7�w/��L�f��p���^^>��N��W����?�=�������g����g����v�������c��1��~����G�O���y�����g��w�ؽ>�~��?:���zsz��ͩ7w����].?V��Z\�\p6Ҟ#�k�LN��'B�|YpӬ$�    IDAT6�"�3�D ��E�ȍ	q�t?����|�`z����yH��(~�ĵ����P��P���mI~D�Z��Y�J��β+)�5:������.�˾�/�N ?�Y�|#+�t�$��H�7jLV���@MJđՔm*���p�d����RC�I���W�Ԣ�@��o�7���U��AP1$'D����-^"�F�U7����5�tZ�_���a�S��f�-�Y3h�(�w6w�l���J���I�g��n��M�h�N���h���R<�L�	oH��-4��Ԍ�ZŇ`����B�obL�NT��>�%E\
�6�$7_"�ڕX:^��SP�_b�p���f��jO�M�a�8u�;0)�!ۢT��:B�rj�S ��u�!��1�bR@W+�6_n�*J1D���zH��(�5��[���eIl]�Y8���b�+Q�Y�z���H'��<(BV��u�ub�_��]d1=X2j���7�7����JGmH��|��;���V�Ҫ��*�-D:��6��W���8�B�@�<��Ν�B�H\vd}���` ��~������a�ʡ!#$^uYm��H���X�d9����B��b�f,���kAЀf�|�MVT�+��Sj���� �s_�{	8���J���U��*��(Yh��� ��h�6m��V�@����N>��s?��Ԥp�A�v.�a+r��L��S.S��ez�;�*:!���t�D ��|mUH�]:[M%�(E�5j���A^�wg�L#�$§?��.!u�{8�dG|�")�5es$&�>#q���O���B�)G�N(�g1�Z�/N:B�c���c��Ti������v�G��JS0���gdM��M�h
�SR�%Rnih1�tYBF>NE����zҲBtl�'e)p�Ֆ� >f��r�&��~r ��oCRfs0���Bj�cdE�v�CR:\��@ӡ5�R
q�F��L��(��	M�ZE�:4ůb
���V�S絊<
ʵ��Mg�6G��8�4�JT����r�GM�.tc���i�uŁ�D����E!��k��F�i��#QV��/$]"ܨ��l_�IA��62��pNCn]�J�a*��p��QKMSS�n:6�98�Q�\���,%BRB��IG:�~ ��\
���L��O`���^צ��F��Uk,!����a)��wW�bqT4�ZH�n�*�Bs�X��A�S0:�i�ь�5�,�4Z�i�њB8�l>Gb>k� w���d��B��N���H'fY�)Ag>��8���(
1nf���B��3�҅j�Ĵ�L���u�i�ȭ"��#	4�M��B�4�Z��֔Æġ`��b�3��U"Ѧ�DL����P�(2���T��q�����pL�Ԫl*�N��8��?5|���R���9�ͩ��w��U�]B��Vm��j2�@�sO�1L��7&;�:�39!�N)@Ӛ�+"@�5*��im�#�hjE�~-��$e�����:[�k���5r tf��p��Y��8G3,)
���o�21�0�K��#g5P�����5L3���_c��V��`u�"�w�����Os��!�cʧ\:���L=Ԙ���!mZuk,�,�X�Z���a��)N�T��Rp��9Bu�(ޟ-�
����D��%n�B�mWs��gy%^��g�=?_~ҧ`� >G197�w�5��m��>֟��A7W[�{�.G���y�+��VA��[����#�ޡwg�]�c�W{;�׏O|p���������!�w6-?\�Dܻ+�����n�sk��	�ukǽ�����w������G�>�g�n��8�v���'Bv�m�+��i��s�h3�,�7��
�v��t��שׂb�|��D!
ݡR�D�nG�L7�p��(�t7�jp�����n.N� ��N���+�u��}�l./�oyZ{�w��	tK����7�>:�?z�ec�O߾��������#��zs�)��ͥǣvԛfX_Ʋ��#w_� �b�����93©qQ�7!�+:���m����TqU��jM�bj�%N�@������<"萅�Sؔũ1N�Mg����!u�����VT=f"l�G�0��Bݬ�� qV���A��d1#��E� kj�ڄ��Y��C6��|�#�Dx~�w�Q�V�X-6�鐉��|UF$���'����B('�46�\\�A�z�������g����v��e���վ��y{�ֻ$.�O�ū�������wn>z����დ?�胟���w��o^~��WG~��v�e�����/���}���u��z����g_����]�~=�ų�Ͼ���G���Ͽ������/�����7���������X��*Y�2;cڗ6H���6!&0ǘDN��q�#n�r<stq�-]c����ǕP���F���i�\<=���㏉x��#�K����ʘ������-�J"�>��J��	1���:�q-]Ǣ˱\�6%L���Gz��V:��4��NW��A�`E�)$����WzH�g�ǉ\h�
4Z�Lm=���4�*�|n
��J6�5�ۙR�o�v�$��ۺhY�)#l��K�V�V����!���4���	D08r�
�VJ��e�RL9���-�%�ز(pl�sn�|YN�G?��S��O?�=�s��g`zา���u�$RS�iC'e6\�o509����b�v
B�	Ĵ� �X�H�8ZjE��^�-]�I@�>G�q+J��?�(�(LB֊$�Bؐ�,��p���^Q|j��!2?���"n�7p��Y)+J�����Dӑ�S���t��|L�r)�Fɉ���k�ڦ��w1Ԙ�����^)L�׻ޑ]m�?���"��/���|r�*!�����6Iߪz�	�n��W�u�:
�h�H��Y���ZG{|=�Ґ�,��3��B0��z]��@��v@;/���	�V�>����-��S�x.�q>f�&[!)-DW���=�ki�'Ň�p*Zn%������9��6E�c���N��0Y��5�$�`��@S�6�x��X[#�@�m܁s��!b8�������ee	�������FYME5)K�J�Yi� {�H��t�"C{�"Ho�JAhLq�)WQ(P�!
��
�MZ�=A60�d�G�^iS4%�A@3�R���eh���n"�l�մ�'���ۤ8�!|�Uh,GV�@ӜJԉ\�*G�i\n|Q�8�z��n*�]���� ���9F����C�B0��91����n�;�)����z`����q�b��8uR(Yg�[ȴ�K�cp�5/�0�ƈ-�&�^�u^.�N�F���)������T���)����mS�r�x|>�P/�Dh�����!�
�rHa��r����j��N4��L�Wxٱ�+Eq6�A3�%�JCp����|:�eS�J(�s�gө"�6�%��ߒ9�cȒ^.k k���N�8�BhQ�� ���~CV�~ZK-&�\j8UOaU��J�%V�M�O'�I��m�S�����D0L�XH�C ���� ����B��e���o*T����hK�:�q����VTsM�RS
� ���s6M���Bk��Mk;f�U]h�(?Q4�[�h>�>&Z��16��S=�ɵ��X�^ 2N����|��NS�"��t>p�YS�㮊���Q�lk��M�Z����qJ�PŐY�*��	�L�|N�6*�H�SV:��Вg	jB#.T:��")�t�S65�eӪ'�2�4�iVA~���D�`AHI�����H:83�!�B'޴'
l�q ���r�e���	��aD8@"�����B�S�����R�eTT?�S� �dפ�/��d���p�J�98�����)rȏ/d����+�V4YӘE�$��G ���hL���L>��,��"/׀4�M�MS��(p�##|R:��`�MiS�L!¨�h�t����s�7�3K�~�B��nڲ�6�P������:�hJ�zR�h�YY𘜩���y�b*W��BD��~jnÁIQ�(-7&�0�PURcs� �q09�I����j�U>�T��ٜ���������9�A��鲖s��P�w:�sa���!�S�層Ŝ�//��������wg��\,������>���;�n����l����7g�n�����������4A����y��n���tU�?���p�\]� Ǜ��s��ڏ �Z�v�M���a�֦�dK^��/Չ�KY���(�^��!���N*�]��;�N�Lq���aY>��p�cу���}��U:V�~����_<|������n��^/��}��U�n}�پ�������֡��}�����3_ѯ<t^>�wy��?�I�~��A���A��ɶ쭮���Y7i9-C" �:�B,�3�Z$�	�J�a�J̶��
唞&D�B��;x��D ��_�E�_�d�O�����I������V+y3��M�M��)֘B}B��C��s>ghRLC&�t��N��s%V1�z-���O����J�D�@v��Q�lLb�|���/��F�(�;�ȆOgz��X�?N;�4�Z�,w}y�W�{�ʕ��w���/i�y{u�b��H|�V9���.N_���~�l�ʕ�l��f�����������ß���x|������_}wa���ƛW�o/���<y����W2o�t_��Ɵ������o^��Z���Oo~����ow�v�<��|���}n��O?<y���k�<b�f9�@v�q�P��b�Υ̋T�.D-���̎q��hj�@\���Q��]!�.KwaTH�������t����@S��?�x�O>v�%AK��t�?w~��
'�w��K��Q��}gU� ,G�8-L����b�)ck��ԧ�ʹ=m��.�V�5(�	ʪaU�lISNBg��n���LW�sP�I%ˏC��&K�����ďO�r��p�1�.G0������\�F�q�Hm��qd���ػ�`MED�U(]8Κ�����i)qR�oֱh�(;uk�u��Sߧ-Á
9�}�!��͖LA�gR �EVԋD����բ������j�p�m/&'��)�'N����i�)�q�F�M��-��o+�Np�b18B8�C�ӆ�w��wy��8��l�t"v��7��͙)�r��W�&��bV�OԤ(�p4N��|�vE�b��N*mH�5⣦y���:e�4��L���V�STp�8�����=)wyu����'e
���_��%�T����OV	2Kt~:u��?����L��j�h�U)�";u���y;	��Gй�Mg>B"��u�U��EcΊ��^t�^8R�K!B��(���&$�ϗbv\�5Lm�L�(Z�N'Y?*�	qK�ۄ
q,ܡҧ���g�g,M]_8�Ҫ4���5v�Y�B��l;A.�&�m�8���I'��1b��"}�"ܪ;�����GVKzS�Ȧَ����I�2���J�3�4A��!D���![�=���c���5����
� D����I�c�o��A6�d1���Y{��R�X������	B������*�*$J��:i�@!˙Ңhq�F�h�hՒΉ�\�S{,��Ё�%N3!�	rT	L��'B[j���Tw�VLj2�dj)�!洮S
������(��P|d��g�:��8|#��)(�����٦���L��i�T��c"(�(<N����ƴ��j���dq,� ��U��^G���u��WťF��t�E�4r%���ǐ���ϱK@N�pdщS���1��VK�)���׉��E�t�BmQ��-J�J���Q�iL�B~+%��N�	�e��a
1[�t4R2�ZYSv�,_eA�-A������Q�O�tH)�!
�">f��Oy�g�����%J�B�>��B�Ǉס,�|N�~�B�țj���ߨt�!e�F�h��#,Z�YHk,*R(���ʇ�bo{�
g�)_WJ�l �b�,�(\
��q������#�t>�W��]��)��Z)p~�:a1I�D� s ���,7��rQN��>���6���FkIy:��OAz��@���\xˉ�RlE{;><%e�0-�
���G��催�E�%Ƭ7�Q��`�h?SNm����]�Y5g�rL��6�笘uũt�#����'��H
^�N���+D� (ѴlA���,�8����t�t�_�/��p:�4�F�AZHL���TG��7��s��`Q-P4�R���o��x!����l
�����7�!Y:S��Z�P��>�ȱ:|Y��W2=D�b���R�ɚrʊ�W�
;�*�o�ߪM�紖M;-M94Y#ML��U�!5~��V(��D�2J���X�tX�O�����É#j�;:@��U��K/ԡ�����P�n�V4�,�ԨS4o�\�^���bb�;新����٭�뫝ݝ��k�\{[��́��ys������w��}sw�}��#G�v{�؁غ��U���-�����㫃ݧ�P;��y�������������Ιw]_�4\���!�����Y���*{�jn�5�]m]�_��\�����{g~w�����닳ý��7�n�k]��Y����l��b��t~S�@��@W*��@s�͚��F��p��pR���]�#$����~��g�=����ߘ����g��%w~��z��'�<{}�������w{�}�ws�͗��x���GۻG���wO�w֯�*,W��(_��h^������׉P���o����@�B�%��O��Ŷo#T�5�B�!V��!0'H�)[3����D�_{ᬬ���E��TM
^�dS+��t*��!�\��L�/dJ7]t�	�	$��O��?BH��d;�u�����؜rG|B����68�h��k�1m�V�t��Y:�o&~�GfE���ɯ+���J\���Ij.��r����7�O߼�~	Ħ\���Y�r����''�[ܫ���wA��݅�����o_z����Ǐ�9;��g���z�ݛ�_���\�&����������G��/y��{x�ԭO�S�v�_��=�����_��ԧ�������o�]�;!�
-���qw@�+�Z�K�}pM�wB�F6y�ǥOz��Ő���L�����R�rY���ޱ&���(�'�`����g��kq���ufk\^]�%Ct�v����e�������47�X���`�z�"BM	�A
͔��z��*H�DsJi+)�­A����:�Fq|S�Q't�&����A[��\���_H��A(
�Rm4D%�M�ű�B�4Y-GVS4�x�3�����e�j#P��5Ɓ����B���T�A�Et�yJ� �6F��a��3��Ջ:��{���y���EY��C�\�%PNܙ�@��e9L���C9L�����J�텦�M)�K�tӤDg!�.�t���mS�H��A��kG�4�7�_9+��B�@��j�^��(J�O�,x|��j�/��KA�7���l[Q���Q�����û�A��[�ui��!���tٶ��8t��1�u��/?s*�f� ג5�ȱ?�VZbQ��Бe�Oňh����I��P��������H�.9�l��<�NǺm��"ؒ9vC!SE�r��v"=��d�
i�Tz
�p��6Y�V�W� �Z����v�[U8���M��Tl�jͰ@]���7���k�.�JCbj�T���~ ���ݞ;v%��8��8Bj-��<֌��.n��Ӥ�髧��4��� J��&[��Z�,��V���)�$����)��_�)��m)k^?��R
����-~��!�lJ�pnRY�8u%E�|��\�zf�,�HG	H8j"8��'�`$�S ��E# 9F�YÔfS�ځ5�L�gj��9�ijٺ*e)���S"�h������p��S�8�p�D�3,���Y�fWr�aNo� ��X�֫���"�|;7$�NV��E��ES�֔�W(�ĝ��J�q��OP�e�.��_/�)1�r�Y�?KA!��aI!'hZ"�lJP�᷁�YC�s��0�55�6&�#�^�A��*7pȜ��)(gh��B�I���E'�q�<    IDAT+GTnQ|�\�F`���#%��ZY,��T3�͏�!�	�Pg樭�CG!YRX>�ܩ���8��1�D�H����U��huɡ�TS6�,Q"��K��5�)����r�����E#�BY,B�u	�UJ�!�,�k"4F����%Z�iMw�u2~��C�|�BkƢ3�S��,���X +�B=��*:�))���)�!���rk,�du_�(��6���V>)��c�dM�V����1V���sd�� �\�V�������T�-���s!-��2\�L~>�Bi:�EӉ�&X��Yng�)>/�c��lӮ���K�%�J_6_H,eW�D�B�(���Y�*�����7�"�B5�W���B�J���S(M���f�R�0~̤Xd
iN"��+ڦ�R���o��T:��c��'��q�x�Y�pF�_!N#f�Q�T��ku:Qؠ�A�7�;��*��O�i��N'������@�Hq(��9�׼�7*D�f�r�ê[Hj�6{��Jǜ~ȶ	�I	YB/R�8�e�K����՚!UHԠ����N�5�I�_Ř	�GT�8c	�����]W��O?O!���d�B���]=�)TE��O�Z���F:�j�&!��&�\�8|�h)�\m8嚆#HaKgsD��9���͔�x�3fѶzr9��E�)�a�xR�?�l�e�T��ɻҗ�[O=���3����O��w�io}��펏I���L&��SIO*�]?8�9��{�p���Ǉ�f���7�4�Wn���p�x`������|��lݶ_j1nY�����������:ON�^޾qi����?�/?;[�a-�o���ڟ@x_����B��a�R!̦|�� �gp�ۉP?_��i*����%��?{��!Yn�>�V��o�����j��r��ͫ=�b���������ڞ.�h��b�����' o�:s�`�=�s1�����z/��%�*��<���'ÜB��ꙣ��M�n��!��4�a/�(�f�5�.q��A�Y��g1���R�V1Շ��NY���pYb��ojT���s&:�B�t�S��4-��Ɵ��r����� ����L�$�t��1>N4H�)W�l��N��Mp4әPx�	�	��g7E em�!������t�Snj�iOL�;�#g� ���$�t������,}+ k��2���^yt~�֫�=�m����������ܫغz���o�������띓��������COCU�;x{y�M�����J�7߾����n=��㓇G��}q����у�g�\߾z�i�������{��u]��㴢��i�2�1��g��s8\d��� w�9��W%>���q�.�՘����_��m�n\���3�>��#��hs��?���.��k����r�AQ�hZjw�ӮC�6�%�
8p�"1[@ �V�2p��CXE�R��-��n̢l�a
�ĳ�7�H�n"+Q?ͣ�ƔNY�t�Pڀ�e�p��ǡ94Y!l���t�>������g-�|�n�-��X\ϳ�ɊoQ�S�~)��)]Wi��P
)!C(q<D@B��h���I�tX�6X#$f~8���Y���
q|C�l���~�Oܹ�lq2x���1���o$Z�;�No�!��$��#H��Q4�T
R���g��h{�j8X������OY{|�@��r�^H�h9�p��H"��P�f�%��v)� ��p��������װ�D��%hg������?��L��D�>�׆;@D��+�:1�յ�)Y�
x�� �jL.�Zs���*� �iK��5�6�E�[�g�}�cX��6�����o�j9+�oF�G�G)�����i����[벱����7@?V��%cұ@�h�zփ�V4��1p�p���q%G �XB��Q���;Z�r�օ�E�yb�q�s,�B����훕�p=)m	���i=G�C�K'iʗ^�l�A��5��iGܔ�oE��%��eڥJX���4�slQ�#�H�q��@����ՓSc�9���O&��g��k��o�@pZE�Ii-�,�@&+���UlR8BSG������W��T�D:E�h��5�l�����r�S�����-���S��Ϣ�Q�hʩ[N,�u h��u?[Q���:�"Q�����iOb��j�T
Zh:������bw�1��z`U	�f����1��3�������&آ*η��t��D�i�O�*ț��K�
��T�T�4d�)ݴ#e:�HS�(;SM�;
���[-����ƒ��&ҩUQdN"�"����@��f�B ��!E'+4����>m��N�E%���@�h�
F�r@2\�}�N;S��� 8�E6�#G�a*D��8�U�T�5&kJȅ/�����_>��q�C� t�$*�r��.�ܥ��1��TV��dEi�a��8���4�#R���%�q�Yd�e5e��/���dS��J�{5�M%b�%XJ�;;�I�CA�1������B�@)��YQvt���<����)��P=�X3���P;`�#+�rD���4�+�Hu�Z�)�S����E��OjU�{��!Sn96B�ΓKdS��8�Bb&;��a/Hd�r�(���1Z�G4U��Yxgc�@|��S�f|N�l�ZK������5�Hܷ1B�E�R�E5И�p�8���Q��:<Y�3D�W���\H��P>�`�o�����B̱iR��xQxW]�5���/�W�㵠��r��� �kj���U��a������?B�(PQeZ��9F̦�5W�Up���)r=d#���������0!�o:��	��mc�B�J��

B<���h����S	�����eQ�X~S[?��e��F���)!��$U?q�.�5 ��t�h-��ɰ�.��J���@�ղ(�p�8�N�I!�����t�m��P:�|H���s6���J�bE�Z{@H���IqµM�4$���׭N��qB0(��8�C|r�?Ҷ}��V�>�'�҅g��Y�6�֍������{8����|Z�����<�L�����ܱ?[>���|�އ���x��ԣ��[W;{G�t�ko&ҙ��3痽W�[?�,K��������Tw�v��p�x��==� ��c����\{�j)�ECf�i�:l���[���i��w��X�2t�'��?��8�&��NM�A����Eh�2ML7�SrW�/�[���7k��G�������[?�ѓ������Wϭ���n]��Z�oo.�AMO+�޼�x�ݫ�^�y����7_}�����H��qB'O�����X�	j��*��2�S��W�����r1Y!V�Be�� 9�X����>�=�N�B;0�!��ID6����ߡ�����5���`~�z�D��ɐ��~b�'�m��&Դ�|��ĉ0Y���,�����d˝,Ӷq��D˖8)��c��?���$ܧ�R{��Pv3W
�mIA�����۰.{;//N]�����<n����.���{��k���ի������N�^�uO��������^������O�/����}~���o_�8�p��o������������o��͗ϟ���۽�gߜ~���?�����E<��ë�3�`�^��~�������,�W.-����yW-��KA+Epe�����E��,v�]]]� ��~�����.��=��ۭn�����n��P�H��=���?e��O�y2᦭+,E*z�l�qXrJ6��1[*)�ٰG�G���*9�����<�QY�5�(Cꍥ G`�b>N��j�%�G N$�T��0�Sh�%��\4�p�����]��������j#����g�
%["nQUL�>�"2���ok�B�S�B�i����Պ���hvD��Hوዲ���8@�	�Cս$<L�ۿ�[�5E=F��?�sο�ۿy8G��:����m��/U<��h���E�(�N�N_9Q�TQæ8��ey-��Ƒi�>�l����!�� �ԉ�bU��ĳuRi�<yC���}���˿6��#O��]� F�<��M����8:�r���_/�woAF�u�z� Z�/ֽ�	�4�vX8.Gu+���B�O'eV҅*J�������Ai��M\��k�6�j����o�Xxͳ.ʲ���w��N���������=��?���*Z�B��9_	�)f�s�ʵ�@�a]No�Bi���HJ��ܯx��_��������6��]_4�C\'�X�Ta)/=ݏ6�e�cE��%JG� NV���B9l�R�acB�v(-J��D��u�wȀVd��vB�%��~_,�����;�F;+m�U�RK�<�!�I 6@ɿ�
pd4 ��GST9&���)�BU���~"��	l��|މ�R�%�i�˪�j�K�u)>�}ï�����thZ?��(�o�A0U��!��SJ���[ˈ$���IU���Po�qFv�L��F_h��������Y��u(EH'@�i�Y����E.�ݜ�ߢ���rH4�Q�8�v�fjS6Pc8�E��d>k ��笑��6����U6�S�*A!�(G��r�Ț�����KSn'y"�@Yd:�j��f>&�?����LR�q�� A��!['�Ҳ��(46i|Q6<���%t��ͱn��n�#%$��,)`��Bô�y���Ѭ+`��B��PS�4�q ,���cή��a;4�Z�Z�.�I�c�C���m��4k MVc��l�b8�M�r�q��-%_�0�����r��u�8��	V�nM���O$)m�)�h��ٕ���D6YW;9� �J6�Z�7E��#�);��Aʅ�l�gL���q�Ԓ��G�l^��h��+ڊkIhzC��05"��o���Č�&�n�M1�!'��Sf!x�M�����S�*�d����*$��&ܴ+@Y�����N�tR���W�nk�2|�.��&q��R��S3Q����Y�Պ�YK��M_JC�!4�#�m�ymD0�Tn�����7͆�Β��	ҋ�S��tSVE|`��Ӻ�д,H�T��j!�l�%f���lr��p�7�Ժ$�JSk�ZT>�)��ȊR���6m��M�@��	��8��Sϐ�љ��ֶ(ZLV��Tt�R(RR!6}!�h_�L�@�7~U*JP���ǯ"M��ҥ�4D�}3��F��1��Fb�G�>Y8	Z�\~�_�@�p��v����Ci�� >����{��!|�� eA��@��æ0�M��as/)�%�'U���P(rSQ�B����UI������	R�Ӕ��З�����#��H����ʭ��]����|��^ڽm�j��9�u�f9�~�eo.��q�������7wn]���w��֍�ˋ�ý���#� ݰ8<�DN�����}Z��<gU�(�r5Lxy��RZ��������N��O�zyv�<=XN�Ea��5��}�j�0�t�d�"ȑ�u��;�����~���9��h|R��7�D������������/:�;�7�\_�������w_�y�|k���ޓEG��YN���]�O����;�y/�N}R��թEy��?��몖�6�}0��攛�8P7��M-?������'k��tXC(gB��hir98񳘖flr&���4���~���N6�࣓T)E'4�`x�;Vi�V���N�q$
�!�Y��N�|j�0��`)��Q�5`:�9R,=|htji�Rdq8;mo��/�����ħ��X�&8�����d��k`S�ܩ��4��"���.n�>z���ޡ����������X��`oM�<:�H�%u�7����[}�������R�sp�u��ū�o�<��'���^~�����:>|����"u��Gx���8�:}�ŧ_����T�����~�鳯�ŧ�����g���Çx�޽;�����_z�����-m�|kl�������Y����r�.�@���|�����%l�h:w5U���t4��CM��	q���x7��ܢ��͎�����ҋ��[��2���EoME֐��:�X0k��T7r�����N�,��3�L)c"�E���$��e�Z���e�Rj#�/w�#�v����:�X�j�ǀ�F�B! ���6So��r����
!�� T�d���A�(�ȤȚQ!!����YSkD�=e��Unz#��I�i��^
[��Bα]�����u�=�\י��^YɪbQu�[�ma�`Иq����?���?@�h,4xж���{ܒEI$ūHY����"���ᔧ��͵���g��#N�̈:'�Lќ�������I��o��o��gr?m(���Qg���9�)�r}a!��U�i���$��F�3m�*L�u��)����+'Eo#h*Q�Y>f�O��!#��S�1%Z�hK���[��O�S�k/v���(K��F{B�S]��M�F�J 핟� �c3� ����޺��*8R(H!�����h%V��Qm�-E-��I35�tf�$
1`����+T�r] E�E�B�=��\c�UA�����W���9?Q�)���E��I�������Su!��9�r�U/��Q�p"��˲�^iJASHHc����M��D|�����'�y�����}�T|"L�Y�KM	Q����,���3�D����� 0�ё�7*d��<?e>�����ݕP"д�v�Mbo��ҙt�-j9��z�L�RRH��j��A'Y!>�[c;YQS��t�n)q�D���NoE�֮�V�ϧ`�g=�a�gK���~��Wl��+}9�t�O�i�wX1����IM�W��.#"*�z)� �
�i��8�AƑ�ƗA�ijC8�!��d��ɇ��<�	5-S	�(P��������EQn��J�a>�9~���Ñ��Ȝ6m*b�t�lWT
�S"���O���M�GK�(pj�P��Z*a[N�C�o���G"K$����GHS?�J��h�@p�C��f�SW�(a�6ӔS��)_�ʚ15cs,�/k��Bj�Oz6�7U�5�*��t��E0��]R���e
/1)�p&�'�%�X!�5�i�]��&A�`��a|�8M!�V�)NSk�B��D�wY���_T-x�r���m}�zm����h�#��$p+���88S�D#+��n��Z���)2�8��-<r�d�.+=�ψ�l�U�©�ioW�eC�ö�i|�*��[�D9����"Ȓ�g5��)g�o�V�d�T)���"�Bd�NOj�/�NdU��/�Ovۡ� ���E��ϴ��
�\oK�].&�H��;
s��#�6�>�Y�pN>�Ӿn�Q"�S>j��X�Ȋ����
M��+nZ�
�t8�G�f���ړDHvz[�n��FVb%����ȯJ���6�'eD�Q`7����p�-�#��72K���8�
Y�K�B9��]�y��D�F�]��� 7M�`̢�ґ�Nm��F�@2S���4ɟ�8U���E;�!#H�&���;3;(�2�wtd�s򍘍����|�OU�S)���U��-��8��h+2�C�W��U՛*���&T1��k9K�����J-IiZ?)��i�h�z�I�Z8�,5#�������;^S�VSN%��	����!�M��@LS���O?2�N*Q*$��q�^Ɓ'�و��4ڙ�d�K���|mW+5x�i�A�.��R��*g�n��m3c��S0��n!pd&�ZL�6�ݥ��3����)��剦��^��<w�x���	����5ŏ�����%��:���߉��9������>�l��l���.����I�x?�zػ�N���e��������ss�UȺ���|���_y����_������篖�ߪ�(G�������]������6y�|}UJ�f*�d����7q��lN�I�c���n7)ݍ ��](Iww�Zn@�z�b��y>�u}���������_���ȇP����w�^�}�����w�������O�<~|�����/_�,o^���Ս��嘮gT��i`8�)N!C6�1fl�(��jc�m���)�P̥Һ����Y�BJ�9U����``|���f�eAJ�T�錓�9,��I��k�3Kr��h��-�m3�R:Q�&%A���n��D0�Jge��J    IDATOnx�(�h���I�38�7n��u3B8��E�U��*��g�R�AHn�h�ΆS�|���������ԪI�:��>j�������g�n./N�!�s��r�����1���>?�8}��'_���w����|�ūÝ�w��^�~q����WW;��'�{������[_�^����K_��O���o�~�g?~��O>{������G{�?����}��ų�?��֯}��Ǐ�/�;�W>�>�`i-���r��rr�E�z[2Nr����Hw	r�kR�����&vC�2HʍG�St�Z�qR��ݾ�xl�\E�z�-�rw�}Z[��<���^�����<�Z��|Wo�R����i�1��!�ga�}�)�1q�D"!��RX��drq�d|2?>�o#����S�R��/�n!�p�)��=	1�s��4�����I�nc�n��ȐQ���b���LYU ԅP�q4���%qd�h���|&�TH	N ��Z�f8��vL�t�,Ƒ��o���p���G��`?xf���d:� �Y�Ta�={��q&sz�t�z��S�98Fm4��q>�h|u5l:N���r���j9)D��u���L�u�%�։�4���524���D��H�?��?��@[�ed`����
�Ie�%ޢ��A@))�ܳ=)p�ɣ�R��/Q�cZE����P-Vb�U%ǘ&P��a�KI�ᷖ�k
�0�����\(�
��A�&1ME9̪���p�����Og&�T杜]]]�ib
����e!�N�u���L�=����f�(D�>M!�d�L-�x�@���
�s@�� �EiV��-�֩%k�$eSYp��@�O�S��&�ƴ
�V��-�=j)�b���j	:�ЄP+J�f���%����@�r-��j����
>S���x��)��[���|G���R��0�L�d�H4��S���gFsz�O��1��;^��z1'ڶ�Q��
� Z%�j�H�[r
iʭᤐE��F3�q)m�i|x�ф� ��9�%e���O?�!R�%c$"4���\ʔ�^�S+����|H]�X�?��
ͱs|	�'[|Y�`r�JO��(|��/]��82-G���9�4Su4j���J_��B��4rkA&Q�_������K����Y��i�UW�t��4+!�48� �����g�j�X�����^D0T� �!h�b��R�)k[���&��`#طh:q ࿺v�8c���_���/Z�&D`�#!�u�锏�	��>~m'��VB"�R���̩7#�6'�d�Ja�e[�(6s�RhJД�F��4
���%���\�
1'��|��n�MKI�2~Ӫ�5�X����̱	�k��
���L?V�!��%�$Xõڈ������[���J��1$0���JO��h� ��s�VSX:XO�s����U�$R�-���0u�H���<�6���Dl�h�d���_i��%e�������!Ĉ��z(D�%^�:�����J��_��,�*�t̏a|:�*j��ȵg�ʊF3��@�U�n1��[`YY���Lʸ��Eq��h�j;0q!NH� �h%4I�ዶ�hȐB�[5)�U׳P�k�D�@�t�@&��h:?Z ��S�.��I�A�j�����.:H3~
��HQ��J�f)*T��)�
� 1�	n	���r0�O[*�VӤ�S�,Dá�>�b�I�΋�%b��t`"[���)΄��G05�A8�M�-�B�JP�/�4��є�����ᬕo76�@�������̤��M�����h�~�� �~{�D:5Y�F|:�L�	��KLg�R�F����o9E�d�"
��p"�7����pBZ�)�C�+����o}�s����#`]�4Ϸ�~[��}���������,���r����w��X��W����%�vp���7����ӫ��?��u�!?�yO7��U���/�u둜%,��]���??w��G�Wߒ�X�3Vg��מ|���x�����Ɂ_��ܪ:���t�[,�R�{����,��@ �)A"An�)�7�v���ry�(�^�8)N/�~��S���} ӏ$���Z��|~~�s�������>z|���ӫ�'/�]\���?x�{�d���ǜ��C�c� ��/��/������W!���ů��<љ��i�.1�r��>D4���h�����{`)�k�(���H���̘#A�r��T��E�Y���/k��A�r���\V|c�h��F�a�A+��1EcK�ݩ�0Z���L�Bu��ҁ8�C��.�y���X�h[N����w�F�*�uB9+�Ϲ7�Ûne!ӌ����Ҧ[�ҋ]'|&w}i/?�O.�{�~����������x��=�ל�<}���k�����Ã�gW���N����=ؽ��Ó뛣뗧/���'��;�~�����ţ7^\<>:<;��Ym����~�����g��Gg/.��?���|�[?��;����'><q���>�������f����s����Nѹv�X�������]�����N��7�e�K(�3#�/U�͈�k�r��4�S���g�Tr�����Cu�Tr�WC&BS��st`I���եP��D��/�K���-�Z��>����T7��Yo�D���q�nУ�<�N���Y� ��F~S�L"���4�C�� �� �v���ۭ��/�h����$*ZbS���\4��������2�r[�@�����MA"P��LKA��/1&2gB�lS�[K�X9c�Ghr=�4j	�7?@8��Nc���s��a�ۖ��?���ԭI�Y���ZQ'|;LGS:Gu�Ҧ��뾙�
A+Z͇lF�Pb�h�F5V�+�B��������$.�r	Rh9hۃ��&crd!�dNT-j�ͷ'���z�U��]��wי�+%L���ۤCT�|�v���(�oԿf�SF�aN;�(�L$�Av��q��08)��\uc�r�~Z�)P۞��h��<����uAL]�m�������S昶�)߈�O��PMS��7Z�r�;��. �����h��'ҺTq@��ԏ>)+�f�CH���J���Hy�o�B�"���(eE���) �)T��Ƥ �	f۫Jo�ղB����g�a� �e�"{E���і�a�Q���P�����@��W�ӏ���s��
�I| �m�s�hR<Fռ��xf��<58���wd��C����E+�Q�BL��
� �!R��G��Ja�i���qz�	8��~�t�q����i���N�!ř�M:�6=�0�~-ɲؔk�����"#�ֶ�m��i�����G��A4����q��G�D�"^��2)5�@H��U��ঽ�+1L��-B�ܦ��4�@���
�X���BL�+�U�o�s�8�)��8�*ZQ8�&��ř��k��8��&��Ih��V�>�|"�8@�1��	Mt��f��%��jq�e�F֊\��X
����/����������LS�8��B�Z��ܦ���3$�Uc��U!�ᔘSo3FC����h}r��L�J�M��Lo��m�	��ܩ�����ypH �� C�խ�#:�S��d၉�R������W:&S��FW'�c��c����*1���К�;#�f1Ŭ�D:,NK���r�@SL��I��Q(_���A88�*�15R�:r:8|!'�"q�� ~f?1��dK���tDK��!��*�?��7��K��V�\:Lo���&¢��<��c"����ȩ�[~���z`U�un:N�LQg�\�QYF�k�FS�%�(jl��t葁�)�(+pB�2>Z�m���!�X9�O!Nj]�R�K�u*1~�p~�盲��)�r�E���X�)�?LN������8���BH��2�p)C�T(q>�I�P���U��2 �ds���G+D��i:E�ŏS�҈ T1�qꦌ&�f)S���,�^�&]"���O������G(�'<Y#��K��Δ�V'E�L��������5ő�d�7�5ө�#
L�_߼�C�j�7�~���ig�$^�iՍ'��r��VT(+7N�8BӐ�F6���.*ܩ��
U�j�Um���;է%Y�F���p9X�W���7��tPp������W�{�>Py~�s������z-:{駟=��=��<أ�e�wu�^%�˃�w�Cs���U�������.���l�D��-�Ҟ+������%��"�w||���	�ɓ��������G�_�p����P�Mh)B���1�S��M%b
�)0�~�6��;��k��0�K�sL�(����7�!_��T���/�w�[��{�Ξ�=��W���׾��o]���廧����J��kU�W�W�W>vp�z~���W�����xܻ|��Z�L��FՁ3m�@�V�?�6
q4]J��f����¡����8RL����X���
���V6���I�f�
�PgK�(Їܳфc�iD���LAfB)��ZC�S4�I���8�q�=O��uȟ�w�N�-�I���v�BFLQ��Z�,�����b�6�f
IM��s��i���Z��	���3�b'}h�b߆VT��k]7??]nй1{�"�{~}�a���ɣ�W{�{�����t��,�ݝ×�����_~�ڛ_z�k�9>zt��ˇG�x��׿��o=8~k�����}�W?�d��o~�돏.w?|������}���勃ݳ�닣�O���o����~t�������������g.�?���Id��㺋�oĎ�k��]�-ܥ��uu,8̝�yݙ���6D�+3��Á�4"+�������@73���G��M]?�]K����Y.�.���>��{��ڭ�
�'nj�,�3�(]��(��Z�+���H�o�I��D�ae�H4Ӑ�N
8z�g#���k�K�L���ȑ�L�r�L9CC�՛,S�Br[W�s[+~E�U�=S8$�P�!�9h��L�(fRQ�)BSȄ �C���t�X�,�I���Z4���5�t�8�)��i:�����t�;֦��t��؆��t|?�U�e�PK��j�q(��5�7R�+$�/Y�s��N"m���RF`ӛ���p |
C0�D���8�B����Br��h��_���`�2Yu��,�R8��.*�V$N�_p<�hu�^S�"�i"{I
��1�k��KH
?�I_������є&�8�z�ӗ�8�p�3�3RL�EGV̎#?+e�=��pSR��B�^Y:�1�p���/���`��f�{~�B����V%�'CRFE�(k��uh��*K���!D��p�R��'x��������o��I������R$��v��d����U���+RB��є,����,$eu��L�1N"�oO���dѱ4=Xi%f�hԄ,���"� �^|����T[����1:LQ֙�#OSO@��%
��{����k��M��+OR��6'M-q��-V]Ԇ���~@ͯ=�SE�щc��Y=gM�X��F��!kmӀt�Y�)>�~�2�n4$>����ST��Bj��U��5��锈cʑX�)�)N�Bէ"�t�DS�8�F�MKI�]*WG��� #��HD�I�BEg,Z��%�֢�j�v|�'�zP�����8䪤���V+��I�87I?5�[j���IODE���cL�)2�h!m��d��e�"�V$	�"KEΚ� [��@P�z+a��E-�By*���FQ�F�Z���'1�~�LE��v8�(s���+Qh�&G��+� ���3YS�u��n�
u�`����R���	��(G�ȇ,��6m�L�*e�JS��Ψ��Y�D����u�V:蘖U�m���0:1�1�HL8�q�\�����+�䈦O��rH��ƴɜۖ��mQ�R��<H"5�/�ⷐmV�T�hZW�)̙���fRJ���j ?C�Y&
I�,���SH'�Z��"7m���.$q��F)h�uh�BZ#�Y&GbUr�Y%�kx4!S9�RR���0&�r�%
�sFY�*�ۘ~R�6�C!Bı�P���t0)7f`%"'�2SVJ~Sd�2�M��M)hlih��rgJA�1"`���#��ed�������5-E'|v�_�Z6*?�2�u�r�N�4�ht�C��Ù��e���T�Ȃ{�PbT�c�ϴrфLY:�XE8��z��\Sc�4�i���Eh5�M��E�;.�/�l��J�7��ӯ\�J�̗+:m�S�
��S��˝�4���v՚f�s���9F`K��C�"�������i�C�ES�n�c:mc&��ҧϦd�M�]����e��Y��6���P=Y4�3���QQ#q��0�ɭ����lT�ί��|� ������/]���j���9�BF
�524 g�����A��و<UF*��ҹO-�r9��Iґ-^[�ocJ�����y�#H/']�^�������>���|�kh�����1�w~}�/iz�_�.��nί�^��<�>~`<=�qM� nv��s���޾C`�����4}���s?]��ֽ�j-����׎_�<���.�[R����X��%o�P��v{h�l)yw�S೤�B~��io)�6�͂��gKj�41���wVӄ,!��.�c�+���������'6�]����.���_�;q��^|�����r������o����y����˛˺՗-҉�b�+�g�z[��e�E�?�h����n`c�F|�,e�.��6U�3��W�t&1p�Ek/��P�86�#�4LQS�:Ig��	��!���BSb�������?$�(L���۶;A�G�Tz
%��-�h�{)ȘSk��r�B�h��<��Is���
-Z�61��/ݸ�p[mB3�3�(���P���S��%z�:9~�&�������+�;�;�n�+�?!|��k����ý��_�=�=:y���������7��F�ON|6����o=y�'{{=z������g�|��}�kO><���/~��??������l����ɛo~����<�}���N_���޹�������O�������j޾G,�p��Bd�����g{s�F4�:~�Q.�tNr�5u��Z��r_+��˯˔K�iLE������K�����5��DdU_���e�i �����OQ[ˑXom�R9����n¢�ɫM�"D�u�J1j|#�E����Nj����M9���̷��G:@����5�kB�f̏P:���r3SV�U8�iN
P(&�E��pfu���)���2��(M��U��3E!,ٔ[2�eʏFg4�C\��u����-�Ә�~8��Dj�߉��҄�#�)^�d�ӛʵQ���O_�zUX�P��*�g�u�1�����	�Xg� �,�r��o|юZ���J�B����0�)fH��6-N�R�kY�3S�ó?��?{��w=��g����%(�#�nʉYW�^�5�iÑ�d�;���U4ϊ\n���H?�$}�;�1z8Z���(Ez��t��	�8����F�D:
�Rj�T]dS8'_�9s��E����"é�n��a�G�B�%�
�BL������K9�U�Qⷖ��z�s8h�:��v,Z�Mq8Z�W�_3)c]!9�q�A��t#��B�����+�,�8J�6ASH��1���e�iC��:��h�bćg�)�K�;�R�f��Yg�6�(��է�>����Qd4�CMRzs,샊��-�r8p)Be����������"�ԪD\����=o��'ҁ��VT
_V���l�sc>?�	'�U��6|��Z����;�P�R)�v�h�G���i͠�)p��4;�Ne���	5 �E�L�O�n�i�M3��#�LQL8C���b�J>}�DN�	�2�Z2���''f#�5�����aj�B�u� ��V%�؆�/AK���빊��j/A�)CR��bgE8�c��:)�)��)�*5��p�0�XV�����sV`i8Y���Q�_V�4+�Y�1Ki!��ሚn�Dp���&/j�eJ*dvrx~Ld��oZWF/c��N�|�p�Rh��
�m�rx��Q��    IDAT:�7���(����'��y:��'�!�r��@�Fʙi�v �N4)�4e�"$R:�i}�S�8�8-D9�*��E�L4QH
��h�G������S�gj:��9�1MqX807�	'��!��Z���)��(�L�(���LS�o���A�,Zwf7D��%'�X3)��N�|,>����0���V����N)@L#�R�9����tfЬ ���3���g-4�����~&kh�§W��JS�Y������am�E�X��MM�r����L
�B�D
�n��A!:��p�`�f"�ImϢʅᄴ�3MAN3Δ�[��6ڟ��!"@�7>#�l)�K�Zґc�`d�ks�9UQ=MU�li|��D�ӵ�@��E�� Y
-�_WUD����n�@���3�)�)�O��L98�B�ۮB�`DkOD�*�mB�BE�[��_���ㄤcd��Gu�C�#��!R���`�B���`��jOz��4�r ۢeId�����I-�X�Ò�5����D;����!�[�6��Rf5|M���)��J州���Z'm���)��6��:��� ��d����I��gV��6H����Odc�D�['�Pc���Bei!A�:5���8�rq8��P>�2S��tѾ.��&m�,��\z���������{�>w$�����=��,�9q�{k�?r�u�'�vvO}��]�h��z!:;����ڷ�����0gļ�w�����y��f�D�FU���z���?^����[���O>��½@.�nO	���eO�H�Q��ۑ����SN.���,����;e����]2��4@��<�������H����ݟ�M����ϯ.�.v�|#�����ˣ��O?}��?]���`����ϟ���},v��Ý��w�������O�_]\���zp�ok:�
����,����ր�ڄm?֮�hm�V��֞;��m!��ڽ�-�h���"L��%�e��a�8rWli'���9�8�*��)�J���hC�����]W���iQH��Y��%a��G ��٢F��a��JL⶜���3!N"�F�tR�`�D9Z5�1�m��V�r���%�G*�,��#�NJ{��_v��[>P(&g�hl�pd�b��� Kw��÷�)��d�fߜ����თ�:�Wh��������/���������ӝˋ������O�>;�w~������O��Ϟ?y���}�K�>:�~~�ዛ���_�̋�����ǿx��|�_9y�[�o�������>}���O|}�n�z�-%���7���W�mh-�~��.p�S�7k䰹&��g+�n�p�7b�5i�Q�5݄L͔x�I�e�gS��.�z�Ѷ\4WT�x���u%-OƯpwE�9Ǩ3H|�n��WU��l�;:�AY��ߪ��Ȁ-�ik����,2�
���Bh9J�eK����|:%
9N)���od�L4���BF���~�V��F�^~�h�V��1U��Bʃ��� ���0��8u1��̏_ҡ�#�g|�ɟr�4�:X��$l�8pYq(�J遱i"�K�)��|vJ,U׿эÈq���y>cQ��u+ʡ,��%�W%=�;��R����7�˒��	V���~u�R�"��3����MA��E/R�G������������%Tc����Ha��U�5�V�%���EÁ��(�����f��T�>�����0���pe�իKG?h���2eB�ã�2��#_��J3Su�-��d9� VD�P���Z��D���c�օ҈	16���l�]�	)�Q��w��{����9�\��2>>g)�:�i�������6����^L��N�>|i��'�Ib��<�^�/g��<���h��RK���1�B�AV'hj���DN����U[�Nj|�l���I�Y���Duk�:Q���Mvp��2{i�:����_}�q��)Фf���pE5�g��4Mg7Z�_��_תǍjQk]�^kE�H��<�:~;@�i�)s�զ�7��+���g�B���H)J� �bW�5i��.>�Z�8�V�1���!�&�c*:�i:�f$�:�B��꭮�gC%iL�4��4?���P�߆�l��6���J�YunZ[��u����hd�'�� �^�M�.�UA
SW9N���S�t�3��>C�&��a9�$�,�P������4�tR�I����#kJVJ���{Y���5�@�d!	��5�\�
X]���y���E���ٞ�8mˈ׃��-�B��c-Ah�2N[��C��ڐ��L?P
�=�O�r�F�DD�t#����#K_H�Af:̵�r��clE�)�w�'�O�Ѵ�u�a���B�g?qL-���Fd#��H$�(�U�_��:L�Im��Ԫ,|-U8��S��i ��%B�	M����0[�Ш���]��տ�N�O�X.?�~Y�59��-�öU&H��h1���j[?�!���nd�Q��@pH�7]�����# /�k4M4`c2K��+�A���QbY@Ә9B�^]��E`��O����pO3c���9�Y�q�E����6�CSք�RΨEk7JD.4:���iN?S�ݘ&�D)�R�
��l�f�t�JI֞�|�E�$�R8II�W�S�� |���6�#�C�S�IB�OS��� 3e��w���T�:�|8��M�Y��$p��j�
�i4>'�5r{��DX��En+�j7঳3	6⋲Q�d)�EF�H��bĩ�|�vc�;i�ݦC�~�9jqd9.-m�����,N=�v��;RR�v�K�-\�1~=�ӘF�v�������F`��N�
-ɫN!~��`�V~p�p�Ox�K�u*N
��72�6�f[W��_�p�_�B@LY���*N��7e���1��F9�1�Rq�*ʥ�������cx�o�L:'+Q�#7����,�l�VJEx��b��1�N:b��z_��/h����G5=�\*��/=��ݳζ����n�O5���CG�,wq�磇7{7���΋哚;�n�==��:���W�j)�ә���y�u�c_^�ɣ�Ã�w�}�ѓ��'����B� U�)Ŵ[`���c-:{eբ�9�ʅ��E� ����qL>�]L%:���F�}	���e��9v�ov|a���r��ۋ݃�/>��C�p�uyv��M7� �W����Z�s��G�;{�L�/Ο�{�ꙧ/�]>��~�vy��֛?K֤�X+��,�SG��ܨ[�=�L!�pr�O�S�����U��+��x�]���~�XY�`n�tFp���,�0|����E���B�YhjUg�X��8����ꍣ?��Lq��1�B-?'}�6%)H���CV��S"�!4��T��ՉN���x�d=� ��8�-�\��K7e�p"���ȟ�^@�����8;]���̻󎿥�ӛ�/�<~�����+���P]�_����|}�rw���ɫ�����_~��?���?����'?��G?;z����������旟����_~������x��?zv����/��o~��������~���٫/�u��~�m�y-���7�Vљl�����"����6¼��mfY6��\)�I��̻�;Ґ���w�Tnn�Hwך���p~����e�nغs�+�ۿ�ۢ��s�(-��b�����oձز��s>5��e�8*�x�F(���V�G �O�8AJH>dp�R�/�)K-�n:LS�)Y��4!m�\���\��׾�q���BƟ,Q�gjF
�86��dȚ���P���5�B��R3ũCSά´P"��8r�Ӣժ��)}�?)Crڄ�0#7&.���l5�6
�y���O;ㄔ�A��㏣��ѩ������|���<G�zP���5Q{�hr�B�"�f�2�(}8f\:MS/�un�
�52|�D82�.�b!m�J'[z�|���i��H$?e��zd���RN]������W~E�O��J�E��������f�T(�Iw��&�c:{��F�L�����7&=mu��C6`���&%k�j�ru�j�Z8�8B��+dxQ��0��D6E�"f����.?S���w��dUAE��(�G�6(H�(�s��s!w]F �:��Qj����M���!d;[�v[����)$�t�Gp\�0 �בҊ����}Cճ�	ߞ���ͦ1�"��d��2)�Uj���|����u�F���(M�cE��,0>D.2�)�=�Q��-s��!��25_V%�.��:�vd��o���u�½��:��3�Y���j B��G���ǽ���i�GuRJ�4=08D.S�3���ҍRTьh_u��]��B��+�i��X�Dd��jp#�J'5k^o��lu� �a8�ㄈbj�A��X�vSW� V@���*4S#��P4���Y�0��9-��5�p�5�8U�m�ڎ���1!�vl�x]#�j55��Y������/�]J|S֢�O'-�r8p�oZ�tU�*U7���|H���VmL!�Q�5R�h�V:��JԼA(~��W�V1�8ˌ?�I�m!�"Y��oL3ӺjZr���(=��^ې��ݫ)��pB�Z���,�vO���"o��v�sp4Pz�T���(����*+xY3� �wG�C�rZ�Prck�1͐K��V7�7�	�E	N��S�dQ�����Q��#��,��	���	��8p�)�ϙd��@L{]������YNu�X�Nd�Z�t��b�y�^b��q(pp"$UH8-E�+~���p����,���m���SK���dY24fjD0zr��r&w��˅�Qs\�'o]B���B��D(�c�d	�sm�'���Lk�?���t���q{jѩh��krZ��)pZZU��{
��J�)�#"�5V�/�ߎ�܎9Z�'��T�l�Y���O��So��
��i�D6���-)��×�8�)4=u�8���X臯�88-�*�I�D�W�4�������C���A1<))c-E�`
I�-v�LK�Gh�9Se��O�[����-����C�($���q:O��yā�EW�-(�	i�	b��1"ty��Y��
q�iu���,�#$U�Q���&����о�F�V:���c#�!�`�~�P:���id��$_H/j#�� ?2_t���@#DV"Ԅ�B�Jk��||V:2�M"dL����G>D]N�N:���M��i))������/�B���3�U��a�����[�Z���{����s��[��>�N�K�̝_��noףG��z����G��s���lڲī��>}���ʇ����\'�g��g�d���uWD�}����l/..O=<��׿��G��/�鰱-2eč�zvj���-�V��������[�;���(��������
�~w��%��:
��T��GT��C�n ���Op�_���C��1'���Է������^}��W�/N^s��\�-����QL�=8����=�x�ū����W����������Nr��)�*d�t�kdB8�hh�t�v��Xzj�����l`:�������:Q��a8"�(�Z�$��Q�)��q0'�M/:�
��X⤯�U�PREg܂[|+�ojb���;�Q��%p��6�Op�d҇?�9�"�8��HMh�r��� ;��t&ʙ�9�KwG���''�� �*���Eh}-�D�\>Zu�<�������Tg;{�w��է�/�?�{x���������g7�//��=��?x����'���׮�/N_�_��K���/��y���������t����������÷^]���/�w>y��_>>:�t������7������K��u����>���Ѕ�K��p��Uۭg.&�s���R!���Y�.h��{#Ff� �QEu�GWEw/�݀�S��r�E��t�_��=j$�N�b.�i��?G���Q�L+�����|a�'
��v��w�5{I�kmDR����|rڣ��@����)�qݚⷄ��0�BF:�FH�BFֶ�*]�A�U��[Z�%�b-����|����j�Tϖ	!�Q�Kdose��ɚj>�פ��.��顽-E:����1V�X"S�)^zmt�!�k����u� �I�h�����HJ���7�>LV�#"��8{zl�@�2�*D��Q����e�#Cn����������$*G->3l��:�3Y�җګA� 3RLQ#)�@D�X+,_2鉈����{^�����U8���)Z�Ԥ���d!��XN�N����H'�D=,[|�O��(��>�i���(��rU���I7Ҭ1�jOKD4̀�)� ��4��!�F
8B��@T)Dʫ�l��0�c���T�SJ#�(�8�������i
Gp]֌,!NW`
v�'8�%U:)F�
7�1�g��2!����>����r;�c&$�Ͽ�%(]VG�(d�?�!Kةb
�ԘZ����/j�/��r�7"�F �8�r��!bS#����9͜EUj�F)*
q<���{�繣�F��H�#ˋ�U���co�u�y���}t[9/7��@��v��/�'��mS4�(�R��[��� �O���O�(Ԣ��*�d�����v���2����:UdymjIT����J@Tj	G!c ��VYBƉ���Ñ�ꄓ	E��Z!r����H4`S!�QX9c"F�mW!�d�C�E��T�݀������i�
ᴊrI���8�[f`�F!��$g��#3�U�;7�Gٱ洁�Jb�!t���H���>��B8�0C��Tbڦ���p��0�h�R��2Ն��R��mY�8h�U��`�q�c��2��R�=��%�5`���FA")`��	��hJg,Z��$k,ј�/��eR0�3>�)_�,��D��_"ۉi�d��+yE �$2HW��MȒ�ӵ1~#>�R�|�V�ě��� P�2�������G*A���F�p��5���D�M!����tR-M��8|����Gk��D�\W��DS���o��u:Q�t���C���@�"ˁ̪q��sjo��̒!�Shu�G�O!��ɔ-W��4Ms&Z'r��d�pcY�g��cZ������:�੉Ve�8�j�45��Ra��	���PY��롃L�h|c��(�r��:G�c�-.1��%^��p#K�m
B�9�d��B���eV9Zg�t)��!Ӭ�pS",�1��l9�j�˭nc���4�rȶ
DJ�h��/ݬS>B�h����%�� ��!��B�R�B�1��W��z r��P4g�t��zK��U��Iy�Pc�h��|�V@�U��T��2l��Z9FY)�2w;�н�']�^*mNi
u޺��2��
�;`���Ds�􍬔��č���_-x�F��F����k��g!�RdS��cnG!Sd�0���P:?��U��I� �w��H�����7�����[��O�u"�Fi�6��T	S##^�i-�-�(���� �KV?T'U�u��*E1�B"4Yjp6�p~|NG���e���I	���dy"��s���K�W��\>��L�8�������`���E�Y��X�\=8:Ђg�G~�8p�^� �3�����kw}�ҋ�3�p����g��֫�c�[�Ϻ�X�6ĭw=_�z��W�8:X~�q���(�N"�~�'=�̢�n#�	YT�9CR0��p���7�7��q�����~W��0kw˿�.��N���ɬHK�n��*���/|s��\���Kw�>������������gמ�\\���/�c_�{�[-}�������v�O�?��ɓ���,�E�
1}�"��R��K�7�Yz�S�Ҕ� �T��q~�RKGԔ�%�O��K_)��p'����]�i��d��&��%��6�?�:�������x���b2H͌�iQ��٢8��+]:NmLn�}���/%���M�P���p�D ���/1���,�9���{�����F�Lg;Uׁ���^��12�F|Y�5ɇW�H
��^�_z���׿�闞�>����C�E{yz�����?��=�_��o~������љ״/���8�7�\A<<xx��?9|������z��    IDAT�O��`�� N<��|��=|����#w�O����������ͳKW���^>���'��������~˅����0Զ+�ӕiՔcl\�:�-غ�ÄO�l�L"p�o�%W:�>,��o�#�&���᫒���a�R�V�]Z�7~�� ?���|^E��	�<9��������B�����C:%u�Z*s=vˍ$d4Sxm�dV!e끠	U7��)��ow�W��kl�L����Dx�rZ#>&����R�'D�Q�G��#W2q�i��7�h�����<Acj��f��C���]3��++�Y&��P>}|�
��P��B��NMS��1JR:��f��G�H©"2)������w�<H���<�������	��CMQ��HG�FY�+ǈՕ(����0�[�.�x9����K�f��H���J/Bw�+q���W"dM�tX��:���=��;f<����W�W�H֏S�;��#Aj-�hǔ����e��_��!A��-���)~�w�4��}��3�>[��������R|Uj��5��8��9R�J�1S���e
7�l�jqb������-_�]*�ƌ��NEH~��#��U���g���)�T�ҜW]�j�S	��f��,%�+�GV�Ģ��C5�.hpG�o��C�-�S!"����q���%�#S�/��BS
�X3LQY��5����t9&�EqZ�($���^>`꣇@S�j�Z�;���!��ZB^/NQ�������ar\0k��w��]�tnj�!^�|��ٛo�IMHuO@�]3m�����!�
)�=[.DE�������-Y�N����wgN����+���BMR�QN�r%��AF�a-�էPӲj�,�IϹ7F�EF�	�O�J�1D�����9c'0��{��%��-�40��Juq�8�ɶ�@#�8��_4q� ��a�Dj��S'6�o��gH���(��&b
��9|&z��V�I�v�cڹ�!�8)���''�V9�蠵(�2��2�,8Nʣ�U�Q�8��!%֞�m�ԕ-g��2��i��?���0#b2Hc�#���.D���Jg�N
A(g4�q8c50SN���u�Ӑ��P�z��^c��A(Z�*V�t(�̢JO���"��?���o]�tX���0B����P���i+���8�"1"�C��ͨ���)�H?��PE �=,�Ԝ'���dkF��»�+O��D�6j`QY�R��<�p"�#�h 2k��$����f�"?P�p�~��&KHxQHN��H�Ɵ)+d�4��vuj�'�������CB�|΄F_Wq�E�o�G�IP�q���Ӻ*��B��i��EkU��Om
�S�`f��r���!��P|�(P4~U��~���嶽��,�m��)mڊ(T�,�d���i]dsf�n'C��F�J�L����L5�oz/d�BD8@�[N�#H�R.�$Ƈ�z(K�3���pV��A4Bs�i8RǴ8�1�'@jU���P��ݎ�8�'�"ԕ�u& �iāǩ��8G��� 3�l�D� �hd␅tbL9H),�x�N{�h��|BS)��mȝp�0���'R]"�������oE~�y뭷d�l�q*d
�B
����J��O�~)��]�p��Z�1BG��jf+QHF"��@~O�m�Ŵ�t%��x8��U�2g���g8M����#�}f����J\���J�����*���lR��ݦ^[,/F�@Z�Z6�ף�n�����H�P=꼾ٽ���˹G{4�)t���}_O{�s���^{p���|���C��]Zs
��NoOK[ϋ�g>���姟>[:�W��o��l��S��Tnٝ�U�v9�ǭ�%�����ߦ�0{�~�_��7��Jg������7��r��N�gY�<�}��G'��8?�̫�.���o�����^=|�����gp^�� ��^��ۧ��֚��~|�s�����kߨ�ҍwu\���'ɷרV�Eۇ��V{�}(*����Advl|H"���O-x�1_TKi�42R8�hF~�[���)R�o��"o���#�Fjp�����=�tM�^�D������_4��o�'8�������[����B�6&�É)���r{���Ҷ��X�����oe�>�i=���;�[�(���p�C	O�m�9$N"�SB�Z����o<}x��/���ǉo^]?;{��ǿ���o~�#~|��߂�s�������?��
}�����k���w�t�C+�_���8��K�/Ϯ?���\>��S�?���n.^�~���������7�}���������sߞ����劤C/7m�
�ٸ\D�O������!�����Y�D�\4߬鶿���8�=�v9M����)܏%.�j����?�q?��%B�1=eX� ��8����%W��M+��b�ġ����,��Z?GIQ!����
�B�Dc ?�2jUD�������G{�c:�!I�@DeQ� �_H� %rL���(G��hx� �.����RzG�/=�TL���sp����׽��v]u?��pb���JPE��h!Z��t��!z4�����B��T�rlW�A~��y�g��9ë�)���1�7~c̹�^���އ�ic%Rㄔ"��(�[�(�`d������/�ϑk���� ��\Q�́� Ĕ[���Q �<�:������S�/�qb�-�~wZr��0���F��!�>��IP��Oh���:a�����rS8>��Y�\��q��  ��w>[���HɃ+/�7�x�o��o�z�-���&����5ϧ@�r���d��"}���T-�E�3šfʟR�&(�����R���$
��g�sT$H�h����ʬ���MU��+G'>�Tj��lW	4=Ha�k����] �z���|
��ơ��E+]-��u�7�R����1��k��tiF�I�͜`R�&_�#3�F�:�d���I�J(D�Vk�l��KFu�d!|�||��~L5���SH3��OD.2�)ӃQ	�?���t��"ʇ���S:Bߏ��Y�D���8��D`��`Q��8�X~k�-�oE��`9�	^����B���_���&�z �ۢ.M?k�DGn3k�Z]�ɦ4"|��M�f���5���"�7�G�-M��)�����R,�ڭT9 ZbF�Q���c�j��D�&pJ˥/�À����L����q0���-]���Ҵ�K�ϴ(��}]�h�s��d_z��^��ӈc:#'�1�Z@�Lr�©�F��)]�3�R���t� ����Q�B�i����W�L<���!Ԣ����=�Fd>�)
LG����/��k6� 8-y����W�Ö��*
�D�0�gt&%$~)IY~;�B���B�QkE�m)�����lMN"b�2�!�kZ�{�i��Vwg'~cj�����*G��76Mt e!p�V���L�8��t
���p8@#���ȩ��YT�6�Q�iֹ�:�r�2%��\Y>�8�5N._�p`ʦ!3&n:٦�r�גns�FF؃ua�d��Ȇ0�Ƨ��k���@D�k�P�B���$5#C�9Y&Ÿ�/��)�!�Ij-AHQ�� l�m��9���S�ɚ����KB�pQ��(���jk)0��ōNRt8��͘�_��0m��nKcΈ9[�1uۜ�IǷ^�A�T� �c��t��!!��m�S3bF�75
�9v�K��J�g��%!�q�C�$-´��ۨ:�a�h!��Y�,qΐ!3�Hi
�">��P��"�W@f:���UD+1'�i8�C�P�VD*��)+�Aft09[p��F4�1�_�*J,Z��i�𳑭��	��*����!�j
���D�h"�U ؊zmF�H4ʚB�/M���AhZ�EG�<Oy:�Ri�8r���	�ڦ D�L�+���I$rSH)u�oFH����oX�I�N͊
��o�Z�*�Iq�#s�oa��	J䳘���x����k{�Ɏ�U���҇�p:|�Z�]K�`xGؔ��S) !
A�H���0����,���qG���m76|��p�����K�>��ao|������3*����t��ǒ<�ܪ\_]�y����>y����|p��ރ{�Oe���b���� �����q:���.�t��M�Ã�Ga��	�m�:��ې+�߲?�t��ɤoʷ��j/p4���́{+ݫ��V�Ψ���[uKր1A��mQ�=�=9����_^}x��m>�H����o������=w��=�/>���2O��Nz$zx������?����g�q{~��g!�ܽ��Q�e2�6�s��m���y�Ǆ$H�OJ"�m4BX!&2jBM��5X��)%�%��!r�\�����-ΏS-S���8)��'��h!Y>C����dD�}��d�1j#Ъ����ƗԆ�)w�S��pS6>�Tncj��E���O��=^�B�Z����y_(YN~�
5��	n��~�ju4��Fjt����^,B�	v,:	#�皯|��_��/���?���������?���w~�??|���/~�~����W���_�xv���~����>�^�������|��'���:�~���˃�KK������������l}��3M%\v�u桟�?z������~��w���jc��W���	q [��Y����桬^��H�Pc+⸽�b�B�Z�C��}Z|�F\ԅ��O?�%ʢ G��(T�@v�R����>�)E�M��~��W������u��N�$g��|Y�Q�bZm�-h�m��V.Em�.�@Q�FF�r�|%0�k���h��˲��m��u�Y�T�'�d� �3j�_T��c�(M��~�BF"���wh�J���T'�Q��3]��[d�Heˑ�s��4�H/+���jŬ�d�@�c�X�q��aRL�mT+�R4�g��>�T�(�Yu[�"P���(�TI�i`tr{���~�ٌ�Q������gHΓ��p�P�ۈ�ڴ���	�����zM�#�(H?�T״B��8�i���t^{8e��F��(�%`��������+��|j@=��5�E�\/m#�]q�Y��CQ�Բ�}��U��7h�B�(���
őE�������U�?�����׾���|�;��VhFi���@>���Q�'B
BBe��l[��e!GK�ko��T����Y��u��Q������ۓ�]��ǜD>��U���j����SFL%:p�ES'��O_Q/��^/ҥ8p�.��~`���\3����a����aJ��4��e"��##HA�VVݎ`�h%r�T~��!�g�p�A��l�k?#�]��׿��b�הo���7@|"�DԢ$��u�r��x���q>�ɢ!�C�o�F�ӢZ~k졦����쀞�A��G�f��&�����c�ҏ�r�M�Djāc�B
��Ĕ�e߾�0YaMd%��0Z�h#%�����Bp�k�!J$E��JtNڐ
�q��.� �PL�*�Đ@ngY��V���^����_op4��4`j�g4��E��|ΔGs>��I�C�Mo��G0�\�-%&G�E9����Zj \J�D�QV�i�&-�zk��ߕ*Ј�t��H����F����0hY�ږ�D#�!��r8���"LK��6�|����C����eQs�uU:rW(��҇�����r�R6ͤ䔒�Q	L&:�L� �#�mzVHJױ��銣�1K��)0!x�E�Ǚ�Ȣ�8�p�����7����!բPt�"	�0��iQ��)��B��c1+ڱ�K��N��Z������r��Ԇ�Q:Hq�R�#�f���>��N��A��2
Y�F
�jQ�E4�Z"e��-<A�8��Zc�E��f�Y)C�����Ob�����_KY��2E_J��>V�wW�4�SK�H�VWh��K
���V�6NR���<$P�p���CZl~��M��8���W��Q���̴��PD�i�Y�S�x��k�fJI�\'�ǁ#�&hd�7��������n!B����[f�&
d��9�B�o�7�^����Mc��0��[�Va-�BDFX3����,)
94)��g�W�3�D��rg��
!�7J
�����@�3d
�Ȫ�v`�h��kN�n��D���RdUe��j��a�YSR�̦e�y�I�ؔ���M�!hZ"���>�{%+bB�2��?h��JsX�>}Q
�CG�ü��ҡi���'Z�,�#�-���ӀS��S�_K4&*]� C��~#r<���U �D6�s�PL:����
Б���y@�/��up���>��Y�x�)�/����'�/o.�N|��sg��}��c�[U	�q^^��>{�cG�����Ӈ����O�s���9}��ƫB��ko���<���-^�Ѻ]p�	}鋿����Ϟ?|u��n�����X��]��1�ͱE��l;ci9s���@D����9-�s��%�����S�)�0)4����>�������յխ�s�9>��W�=8�ַ�����_}���g����lӥ��飘'�n���<y����z����l���Vz��T�ir;Xk��v±�6��Иh��F\'-�=n*٘�&p;l2k�k�f�T�� �����yS�J�J�2N!Nu��!�$!f���)�LU��-�qd��ΟZ�lڸn��*LF�_�=s�Q�}��a6'|�[T�ؾ��|JOb)�Z��jC�O�8u�P�@��8,$pM8C[	w)ÄLnG0���o/�ጸ�"Ǫ�с���ϼ..n����#���WN�>~����������?8~�g��w~�KON�������C}����w������|��_<��{�7g��K����gG�n�>񹣛��kׄK�B������}xݭK"��Uw=�.=�#���e�v�2�K��j�� FQ��%�@�.FV!8�	�V�������g���bu�c}��cUt"��c���ؕ��Rq寿����&�#ԥˢz�ԁE���2BЌ@)�'�,�&�����!e�u��6�L�� �&��q׉�q�hX����|&!)Sf������
T���[����ʹ�Q�h8|��t�k5V�!B8�����?� 1e�,�Y�F|�5�#�̇��5J��i���82v�U��z��:T��Pfu�\��<0�|©�%�	��L}Ƀ��R�͸_�хCO!k!��L]>D��)�@�3M.�ً���$�K�-BK�T"�7���7b!pfʗ��a8I�E�E�뗛�S؞�X�?��?��Y�v:���M0Jd@f�]r��D�ho� m�ny�i�&���.�ѻ�o�5�!Ќ�paB�[χ��@j��E_hVM��gx4&�o}�[z6U���pc-!���($Q�*�h�BD";��{�t z�9�v�&�P'�G�ZMr���U�^?�d���3�~���;��� ��q��:�P�΄R�ej�F��:Nm�;ppj����3����8RT"<�є!�bC��f���%�+'�/�A(��=��9@~N�(�>��Ieu��p(�I|���)�r:�;��@��,
��
S��{b}�RÎ�u1��G��|�M�)xDJ�Ch�Ǚ�&=δ-@�0����r1�8�9�6�3K��6Ǌte*������m�Ƣ�j
��ڒn�C�0��N�����vA�� �R|����XQ`=(đ[:&$f]��@���fʧ��m�n���lZcF�����e�o�D>�R�̴�	�p>�׶��	i�)�iTM�0�i,~)F�f�H��L7���h��L�*Me��vF��	��#O*q!���݈ 1!�L���:yR3��@�[���*R��n:U�H<~:@6k�HA�(���s�R�s��P�"�*
���v���,?r�E��p�fF��/�&[;f:��8c녧`�� Ʋ�7V��B"ÛU]"}��V�p땈-�}��t��tȦ�G�fQc�M���Kh�#�a�%Xb8�i�d����2��N&��V�-cR����v��+`��b���G5    IDAT@Y��-�P)�Bc�^�6D�ik��$� !��:<��<��p���b��+�|��K�Od��'}�"�M�c�yU-)�X�5�eL0P�����E�,R���R�疷hBħ�}3S̖P��ƪ���X�p�;�z��[Q�Jt�D�$�I�cZ�V�@cիb�!>�BM�K!U"��"L'�S�U4UW"j	����d#�h��,�?#����%��C�EkFT_��JO�)�tx�3v�3�gX��S�n=�܈#���2����9~HӪ˭����F��|�`R�N! �~��DbZN\4#Nj%��^M�tL
�@f+谘BZ��8�� ��i������UI�є��N"�#s�
�Ը� ��O:P3r��J�*B�FN�*��G�D"���t��NS#N���ۑˍ3�8p�#��FV'�
q�F:E�����u�'é���Y���i�%2��tL��ړة.���hj�[TE!~j���r���r�z���*]�s�#d���'~:��#%����+����5I�n;�{�`JG+Tz�,`Y�h{4&���<ބm��Qw�==\�?�x�p�5�9涙�K~m��n�	]ލ&�������o�����s�����S�'�G'�P����/Ϯ�|�����O_D{������ŵ���{�������ɤe��ۢ�Ճ/�����������}���ܼ��kW�?�5e'����K�nc�1C�M�����W"�hg�Հ�UY׺~hvr����#��r$)��w��i��/�=v��>����.�<+v`|������������z��o���^7�n�ݻ��N��'�W=�zxx����o��G?��{���K�m:��"��h���9�!V�R�rHI�I-��9q�h�"4�tB��s�BY:#���5�Y-d��))Ӷ(<��\E�ĩ>���g�Б?�i�?�bfC3�����*8]Af�|�HY1��p�����K��5%R�W�����1�.��j�qGs���{�P�����t��L"%�6�F�\�i�1uL�kЭ?[?-\��]��?8��}�<��ӛ�_}�����ǻ?q��w����}����9��N�幯�vm�9����e}~y�n;V�o���߿�+��/|2��+O������?�������n �H�cQ]TY���H�5�v��a*ĺ��Z��k���>k�b;Ӷ`�S�|��C��l��?�\19.q>��N�u�;>��7�����n�{��'C֝S[l=u������H�X�����aTX݈_+�^<�\Gn��T�خm��n��45��d�2�\)p�$�;�@��$�fi�pіVu1J!�o9F��J��!���N*��,�@Ynj%�!�ȹ(���_Vˉ�׳(���\�(�`:��&�Ä���R ��"�CL���,Z�h�4����lJ�#}r9��h�B�h^3|4Vn���%d��m8A米��w��y���]��?g���D�/��j�+-�)J��S��|�LGHĨĖ��z�az����'�F��kZ�H3�z�.%�\)m�����.�Ǻ�'y.�7�7�����R3Z��Xh�a>ugu!��8�V��j@
�);�!���s�FS�ķ�v��9B�	4m;�t!�p�@J�BJ�<�@�Z��?��?�#�6�0�Q�9� �Z2��i���[����=RW�p�Z�S�ق﹣G�t:j�h,_��d8���_QU���Z�b���nϙ���5��%�+�T����
�խ%ffu-�HA�U�s:��I�AH�Z�	Asb���a:N�J�ј�y�!'"ZW����u�Q�Q(E�0��!|[������@��m�s��%*G�=���'�@�[;^Y~ +d���B�z����_x�Q���"r/�ׂMVK]�M���lT�z�Jbt�UD�"��� &��8���ES%2�f/:���,d7�S�J�	��iTZ�d
�r�T�Ө�6��>5�Q�tRB��p �(>�K�m1��ЌR8k�X��L��t��m�?]�SҔR'B��"H XQ��9��pJ���Tzˌo��LAk���5V����;-AZ#$&��L��=���w�tU=��iփY�Կ�� ��2�ɩ'>���:�A갩P=��3x�S��7S�i�n�K�O�9xgHkGC U��1��~�ES�p(`���O-�͘&�hc�4C�Mi��|z%D˄��%��i-5S��}0�%.e�9��jY�RfO�\��O�F�Ƅ�\�Z8�L�8r��t��''�1�&��Y��GY�1��h5�'3�I��8Y!���k)�ik��K1���p贐
�+���m���J��5^E %�A�Y�)�ϩa�R�����IOj��JL�S�QJ�M3�>�!����"w�9֫V��mQ�JK�2n�'������Ԍ�r�&4�)�)�@#��-�h�K�83�v�jM�#��鬢=���d��Y��]zRF6ȯ��Af�65R&�Y�wx�[��&هঔ��>4x~��bZ�)�rc���R����v��K���f���4�Q8ˉ�]���$b�	�+~�-�?󁌣J�4q$�T��7��*�gB��G.�ȯ4��|��eL�Be%)'�Z*W�,k�819�&]��N�\~��Ʋ4��epȀh��s��ե`�����s*
�7��SJ����fK���Y���7!VW�8E�k�sR�US��@cxY��HP��q:���3u!�I�R済28><�,�j�I�0#�rL��J�G6�΀�.��c���%�6� Q0�D�n)x���	͛ ������4#�F�r/:Qd��Z��1��6�=�^�)>��Zr!-n�
�9�����h��qR�|�������(Х'kN�m�;`�?��YN��:�>F;��`��wϮ>=�4���#�G�g|�,e�O]����5��?1�a��m���k|)�/��|tv���������P�YT������j��#U��SI6o�ÉQm�n�=�Ļ����7?x���V���]\^8k'��oi��b�Ŕf�bc���}�HNH!����(7Fp�vIӇ�ܵ� P���~hB�Gє�Z��˫��2��c�=9;�7�|�����=y�����ol�o89^<w�����o>~v�{'?{~���&�����lj��[Wk�4��ُ-�BD��逥1��>����t@��=@��ݜ=h��||��KI�(<r �Dsڥ��9,&�}�*�!CnZ�����@�X
<_��� %��~:�$2��rIU�3x���,��6��V�'<AYt��C�,}R^����sp�rFyZ�������L��g�1�k�����4dt��̸w?��-rx�y����'�]?O�]�T�y�����E�����Z�����᫧��O�>~������ˋ�H���[?ݜ�����ً�؇?]M�����O�=΋u屖��sW 7O���3��g�o���]���T�Gy������i���	���E�4�L)�ڀ�!��ΕкЀv����ĺ���'Y���:��L����=�	���t>h�i��-��[��7�ڪK�k�e��$B�0�D)��˂(��5T�An��2)�
�[�'��-ɂ�N������;�ڈ0!4�L���%!�6�9��U8���1*��*|�)+�`�U�������~$�i��Z`Y|&�8D�t�`K�b�.T�B�%��l�K�~��E45
�~`��߯+M8�b���lt(�4�I�΁4Z�D`{(R�/�!@��NH�%�����y�'1�h�6��K�T�h�M�l���F��$"9!��<^���g?{����"7j	GHϩ��o��8�G�wp5
Y�V-��76��J���������`�H1ؐ���'�F8)�t�h=��uD-�uk2��Ti	R ̹Z�0ʂk�X.\?����$K�18�'d��S��3Պ&�����8�a8��#d�E����qC���[�e�����LǤ��(Wh���L�kWET��W0Wa�.�TN$w=�u4�p�/�u8j�Th�ooh	R	��.!��w�S��*d$�&�;�W�*)C� ��,�n�¡V��_) s0�g�a�S�H��X#�,�h
�cT�T��B���ʯh:��CȷW#����ײǓm���*z�:LN���z�ra�!N�6VW*Rs|��w^�鍎*�L�8r�jR�+��,e�Ľ�9�3{?r+BP�H�4$'���H�2)�sD�������C�(]�9��Cg��7���� 5%H6�n���%�r��ߌ/�H*��A�/*$��J�넃c�S���Q�F�]� �M9��є�j��%��� ٚ4�#��Tј��Z�Q6Eh+��K����q���F�…����	G�+��h 5�Q������@S>'df�J���-��t��0uˊ A@���rd�����8�p��୥6p���1��4���Fe�e�8{b�&1ASNYY�q�.�&�Q"��D�#+�p�@Y��8Ζ�d�nʫ���H������o�/%`�D˯%�h�6!�1��ߴBMCJO��6'�R�7��� 8+��Ru�B�J?�t�Y����'�&�N)m򈣕�J ;9d�#��7��`Ӣ)�9�|�:�����VQ	���F�F=p#T�g�I~��!�L�h"F BS���5L�H�"L�"��1G?������#:��1-�'�?~�eMQ�L3d㾷�d�B�!��J�0��A����J(T	!N����a�tYU�(�)��E�?�S��}�7���+GaJ��T¾�����B��v���#������L�ȣ/%>�c�3�P��6� :1&��%�M�V�1�UQ�Ʋ�"
���8��m]s�ࣆ,ڸ?���D"i�16�3�JOPnQ:�a��v��1��-.�_E	G�#��4g����jR�=a�m��8��i*��i�W�G��5frᐢ�ȭk_7��M�v0�������L�� �mg\9Ӫc���B"�U �`��=>N�Ír;�M����H�*֒)��T/�6�ÏP.�cirKO��m]��53&�?�^FS:B�������Z��b�	�{W�Oc��D8�Ь)#**��H���h3.��3��*DS�O�8����p���N*�A�7%�>��H��=�<v�W���zwƭCr�����'�>W�Tb+��O�[O'�/N|[���;j}}���u��\��\���U�۟�N,'�����G��C��'W���ڣU���SP79j�B�})�~2�ni�&X���:N�( -�Bp�������t���n�����&e�k�]�ŏ���~4�ѭ��NWѲ
9���kH��0�}��ō�wy��)������'����g���yztv��-8�׵`��>:�8� ��==����yU煉|m�����5Ҵ%�Ws[{-�����r6������|�
�=8~!ѩ#�( ��,5>&���Լt�m�/I;i����sR��cT�P=�E4��
m�h�� 1�5/>�8#�g�lt��Oϣ��J���t�=2k�I�J�-�B�g:���K���A���A(5`�C��}���7�����L�j��I�W�d!��N�cD��f�z�[퍫��_��W7>k�f><��/}�����ێC�n���V���=��"H�o���\�	�a�qJ֫��L��Y�q����R㧛�"�lT]TKz�)L?�ۜ�Rd�g9�8Bʴt��D��{�`���S���5J��~�����}����ݓ춭��L��f���7������s��YUI3[�*���el�h��eB�"~�%"�CST�Y!hF|#�N^��K�4n��;��KOM���j����d�Ⱥ�E`���P��('�� ��� A�I4��gRЬ�X"&ߢ*�I�N�8��־Q^crk(:LN��B��NSӢt�3��b�ү�h�f�fZuc�ĥ��1��XJ!)B�r��'��3��@)��B|���C�?��?�t�G͈8�\A���t��j�M�Dјv	MQLN�����W���}_EK�HY���Y��)�F�F-��S��9%�l-�������_��_�RދA	uu�*f�r9�ɂ�,�84q���ȟ��7���hZ/g�^S�J����*�p������+�Dv���AWB���t١�;i��M4���i]�ɶ�ue
'%T!#�1U�8�R�1j�G$�T�(|u	�JB���2�T���
�[��n!r���3�)��o��/��/:�ɐ�a��F>�4J�f�PrTg��zR��g�>��#�RT���pl��3� �Y�n��G�S�hYV
s]���q�}���T��m��L��[�5o,� \�i!}r��V�)�"���U]������V4�5 �"�s��B�.A���JD�a�G�Y�]�9��/ZU�sq������L�$�@Y�v�1��P��p�F�V۞��xQk������52��(���է��F%4lD�X�#������2�FxG���7S�Ӵ#��ޝ p6HS�rH���(Dh���E3�B9@|�D�A��T��L
(%�Z�݃�pc��YV]I11V]nY8���F�}!K�Z�gR�@Yt8^ct��~�Js6��h��)�X�U����"N; �� �3)9�����0��HQ"���G��
򀜊Rk��&kD�M�M#�nxck�b~��5�@�R}�[WR���_o~)e��,+�� 5VtR��XEx!�u��Bl�@��O��FH�v&@J,�*8�Q�pN�z3V��\T�����L��.����3d�l�6�Z�25������d@`�h3����:����!�i�7��J�S
rSxE)Ki�F`8_�qjՔB`+"���D ���T:���Ɨ��P�zp��I�An-�-��,0|�	����C�vsN��r���s^-�#��_�% U1F��Q.Q����PKEV	�k=�!��̔��J'cݞ��M����R��8�+�h[1=�4���F�h⥫;�w�ٔÒ��-r&�np�Z�WG�V^��H$b��od�FF9�#A fє�%����ϩ����)}
� P��
���fR&�R�B�O����g�z6΢��U,K��$��y���t:R�D�1+�o;>Z'[�v(ʦ�V��(Z�~��<\]&To��B����ʥm*b�!��唋 7B�g�E˥,��)�8�z�r��L�V������8��7Vw8���W��9�%�����Ռh/Rx4��G��M��l�!ـ�M���	�4���c��ޯ�P��L"�z�c:Ǻ\��FVKF���pL%z+G�{o���rD�{��N|=����!�l�U���,��j	�B15����B��o����Ao�f�1u2�����b��i�ɪ�XW5�va}/��myz�$\u|Y�ח���n�km�)>N����ѩ/�ݺ�����Ӈ�^��[���������ճ�+��<�}���}��������m�N���z�&�vJy�õ��3�f갺����Y���n,�Í3m�m�6���b�Q� �.�c�����*Q��tQ�~��*ὶ��C��ʫUg5��н����=����j��g�.�>���������� |��c����>�����Ǽn�^��L��"�(�ob[��wl]��,��cD��S`�8�������EK!��G��N�aڨ
�s~|�׉��e5�ԪD�8�p`#�|&:��۱v�45�3�(7��iuSZd�����ak��'�i���>����o��,��C�GvOx)4S����N�F���q�o���QN0~��v��P6%L�[l~`#�����B{2�u���;�ܫ��y��ᢘ���^]��Pӥ���䅗�f.E�G�c{��:ϟ_]\�_�/��Aw"'>��+��ot�ΫF�u�Q��������;��s�B�}��ۛ�=����>)���zh���f�ZfY~{�c�F���G����ˣ����q�D?�]�*w�Ԍ���T���7=qŧΈ�E+-�ՆW�PB�U�'�TϘ�V8mD>G�z)YQ��f�|����ԀR@�    IDAT����Um��*���m$Z���U� U���XxM�e����h��D��|:�qx8�8LѦ
>?�ʙ����q�
��k������0�T'|�2G�U��±G�C�2N�=��h�Q��I���9����_��C���Fv�����sG��184�DP�+��;�[!��)�ו�A%���U�i_�y��!�̷ide����7cjF!
�FY�=iᦩq�8B!>}�����?��O����k�#X_W~��r�t�����юي�;�3$P���TM���|&�[���a�LHu4α����j�r�V�f�9��VT�j5�2���O#f���H��Fm�q�y���/A���Ko-|&�r��J�V��g]��E��)�M`� R<=�'��L4�_j�?��Y������DFM�XcBE�4�¡qywV������!�4E1���w�FvD~��|d)�[�,}�*ĄS��tL�p�J���t\T�h>�)��r�*Ŕ~��3dv	�\4���+��ֆ�}��y�ҬIjh�#��{�J��o|��~����w����% �C���g�[D�����#�ه|���;p�Z�D%jҔ��ɷޮ ��*0����(��l�r�)�ɜvx6���д.KV���r��)�����C�!F�������K�DY@~�'�\�� d�#)��{��7&-}�Lі3��MV~%hF0N(�Z�9	�1�pX�E0E �oW=�&TVdS� 8��� b"�^�,H�ESh�)5��bQ��ƙP4�BFV�,|�p`>\�q4�o��E+����`,>"h_�Yr���X
�BE������%�Vsi��F����1���1`Ӣ|V�B�QZ�����m��( �L7���bQH)
� Ԍ)�N=��tE�>ۘPK(��������jEarn$(�,#P??H��	E.� �1�L�r�vIQ6��ʼ[2�4�j�)�8L�Z5�%q�@!
�(�`�R��aH��ߑ�CY�W�c���)���@N�B��RK?�q4E�
�1!,��.4�F\{��Gk�Hk�iQ��C���P.Kc���2��!pU8�MS�D �z�h:��7�4��!"1&'� ������
���Y�tA�Һ����Aԭ�ғ�P����J�DH�3~����t_W�Rp�*ZV��D��S.��i4��--��$h�b�C��åo��0c:��LYdN�1q�UIv+gw������G�VM�6lB�^���&�:��B@�	�V�h�����s�zh�I���a"�8��I�nQcL ��@F��B��}�$�!�!hF&�8ѐ��VS���j����h��U'|�����mt:�Fc+��k 88'}c�Ȧ[��|��+�Ȥ뭊po���д*�c�S%Nʢ��1#�8�)'ǡ'"ʯV!�
�b�1j�#Ի���u{��~��S�.�I���
=Ӈ"b�vqVC�!ˑ%7�qSZC�tF�Ze�r�O��PJ��c&R�c�"-ǈ0#�Yx-�k�!X2'�C׹C�͵��a��@��|�}��;���Q}���f]:�?��&��;������N�OmWţ��˫ӓ�M�G��>��w�]<���.�G����}�N.|F��v���&X�����ū��6���"��֥��>�&�g��ږ��h�M&�>�򍁍�Ïi%��h٨I��?���� �o�tb	��\��{ �݉?|��8Rv���^^?�zzux��!����?x�U/|V��&�K\O��ɋ���^&�$��T?Ze�Ic���؉�vaj���o:�d�����d�IQ~�D9,|F�~�%�O�*�!9#(��v{������42U���D�!q��g��B����C� ���r�1�&2H���|�����ES���A�R�;p�,$�ix�����ڃ���5m|���jTn2�ĔG�?]Q��v���6��S����;����x���֛c��)G��lnqwQ�����h^��gn_\���n|>|�������5�)��\>�~xz�ʼ/<��<>;�u�Dn�.n�֘>]�����ᥗ�h��=a7��|�M7��O����������w��ݖ��h#�*>e
��F|���ٟ��у��8�0K�K�}�>����'�����t�Z�,�|��O~��F�}N��^��׿�H���1��vk�/SI���^�Д����%��� Q!:qh#pj�#��жeV΄<>�(��J}8C+E��!}�B�����𶻢9/eU]�X�|�q��솨bȪŏ/J����U>�N��8ʹ�S3�4v��&�����\��T1e�!��J�r*�8�3����,�[ ��~>0���+T�II\Tۚ��_���B��
���'��u."������3eT8(�h�;��(����8R,�.�r>�%�K�I����r)��m�t!~�Q�L�h�#ʮAV���_��_���ۚ�'(݅I�.�^��F�B���%5�B6�K��z�N-�IQ#\�i�OV��h�����֏���쉨��x�ې*�C�e�̢_���
�Σ)$�_�f]�+ݶ(|8~�p��Lc͉A9�%��(k�R%:[���F���iO���E�[�9O~���Fvj��9c?W�9"k~mOc[˷C�U�	�H�r|zؙ@J-{�%�tS�#[�(>�N�B��)B4�u�a�%
J�8��<��aO��h���9DHI�/���"�?�Bd#�4K��H�\RsPH�����3Ы@nk���,�n�(AE��h����×�`�׿����\g��#h�.2�����@��B=ה�J�+W�Y��|:h��Z�
�P'�'�a����`���N-#dNZ�ZEuҒM�A�/�"��AZ5�k!���~���bh��+9eH�Fk�0)ӏi�DC���d��L��M��1�B�4ܒ��FU����JcYqFs�( ��Ñ�w����P/����!�f�\Y|����;pS8��S
�B9�Z2�PH-�ql��
&+���z0�������=��k��OJJL�*�g�4g�&1�X��Y}xY�Z��;8A�^2�	�t�`-	�}��K�LM�eH�@V���2q�I����
�A�΁D��b��G�����o,%�ȐjÍ��M�*SYr�<뼬�JT'Ȳ���4�v8,����L���arpR����n�k2�QH��r�e|L�}��B�Å�ْ���ƯUHN��RJ�\����ꄦi���P��Kr
���|��98եϟP�GǔE�a�����h�ÉLt�������Q`�ɭ"\VU���F)�8,����z�	-�m���r���&$����85|c=�1V��ӄp��|�8��N�w��XLN1�[cQ��B����q��>������8��K3$�I�$�4~+JS�$�é!2�t�p�������F��*jJgl�Ԁq8�0��pN�|����!i��2��[R�b$�'�*Ǚ�/�6Q�&7�4�)������8���5V.r�[׷?�pH��g��%Jsjդ1�q���f�m�i���e��sF3~�M[H���\�X]`�4P����=HMi�\>�ޔ�p�63_3팱�o��$"C�a���Z����@0e�ִ5M��A��� �l��6L�7/�L�N"g�)�rn������^�z�$D�o2MsF8��YB��7�Rn'KA��Gb����|�~�G�Ís����ѩVu�Tt?�42���[���(�=�jQ�	�C|+��h�q�=�~�f ���<�ۦ.e빧�mOC}>�7��\�O�z��fWc��ڙc_-{}upq����gO��f;OO|��}�������h���NtU��!G� �ֽ3�K���՚������"54`ӭ��*뗟9.���ޞ�$��+��Q o��lq3a����X�ٟ�-�HyU��~\���x}!���������ym�:q����y���78���3�]_k�F��󛳓\�V���
�Y/ks��0%��o�h	���������?�W�r|��m��U�G "
�X&�#�1}I0�zMH�L�1��hjv'�-q�� ��������O_�GgO&R�&dj�qB�93�($Y�-�!�2� o�,Z�_*$:|����1�Ek�Z��m16��CLEˍ�����(+N
� �_��»��v:m�,�c�$���dq�������gO�Y\�%�������7�����'��o}����8��]�s\��}�g��7&����^�J8i��]m����������ȍ�����o�t��3�i�ބd�p��.���r�8En��qhz+1Y�\�FS�#�-�g.k����*�n� ��ݕS�n��+�ϩ��U�k�	�t�κ�rTŤ��k)9B��E3�*��w�&XV���gtج�T���S	}�dA�������\Rh�����EK��B��C�/]���b��*������d�iU���Ñk/�č@�6�6V��Z�,9�J�X
���8�!�!�J�t���DB�9ҁ��8�J�/���@8�њP�IGk-�Rn4c��vLKNN)~��Q���y����7�I���:I<�1:��ii�JPh����¡�a�ᐒ"W��Z��ÿ��@8��]��΍|�B��	��!իϊd=z�����U��~e�{yKqs!�:�v�+�z�~-͵�SoE6A�r�+�+� �NC:o1MU�*������6؆�	a�� D\+���=l��h��H�jv2[!�F�"�*p�|��C���֞wY���C]�LKfm��j!s3��H��R��m����웵��$}Q@�(c;)�8YKv,ٶ�( k]�9F�q�\�������R|��8�@��RHi|+u�@d��!��E5�t�K��MvNz��l�'y
UB�����g�U`���V��A�jϘ�T�t:ȚGֹ�(ĀF)B���Q����(����`���0���SW	��D���Rp4@P'^������~������e����<�6��,��¶Ե�u5�YЈ��/_c~���) &�H��^2��IΈT�c�g�2�>��:��պޞ�hF��t|N�9Õ�9�l��'[F
��O!��R���\H���/%��L�L���IY�, ��@J���X�����Z8'cSkQFFD�a_n��2�P�W��`dS�U�/�wb���i=�Ώfʷީ�Zx��R��g�$�r��	io�h&��V!R����)��K��l,�*��,��:�X{���L# ���!F`ˡб����a��L����12"B�8��IY�;B~����#&?�)%~`m;(��@
�"[/�)��6�ӆ�p��f
�Bc�*�@���8;Y���T�匟r:|��9D"U	D.�|&��Ț�8{��!�l�J4M�8�	��e���F�b:x�Br��^8f G�rr��02����O"�2d �ic)���O!Ȧz�j�k��"3e� ��_�U7�|dc�F���l�\&!~���2`�"��;�wň)W�C��K�� �Z@$�I���z� ��(?ˏ_zxu�1+Q3�p%R�@Ҍbl�����L�@~��du1���^d=��8ӢI�J���'r�4�GAn��h�F�5��������mJ�B`S=�Q��@L���Q���6c!#Ę��	�h%��ut����8kt�2��h�x��M�����u#7ʵ-irԅ0u���!6���i�J@j{�CH��S6�B$v�G\?	ƁӔ�Z�|є��F>�3+w�956jڀD3�F���������@Yc�J7���-��B�Fj𽦩�hY
3r$���S�cZ]NUL岽H�B���8�Id�9Ղ��ƺ��X�c�.�����D�sP�g����S�E��s��k��~[LG��F8���c�2����T��-�Q�CVbk�iD��b�('K�ȆƯ[��H�C!�Î|���?ن��%y6ysx}��f�>�N�ӽO���kb���6¦Jm{ ��:�\=:�ק�Fg*�߫$�7��l;=�wp�n;��G77Ϟ>~v�³���#��t[�U�c�����.u)�\�G>��j�z�	�6�%{��őekiwo ����o���_�h�M�7���4u:u,��Y��|��^�� JD��1�F��������]� ]9�7G�玷MpP|=���'/�?:����>v�_}���n���Ο?�w�n�171��7'�7��|ʦ�t�8�eUχ�s@Sf�3"���G����2�hG!��#RT+�6�TS��ڥM?ZіF
Ȁ8���9�S�� E�#(-1_��qW8tL��t_"�qr��j�Wnds�K'��}i�P�>��&�Yї��YՒ�R?)ǆ0�B�����.?+�(G��Ӏi�:�G� =�)�N��L.��Ċ�V��/7���6��50��,�4�e>g��&�ق�q�������V��������o�w��mo�L/������w߸&@]����ڊ�'&�P��V�;`d�`:�v7��Q���U��?�x���~��7�x�%HWS�^:q�DB�\Q�P�D GuY������a��߫&���r�K�����v���}�`��g��}LӽG=��}$c�HI@3���ڊ����ԇFM�I��V�c�������'��������8�9ȢB�&!���L��w8Y,�U�맔���5��dȦ�j�"^
��K�/ԍ�\�vغJ4�)p(�)�_Mo�1H=�T"B��zM�L�����hJ���
�R�7���Ѭ+�)M.��9B��R�Q9x)�DFg��a�0�݋����>�\�]Ճ/H-�83�)��t��ZWۢ�V[ ����L���e8�s���C���q��U�ь�`��/��_�@GW��Ŷ(�'.kՌD�x�iψLGHb��pH	4Q#_�z��j�{��֛ig))GfE���i�%��xk�$����>���g�g~�G�)������P���k[��=������_�!�B�z�i�6L	�_"~+���!
T��^��jS[��l�f� �t7�eQ5Ɓ�,ʨ�pD�/[w�cY~Uy<3"2��'x0��L!��d�'�oyB�	@b ۙ6�[�ncW�؟s���Y��j��������;Í{nވ�,��:��0չ�k�������e=T��dA�����$�U�:"�#HѰ*�:,ѵֹ�)u�O��:ѡ�@�t��V�i�e���|�Oߠ�iH��zI�4!�R���O�����P�z}����^ȥ[����oO,��ģ�s����6�Q94�ʹ$)Hw���{Y.I�����-�mQ�!�h4�����]��յ�'���[��hF�_�r�U4%bh��p�M1mqRN��8qR���������;7�E3�������'��Es8��T9B�8��5Ҕ�E08q84�ɖ�� �D[i~��đ������U�T4��q���k�>e䪣5e�E'��i�$Q�Z��C��|��FD!6�\S��S�� ��R�r�YCV��cF0�C�6�fQv�قISn�����i��]t�8@�8����5D-�E��M�����ß�_Q ?kT�
� �^K���^�R�**р��� :2�����`4� �ȅ�	U��k""ė�*��꜏p�+zuڱR����YC(��Em��ϼ�$�B�|Y����P��m��_eE�JtR�-0r�6�H�p#f�1�����Z2�-�f�M�z�b�J7-Krmc!�����ku �J�%
mu�)�)�a*=$���6m'k�l�@�U��r���8"@N�H�7e������ds��R��I���]'�����G�����HRrk5~��?[�6L1ˊ�Ǥf�ZR�#s�U:ي��U�2G��O�U��v��S�4�ݸ8���_�BpH
�B���K/�N� l��6]�p���D�p8@N�ZCVz��#%�o\���[�����_e�J�H��p��W(j%���T�QX�pLv;�xU$:���]u���5\b��1.�    IDATÿ.*���gޑ�C|kԭt�u��P�+�)�fD[Bt��b"���>��Lj� �_"eѫM
9A�ڀ��5���Ǒe���S��{�rP���ɯ=���Nh�DV��~����&q)4�6�)�ͩz�>Mk��SN`)BE����]�{�|��
ot�ɩa��V��y�BA3��������LM(RrM��7�r�C�e�K�g�8e�8:��D�qμ�l�YL�Hk
��f�F�k/B饠�ұgT�&X
�u��߄����[z�ON.;��j�n;ob�{n������>�
�����Ly���ǔ>}u<��hWo׿����8����[J>:}�g���IG��IЧ�>���74GP۝�V�c�ތ;I�yplK;����Q�B{�Ƒ�=�߹�o���r�HUB
QS<�y���ja:o�"8'���٧'BނIT�;r4S��b��q��Jzw�5�s7l�y��g2_�����CSD�x*���с�	6����|k�Uo�|N~�p�\v>��1��E���{򘜩��vc�6�.���W[�B�ڮ
�uZ��cB�'.��7�m�8�	�g�#�bjE��Α��!�QB���-�)4��J�??Z�m�ԲWpH�����xO�J�G�*1Ro�������B�`D�֔$�Jp�%�N���ɏ �OpS�g�kU"@�G�������R~��ŋ��7�(�y||v�f�Wn;���v�+�~!�[�/����z�U,
~��5����y��S�^���~�7~�~��n��v�����X���E��J�u/25�����r� �'���8|R�3�r�s�uG2Օ��A����̿�ۿ���,-M�����y�LM����<����M�J��H`[6��V�E�T+98�#ڪ�k��א��d� �g*��B�ئ��ȓm;��9U�a	�D.�&!�O0�PR@�є�S9�;*��.D��aZ��J���ᕰF��W��E�}�GF�b1;��tX��������
���mD0d�{ȝ��G��TQ>n�@QӺ�ČSuM)�9G��{�)ZJ`���@#$'K')�05u�ī�ጷ���I�`�L�1]Kd!������;u���ΑG�(����,|��K�L#�
je��uہk�Zt�1���Q�#�|?|�q�?Lг��^? vq��_}k�i�V�>n�:G�ot��>5wj8FYp�q��`E�!�U|4CXQ|�(���OA����9h��p �����3��[oh�����DQ���c�M9��l�xks�W�\|�z�jY�����X��uWդ�iYI��؎,��C�dG�c���bB��8c��Q��IepʩqL�����(�:�O�!�jع�Eˇy
�*��	��A:�j�sP�h�lw�J���4�~�5Q��=��������C��S`�d4����8B��PB����i��:׀�rԬ�~M�J����J�����৏�N�>x���c��u�\�pj~�/��9�,2��@$��c1og-Mi����8p�P;����fei���3,+rj���
m9�h��|��7���#Y�� ���a��N`[��OG��D��)  �~j�A��T�݃��9��8?pL��B������0⫢y�!t�>
������+1e�%�TzKK���9)D��7�q��Zm��6�㘞���������)d#/7���О�m��@���S�N�X!���� ��������<�!}#��BU��s�M���'.�Z8��%����X�R�r���[z4~B��7�$��N
��q��^##p�*����"�x!4C�D�94�^�,��AF(������sⷙ1!��i�;@��U��qR+��"̶o��Z��Hu�Ak!�[Q��6�
]���4!�+=}�TȠ30D���Ωtg~��e%�ρ'b�H

�8�\�Y��Y��5�"�3�~��F��t��DHj�&%jh���C�h�ɯ�iHE�5��d��-�x"B"sL[H�hjhMY|�ե��p��C3����#c���k��N���V:��4��
Ͷ�j�锈�m
���^�ڨ�h7d�!7~����I��P^.~䘥�ȯ!��Y)e�l��f[N��LV`�&5�rр�F>e�R8���Y!�{+�4����4���<g�u���V��7�tQVh>B���f�@c�:��L�+T�u�t4[3��&^����O�T-��T�������ZVY��[/�V4�o:�d[�eVi:�M!����J�������3�m�\�����*�к\�@�ƎL')!8ªX���-?�5�� Yb:#�K��}���┈��U��Y��m�)��|���ěYh-?>�I�D�8�F���"�y��.}Y��<5�Y��!��V|v|���)S�L���0>�b�!�W�l!��t4ӝ����Ӭ�|֘B���М?��M*.�'�����ۇ��9W|��i����x^!~�^�(����Ѧo�<z��͍_>뻛��������lwO>|r�ć�~{��>���}��O|��w����7~�B�n}���S�A7w�x�.�u[�%x��$�u�M���E_Ȭ%C�|���B�ϖ�`*ȶi@b*�\YN*o���!�h�=���]����t(;���AHi�٫�,�V�EU��Q�才{����O_������_�=�`���w��!�x�C��%�R�^��׀��jl0��J�)�o�9e�1�ү`��8B�C݋r�ĵ
/�m��?)�E*�NN����H�4��JJ��1�J�K\���`8������A#���R����#�&����4�9E7�H!hHɦ�?Nc�#�)��$���*���^���RFfә�Eִ�)� ��x��H6� �B�R�)t�� j	J4��f�.�f%�QvU���c�~���G��v�/_�<���K�s�7o_~v�#9��8�������o������>��裏T��w��<w���'�|�L�������>Y0�y��n�>�B^�-��ƀ!���B�$�v����!Y�J��n���h��׹�Ǉ�h��/^�0��uy��Y.A��_��W�={�΋�ѯ�􀘜��xW�֖��6Q=��:���f�9)|d��M�,ޠ�"4��K�m
�T�C-%L%6��	\��!r_��r��� �aHMV�/D��iZ9%L��C�P����)�ǳo��!�45��h W�c��-�ID�Sc,�%�I9�-��(�_c)���trؤ�q�ݴ��U1��"U]�>��,�4q���T�5��:Re'�}���v����o|��'9Bg�e����1���3\��5�/*�\��9u"Zc}�����&�.Mj�!u.1��^%��|�-Z��O�2�ϟ?��?�������u|��*.^���3S'	��v������o�Z�����sÎ?
ђ�,��U��qn]�e)ц���}�Nڶ"W��������w���M�P�!� X5��*r4 �r8�Fg��D|�߽�����}����,��!��Z�Ȧ��5����m{��'.E�%;!e����z��od�l��U��p"��͘R�v�]^�5�A�^�|�iϝ��q��H�t諕,D�tzٰ9ԜT��+�6����ҏ�aC4C���Ն(_��*�u--Ai>G��cZ�R
�|���h���!������m;ж�Pc��m���o�UԵ]��|�/��%��ٺ�m!b��A�S��吥���h뼉����4� �(P �+��X�a���ΦL�HqH��]��PD���I�c��B||���)K�[���v�i��V��hg������?���U�4Q�S�8�9��FM��Z�p��cʁDK���P'�-W]xH���K��И�C��w|mQY��I��l��DӁ#���I����xU��3��R�\��Ԫņې�r4��O���,q���$�!��4���:s��8�,&[nj�[)�Pw\6g��)$[��)���S����4C���c��,�*2�uHMo�l����� ��U| �,��,S�(�(7�M� ��iZ"��~W���|7���X� �L!��E��֥dZQ:��\.N���bgZU��Û����	r�.N��)��C�������?��w����,!]��a�0?��8�@hEW�4[�i�ݛx��B�m/�A��,4���W�ϩ����!�����WD�X�i�c!�>BP���Z�@00ס�i#�dZZ��6BH[tH��C\T"AN���7E��KǶ���M�3�������(pZ�(���������s"w��b6�D ��^��J��.:�Es��s
���lQ֨hd6��vз��B�VYS:j����I���Jt,����Q�m�bJ�_
k��#��)�c �M����|���U�X��p�+�o�!�m�d�6ҏ< S@��?�6P�iY��ƪ�ĩ���aD���劲�e�G0r�Ք_	j�qj)�֒�rd�DBX�겫¡�)?����NE��ڨV������K�� �����ڨ�e]�t��*�[E���J�}��#T#�V'�/JA9�����Gw|k$�&`B�,���J���wv�����'��7MJ�"*$�f�@�_�a�78��!�s(s�?���Nh�Y�i�F>\z6~S�j��#Jِoo�bK�����#��~	��=�v��m�˗�����/��"�okR���w�}
)��ݫǯo��n�޾����|�����[-N�Ƿ�n^��Ӑ~A�Gw�o�����GwO���|���E��ִ��>�gO}k�1�m[B7
4uȼ[�oN9�zG�m9t�[�}���#g��Á�ė�
}��B��gq��+Oz��a�'��|����@C���4M�m�)5ky�����cH'y�YTo�;-%B���/����*�I�E�R���z����e �!em����,�A=G ��Ub��)
��1,�8B�,���r~;Ė�hYB�)�QfM���~ͅ���"(�4-=�р�֒���O!�����q�S�M�MYMV�ЪK��!ɪ��x;�	!U�!%j-��M9�FQ�hW�u-�!#�V����|E��R�_����y���9�Jȭ"r�b
q���p֐��v��_�gn�En���n�t��)E޸���Ɵyv���k��[����_Y{Ȏ�m|��Y!�k_	S�w?�r�K	w�O}KK��~.��&[��wZ
��H1�ek�C����K�G�Q$2ċx-M�����|�ه_Kמ���t7s���տ ��㏥�?����WF�r�"���G:D��D�g�Ǉ��ء���wRR�� ��pZ�rI�t�*�ҷڪ�
�9�M��	����rO�qIpX:њ�I�;�"�B�ZG!����e��4S�:�#d��|����m�����($�P4�D�̯%�5éQ�>!���(\���,�7�Á�9
��VV>r=sޓ��8E�*B;Fl���`��[W�)�@VKͧ.4�gl>LЇ��K@��w������&�BPK�9K#�)4��Uעj�V-���윣�KT�ԲpjDL�	�^w�!h��wT�ׯ�RXU�`�n+��vO
Ĵ\��G�#W!��V�"ʇ�����ϡ4�@nE|��@��Hװ�,[�a7Yk�p���\Ӈ
�%fY��r��o���_�:�ф������OEԭP��!�Ъ�,��c��
�U9�%aeYNUS8k?��k�5�9�=�a�$Z�U|���Fp�d9�����1'��ɤ� �m�Vu%�5�o��!;��(���1�9�����d�I�RT��X�W���&;�m���)�C�8v���A�U�J	RӃ�6��吒E�Phg���Xu�?�:a�V�U+��7%�b�RT�oG��k�����*j
7 R����h�p4�Du}	�D뭅L}�)G��6���� C�p�����v!�,V�V�!"j�UǷ�ja�b��Z̈́���(���
��\�6JT�r��@�'�Ɓ��F"e'�Q:"�3�UQ�/���뤊B�FMJ^Mɪ~����Q��@Y�v�L�L��)%��a��he���_��NL��wXjF��sj�o�N��k��tH��`�T���� !�-�S��F����r-G&�ށ�G�.'�I5E����Rڊ�,��NrB��	䘆���@U ���t���ߧ��¢���J�4�f�+QbG.�*�i�9U�)ʶ�M�R�-�\��562�K�#������`�ʯØ�j��ԧ�J�X��Qbʦ�~�ρ���r��j>�`��&�B�۝'mT���NSJ;�iP��rMW%fSd�u�U-�U��p�ﷺ��cPhɬ��d�ES��2�C��/߈�|Q�F��W�g�:�u[(�NT������\V��h��Z:�)���Q�\���K�����B�-Ȇ#�I�I�B�bj�5�{����,Nʉ�V7�ߐ+�W��v7C�K�����ڨm�.�t�1�Q Z�*�t��B��'����e���&����j�@����(�N�ʙR0�d����\kI)=A��K���dq���@�4#P�U���V�R�'�B��gLj�i^� K�2��TTb��J�Vb!�Rp�	�W:�JB��7���45"sJw��ؖ��:9�*�����4��S,`��Y��_������)��<�V$�XiRU����;��r4W�#�J�T++k�)���2�)�qR��P�V��8��"pڴ��9�-�ܢ:Ip48�q���U�v�@ZE��m��'��\�ׄz��8��1!�@�ad!���ڃd��-g`G
�<eYW5�ZJ4"O�D��!�A�% �&U'U��C 7H��8�ģ^�N6v^���~l?W�M��ǲ����g3o^Ͽ�髜Ň�7�}2�x狝�:��n��p����߱x���~��'�c�w������;B������W��W=_����W����~������Kп𞴷̶�y?�s�mE�:�?�jGӴ����j�$�BU�������҃���v|�����R��4�#>�gB�u�ӏ,���r�j�(��)���Vx�}�<��FV���Btգ-�!]����|�P��p,�<D9R��q:�'|N!���Ip4R�N'���%��Ț�6B)�G�y���dm#k�-���2�Hʊ���V���i��9Dd!�rX
�BF�"��7>M�DQ�_"N!��e5UX�B���i�T`�K�@
͇�$N:��i����60�ҩ� \�ѦV(<[:A�Ѯ���拎�I�݆�)���K����<��#C�:�:�p�[�˜���:|���p~S��=:��y�m��Y�.�Z����V�Of�� =�s����˚�������G�eP�z���2H銸�X"]���15oJ�YbO��DФ(���1>��8�����ZS71k�D]��-�G�������'��������瞳KVϞ���H�J�Ⱥ�QF�}ā�r"j�,o�B�9F�2�cw�:���*�6�	����D�Nbh�G�𪤜�(bD ��i�#ѴӅo���U%B{Ruӧ鰡	)��q���켗+��n`]�gU,R��!#�c-|�D��Ḓ���
�������I9Nw!�z�����U*W"���@6&'YS�| 2[WB�'�N~���84��/��%��Sp��b�]3>�H\��W�T��r�?��?���/��E~,���>��:�Y��4LY�ƖI<�3����ȥf���h����}.�
������l-.U=�x���h	�����G���Qž���w��ڃ�2E@#�76A�F�M0� �DE�z��֧���vOi��*���L�ŋ~z���2����Y2�8>��P'p~�)��pH�Ouڠ�=;�`9�X���ϺB3 r��th�N���ݒ������f��ԡtԞ={fiVm�
�����+G�l���P�sΉ�/�#Ǳ���t�B�    IDATԒ��>�����i)�h��T(75� ��pL�
N�ڔo�5V
k�����~��jdK���k[�c�(kX.�*V�(��H�E��Z20��v�3����_0�Z�mǋ�����	�D�����y��]-K֞~D� BPn�+��H�z	�j�nm��Dj@�G����#�Zz�� 'ES9���r�D;	e	��)�ҁ˅�|D9���H���f�7_Q?X8R8��� mt°ZHRk@z
����K����z^�8�Q�ܲ���5���KJl$�'.d���iH�rʕ�8ǔȞ��O�4�-ć��ZG��T�t�=��+��H����b���$U:�˗"TV>ܮ�j���sj�,�(��z(�4�O9y!|b�F����߅ �ØrD�|ќ�ni����D����D�բ`*�,�6��t*��Ʀ 4U"��p�&���9N<8�I<�g��5�E(�������_n������ϩ�4[���[�PK�4Ja���@��U �%KԐR�%�9�D#�[2Z`L8GKr����q@kA�f:J'�r�9�)��ZiC�r�k"_4$+�5�~��4�·h4q���  �'N
G�Bhp��u��-%��1#B�SJ�KA�|�%.$xf�����l%�u[�nM[8��f�1�"$EgRh���VN�'�hcñ h`j ��!�K�re�1��!Y���J�&��cF�C�[�R �Z;��a!�.Q~����!����4V��O"|����&BpSdcYמ%B8j�q�+��d���~Z�i�gޱ�:��.|8f���DN�aJ�#�į���Z��p��h�9pL9t�JW7�PS���s���#Jh���#L?��h�8���P�l$MnQ��\�\Q!)���2'������D!FULeE1͑_�*��2��d�5î��%毊i
�!|U:��0�ó8�^�1��l���(-}��s��v����Y��zUn�#����9��88!��-�rE�B�³�㷐�q�-�Y�q������aoI�WE���~���'����%H��:��"�2kP�r�鐭IH~�Йtb�XW;�u���� �M�|cU���恜Jp�gMk�E��BYq:��5`W+a�P���T���E�]��~��W�_���8��$�?����J�7b>�������!�+��_�<�2����?����z������u޾y������On?����xZp���;o^���6}.��K�����1?9Kh�-�Vk�NZ��>S�N���.r{%��g�![����AZ��c���,��z�����go��~�w�w=6����Lᣏ>�x��	�^�C�r��x$�1B��m�V�E���K�7��_��sH���Ѓ��n����<M�6�j��	��P�tB-'��[i̚�`��S��_���蔧3r!��!����V��_]H)��,b**1�%&"ڊ���5���K@�=���:"5���$�8�3��#	�V�-Wt���}QV����O'p�B�	���dE��$��MC�aR�.�ԮE��|EM�8�X#�k	���WrY!���F���\Wlϡ�_W|:��������N)|A��4�{d�k�TJ�3���:C���4�"ͥ!W�rv��dCs�z���J���������s��>���^@��ԃ*�����:Ӑ�J�=N7OU��l��GK�TbR��-��Bd�����Ź���_��'�~��\w<�v'�g�����wS>���֏TZ�/����^�0٦��w����g��Gf�~
I<��F�T�%1�;���ښ���n����)�}�d��W�Mo�VA*8�����ـ+A��qd�B�*x���%�p���d���Q U	�D6;o	��@���p����I�`ʩ\�ϲ?����Hui5�A(Z�YqL~65~�eE�%�\}��P��iӬYV�t�w�'Զ[�*j�ʂ�E�~�����v�۹��ԣ9i]0.�~Ԡ��o~��	�]<���Bj�\N�~t���1�M]�;�r��j�^ GWh�(�7&�淾�-'@�ub�,Au}�Զ[�d��j�>�y��)�KHa�TT��2u~b"PK��e���31��� 7�Oӝ��,C��0�,�c����qW]-����(Y�l�!d�P�W1�7:[r*�i�r�ahC!�,�~��E�  �B��N>k#d���ٟ�x�I[�.�Y�R�UL���x���U���t�V�J4�X�q��!��uQ0�a*��!�f�N�|��;��\�Î� ��nY~;#�2k�����K��z���1�)
�g��j�r�������nH��L:9tp�-�=��g�_��_u]�`Rۮn�VQ�YSo ��� M�j�D���]�r�ur��U��;�E��t�5T���60]�R�%��[L����)`vdM��,Ĵ�D���@�@L9�M�j���Ee�IlH�$�W.\E��u\��8�);.����=Q�Ԧ��r[��6��@V�Q��H1��ޤBt���־\ BQ�_)#�2�\��%���M�NNSJ=Ё��h[Z`�WȴrlY���4�,�~ ����qX#>'�B,�~;ܜe�+J-�q��������C��95~�����{�DDm�h�����R�-$B(�5Z���R�['���p%�m�f�/T�C���Y�(�C�����V$\9d�l��#�Kt�R�9F
G{B|d��>~ͯ
�P���D�W[��ꍃ0��B6)Lu�-��_�8��L$�-ˑ�tZ 
�|��u?�!0)S�L1��tR�[~ �c��v�8�=t�<-�T����"\9�"'X��wi�����C�᪑��t,$f�(0q)�0N+Ť�y���||��N�-?~
#�VB�r�R�#���b���D���|�5S��EM��`��rM#�F�>�Z��PEY[T������ܥ�P.)�rA��*ǩ�i-���(s.�t>�(��"'���XzL����
��=�4�=dH]�^RpD
��`�E�a�D�5ƩOQ�TtY�+4��� �O�=�O�%���`)
�P��:a�	��
���C����b
G>T΃Nٴ~³U�Ɂ�X-���M�`4~���-W����LS�uq�u�T��c�f�p"/ԩ?�qd��<�4#�F�`|�z� �2�1����
)�C�t�%#�C_�o!ܨ%![�>Y~#2��I���q i�Q�֖vPL��_æ��hF������ �W�|�@Ʃ�i��J?<	qHUH(}��_:�ҏ	�I�ͩ��U�tXQ֐�7Z��?uK�*xf��8���z��3!o���W��.����ڮ}r:It���Y��V�fꖲ����\��.D���h��&R�,���2��8���
�Y5�j�����P�c{�4�ɒ_${|�x�yK\�I~�ݷ�vA�J=��}���m�8���ܾ��ΧSw�[yl�ݍo|�ү�}%�|��-��7����n�S����~p���������ߓa>��Gw:�y|盛nO����q+�f��~��~��ڳoՏ�G��<��|��-� q.�B�NH�D�-E�{;��&�H���1=@ �R?�3?����o�Ѽ��２���(��)MG͓����@
�0�W~ųM7�����'=.��KWN!��b�*h�6� [���̇S��9����eq�,QV��6��P%GJ"��#d;F	f���Yn�JL3\ݲ�I��E-5�hs0��pX8�B��s�j��U��Ŗ�R�+Ӫ!���LM�xOj���U�JPh����K�X
[W�1�	�����ve�0'�B��䏐�>�՘iN�Y[�ܵ�*�b�F����A��h���� R�! � ���tu{Qs������V��I�!�w���t{�/*�r�bt+s����a	*'�iE���W�h���Q��:�i��B!��r��@���(��|��gϞy�K�-�]��h��Sԟ��d�W���[Or
X�G��F��PfO(�E�� �E���X�Pݴ~�.�T����8�o(��(�^�(Ũz>�ն����j�?D�t�r@���&��h�YϬaj ��!7���J�x!�'�ռƖΑ"�����,QYhiv&9;�[i�t�PH�-Bp����:�5� �����4�B��e��ǟȑvrʍ�(�Q�t���ibK{�no;g�m��>��t�8�������~���2t��4���;���K����������1�����&Ԣ8��95\�cd`J��B|�@�ź�����ŋJ�ҿ6�W�Ǵڐ%��u��1e!�ĉ�rl�N�q/��E� �,�r�dKm��Z���q�VG���)(��E!z����lm�Ә5�RG�r�h�oI8��'O��-�Ł(D�,KD5���P�,})w������9|��L�9%��[k��n�C����|�����Y�H�9�������?@���J�k����>����.R�8B�;1�h�G	�zc�@8hȲT��Z�`�U�/�8CJ�f	����r��$�%��m�O
����٫��jI��:A&������N�Ƣ�k	G��`��gӎ������#��m�����Y�����t���h����r��:��R��ں6Y���NHA0��z��q�i�,Y�d�,m�֧����U���<O��LY���M���tn`�"ȥ �1� p,� ���5�K����)K�{e����@���U���P^�C.B>kh��C!�(~4xY�DVJ!N��B�L�v�O����)��t����"���L�ɚb���)�b���N~m������]����4e�H�7NUL����_q�G�g��h����h�V%q��1=��B�
��E6���7�.k�h~4̪����ڀ����J4eM�>ڦUW�/���U����*r��
U��1�ue�,�Z�[xH�W%ԥ#D��L^9v��̊��ȑ(j�+�6��p�f�M����
�s��E�z��ö�!�cv ����\NY�QH��B�ս*c^�MG�
u:�"m�)�#
1J�^q��dKa�L�G�9����Z5ev�S!K�T)iE�
	a�hp�Bv̜�xO�N����WD����B6�C�!؁ �[�P�J�!>IP���n���B�q8��P�ϖȊr�[�r���k�U��d9n\��-���5�Pc.̈́C8�Ƨ` H�Y"Ax)�-%��DCHb�|u6M�Zp>�O�>�i�Y�(�&ĉV����$�#T�Y
UO��-�S-���JI�P>��8��q4��(!�*+d$(�>r`�����_Q�F!YF",_�z��[�)4)S���ē� B�(�[�zc���ٮ��8�Ŕ'�vooZ�E�B5�ү`�1E��������@�SQLրW����5�_�Ș��/�q���4�_8�WXW��5�,>�hU�����W"�"����iO0k�ު� �V�>�J�v)MES���H�7�P��#X��#�<��u�`?�z^��t�Fd�05dy����㝻󓸷3��J��ZGc9ME9�iXV�P8��,GZ�|H%8�h4�h��l�ۢ�A.����FP.$[��b��K��t��=��ڧ��w/@)��yE��C��]����D���&�{���f�w�/�؇���}�W/�������c'o�����4�Z���o{W���/_��ɍ��Go|�雞���}�����鋢��?
��Z�ZN���R�v͓�"X���8�Y� ���5<�>B�-�7���<�j�?�NN���`��~��~��Y3�χB��O��y��[��8�ꐈ�Д�~<[P��'*)Y�xWԓ1O<70������M�R����=. N͒IɭU�yx%��B�q����-m�f��m�h��#�=N4VzR|��W�Jı��i{�ib�q&h*�R6-�f��ɇO�C����ٜ���T�-���*��&�TVkLaj@~%�DkZ��$�5=4���%;?�))�x\M�q�S3L��L�t� � ���/�x��
D3F�>�#%'��΢�e�s�\���Yt���"��6Mm>B|Vc�sbD�kM���1r.8�8hS����A����2��@������{�,t���_��:j�Ήt���R�v"��ȽB-�g��K3���щ��tK�_3�5 p=�g|�%Z,N��X#��Z5�5[���6�����ׄD=~tg��裏|��~���&m��BO
��#G}�Mm�
��D1VF��-��h�"��=������/�q¤��!z�0Yj� ����I-n�^
�t�EM�J� )#h	�=�~>n�"��e$��x�h-��. (��O% lë�6���϶o-_!
|Ci>��g�E�:9p� cr�A��m��8E�ަq�-��a	v�闸��.�&����*��d)� !�bP�%�L��t<�����~�Sŏ60}W>G"r��4�H[i��"pB�9l+�i��ń�g!��k͙���?�(�i&��.@�|�Kаp�Ĥ	4p���\�R�$A��USJ}���QW~j���"�s�>�b�5�B��q��{�gSG-�zhYw[?�uuDkH75賘�9-!?�ڃHTBu���!)z�����GVݏ�/�_뜱�6�?
�	��bv��C'A���^Q����u :R�BP|�#��vLW4O��[Q�=�,A.}��%�DS�h
�A��RJ���S��Y���4OBP��P�J�p����WG�2B��>cꖲ�ڦ�=b���\�Bp�N���j�&&q)�z��~+�(A�cD��h�#� "@(i���ï���{e�b�4�I�w���֫�N 8G'�6Aۚ1��Jq��I�	r��f]e�Z����<��ń�ռ]r4[�r�� 4&1����.�|?�����!�v���-N\�=q���\��z�ƹ�� 
�(5��A�_J������|d!��,���|��8r��&d���i�4�����S�U(0B!R��9�h
�D�X{B����x��R��g!= Yj�ax:��
��vh\�N>B˔��Gzշ:�N�đ�h�"_
�C-�5��©� �8g��#��Qc�Z�(v��!BY�/
)D3&��i&���Bz rZKU0�%��oh�>[x:�u1�sT�/�Cʨ�i)שU���O�t8�M��Z(k� �k !|NR��c�Y%eZ���=�Quͣ��ߊ���Tt:1�*l�;���2�S�D�
�`Z��)kԀt!�1΢�E�%X'�p�5ɧ� �ג��V�c UɦY:����RW���*:1��R������B�-�f*$��,ʹЦ��e���S�7�sM%2rQ!��[�@L _bK�s���h8�Rk�Ҩ['�q�I\JӇ����adM���&�d�Um���L!+�c�ҬC~N[��qZrE�eC8��8�f}$E�5�~�=\)��)�*Ti�&���ՒE��V9���A�T�@d�ZH�E�e؁�!)�9mN:���?+�/�i�������5`�@>߈�fxU�_�*B�%��W�s�W��l�$-�ģ��+�#?N�pvq�3��gB�B*J�
�EK����(����T�>��b�3r��B
��0ܴfB&;><ٕ6m�TLM�U�S	юx�d�I|~Ek@JY�Eq U�#tr�-j*��MSN�Th6�zH�Z�"Z��J��Q�����O���7ө���-IG��I���o���-zw���=�_��GӉ���~��6�cQV��XN+jZoR�"M�m�H�3Z)���L�b���G�7N��]3M��r)�����Ǉ���/^Z�}�w�)s�_���5�=����So��s�����2��������w�?����מA���W5?����~�����P��!~���>��������/�D���W>��/���|t���7���ݾ�W�Z�����������S{��[ڃ�0l�����o� ���.`g�o�F)1E9pK�ԛ�sˏC�H�!��o}��N�:4�D>������6���    IDATG�;��N�?��?����[�\�z�F�G��v��I��ρ�k �U��s���K�G��s*7q~�eU�m)�tLK��$;��l+Ѡ�"7��Ƭ!�g���X-V�a��L$HM�&���Du��U�)�I'>[���j��Ia:��%kj �*���Y�?Z!g���BE���BLٜ�p�� �F�DJ��H{ث�Y̢l�5�8�݈3�Ȝ����pN�v�f�[VvZKn����S��\�9m�{H��;���(�롋����\强!8LR:X�Z���׿�_B�7ϟ?����=����ɑN�~�i=�#�	���sˁ��/Zbjҁ=��*�Dh���ii�����-Էe<�1����ڝ��~2h�$�H�b{�W����+,�nrD{dS��X7�C ꯶�rYB�!��tY�.��Mi��,7A!|���2�p��`�,���A�Q])p��*���)�*�+M�1��9l+ȗ���5�]@!�!p�[µ�r��6�����oM;j-���	Lu1���&��9|CT�%�����*�A6�h!B��u
%��[�p���>����y�@�v�����o|����*D��	f���)� Y�p�.��"+]3��v���B�+�(P�(�^Kl���}�������o��]\���6�՞��kO��.dW�P�Mm�A�Bw��rc��&����N�m�O�P�B%ګ���]� ˭�h1;W!h��u	[�O�^�x��������N^���Ѐ�a�>�u�td�"[ߠ/j�5l��Ϸ��o��x*�%��N
���"d'1m��m@|�g	��I��s��(����Ín�6GuQ��ߒM��p��A��u�B�:8�c���B@m#��;RB��T�����HQ�Ŭn`���K�`j�!ǇcҴ!J���N�5��:�~
�2�MV����SV�)�g�H.����!�C���EPΆ�8�a��t�9�p��>�HT�B�D��#��iCE��VV'��z�s�֨�t>��!S(}�,Kp2h�NG���Iǅ �&K-��F�:I	q���5,�_�*A'���J��X����!�����{,��U��d9F�MH�	}�y�Z�%)���1&E��=�J���D���ɱ��#e�I�T
kʉ��$eZ?H��N:��ɯ%�\;,�y���	f'%�0�(K��������	��c��Sz>�i�D���)߰.�FKpr�A���ځ�8@)����BQ��C��Hն�t�DL� 5����F=����UK!#�Ιz���S���Ǆ ��<O�<AHN�j,���e����*j�d�����^���gM�ȩ�Ko�SCnu�ʚM����ޤ�VkL!�z����U�Lc�88��������F^:�TY�1�r�#8�;�I�E�"�!˨t��_(�L:��Q�,$Z�]�Ӊ��1��m{�,BjIa*�ɶi�ea�N���X��)�ۙ8��t��Y�?��BVbY뜥i\K��C���)�[��L��2����*��B�{GA4��l�l�@[�,�`{���ʗRVN]��t '����cK�n%��OJK@Q�0��-�PJ���xL��|�e� �YS)��8AN!>�&�,
'��H��F��pRC0e7I*0�UTA�@��]S�[Z��VL)�R^��aj䳧��g>�j)a��F�>��TJ��cď�ơ�VJ��� Y�o!r��DL��4���Z�F�4�C�[V{���v��r�=�B�6mC��B�@�����5�lJv��5/*������ʭ'�^�j�*�%����8~�/Ӡ�^sW!~:p���߉��Sߨ�m��o���e��8Rث>�)���~R��Em�hH�9����x�όt��P�G��%%�ݙ7S޲y�I�]����eT�/�t�Z���R )��e�hl>�9�B�m��S+�&���I����f����v�O�c-6��p��Y÷E|����`oe��vt>��{r���@O�ۘ77�LI�X�_�<>�����w����;�wo�<�q�Wo���������#��4o_������������W��x�����/~޽���}�ӗ>4=6To�.k�?}�(,��Uk�� ��K��iEҏ5�[�o�1/*��DJ���GJ;,����j�yG�;m�8���&����쀢N{���^u�V�'3�������_�ǐǑB����p���;��;�IUh�2�E�Չ������(�Bx��r�+��U��	Yfx�ђ�ym	>&Z��Ս ��C�*ib���
����m�	�R��M�Ƚ�)�/1��
�=�ᨙ��b��fTL!�Q4D�ւ���j�����U۱8
<����8s��<p�ӈϿ&���)s��'g6|:�A�s�E�d�>B"1U��f�3�0�Y
F`֔��p�U�Գw���N�p&�q�f�	��b�ٞŉv\���
��]�h���v�ǯ}�k�]�96P�Y4|T}���o��ok��L��$q7��|oi�N*=�[Z��)�1�MGǴƖ���BS��3h7�{��g����~��_�Gʪ�,O�Kݠ��F�c+�`ՠB�kJ�ů�x�"�z&�
!BuLYJ��
n V����X�=���0e���^'�Af%�,�,�5�	��A=��Ƒ���IS&h�ttRJ�+ѶH������!|H�&A:�m�-P:fE��*�lxm�Y��55�8X��*��7]�5 ������I`�>PbQN�R�"��#p`)�P�NG�'ǹ��s?��?���s_I�qmwF��&��苪�ONM���1�r��S)��rD�4�N$�(a�ӱ�cS��3���m!���kRD���1(��^~pWzQEqV4M5�#����.~�E�s��!�#NܽU�M�4RS��[�!+���UN�60�:Dk+*
�F�� ��2����5�6������ �������J!d�fC�:�q��
5�`��.;ْ���/���������e���,���w�+�VQh��RD>��g���s�Gzd%��l���8}�FY=Ȣ��JCTD� 4k��Ņc]����DdC�P}R0���gӑ�h
��(&S#)��O�z�CbU�T�Ǌ�j�%*���Z� �l*��7e�v�t����1���Iuq�|��@#`J���~!Т�����?�s�Á����P�օ�X�k ��� 6��m���<�p�*������C��eD��bѡVɚ�M
r
�k��ɿ���v�S{��M��)�u"��Ԓ��z��Ƒ"T'un�J�
5e�%Š�J )����-��l��s0�s�f�C�]�)��)�Z�WBb%Ѐ�ҍp�:4-M��ZY9��I/Wo����{�,K�<�̤�Ԅ��@�	b���Q��	3��� !hhꕙ���>�����$+�˖-��Ϲ���M��j���U%�c����pK�NUP���r�Z)ֲ���,}KK�!� Re'x��N���XJ;s� �+��VjY8�]a-p�zi�"��qn]-��BVUG-A�X2AR�*qY��u	�oK&�y"��@�gpl0q�.b3��u����T�F��8��`x�<��Z2����������5*�iY�63��8/�𙫬�8)�e������Kx�N	΀|3�[Ƅ�;L%b{i;���!!�r5�+�_�|Y��Z6�*��n0|1��
�8	-Z��[ǌVǺ��Vj�E'��BU�A�3Rn�Z4o	/�<�8�ܙ����]���p��C��FĬskH/jr˼r�& �],U�)��D��K(˔��oZ�F��Ȃ���vɜFRVE�%���Ɵl"8:p;���R�Xhu����b֓��8J�ĕ�LPjW��Je1�I��m�}����D3�N	"�4L:b�Z�I�jD0�妕�<pd���J{�u��� ��O�x�(t ͟攣�PPص��j��9B��DХ���Ⱥl��j�����7X�hDFX!p���𻣒��R��>`��!��ł��R�dJ�����)��ȪZk�]��Gn�;��̣��k��B (n�@��R=m�ZT���G�T��@�`�J�31+�/n�𪺋.Wut��]#�1�� +7���D�B� �V(��lW�玻l���S[a�L�'�x�R\!P���ڜd�����B��ƣ1��ͩD,[��ڲ�[�# ��j#��M�眥X-,�6� 5�b�PC�B���y��٧g��,���'�S�ȣ<7���b�r5?��6���H�����������_?=�'k_�8[W��٧����Of�g=C>�x���������oR��/~�_������7g_~zxw�>C���>C��!���ߴ���LN�[
~T���ی_���1����K��ɺC�g�O�Om7U?>L'�ޗ�ՆP�C����ݵp'�L��yL��X��! �i�"k��H
6�]
��9e�h������(oIn�X aR�\#1_	�Y����cJ]�s�Á��w�b`�TE���D�a Q@��{,�`�-�Q-�ᛙr��À�V�T���]��-�e��l��D]�D�i6N����4	ܨh��1��y�T� La�xC�6�/e�>f���Rj~L�ł�����`kԲ�\���nYU��$�U�RA^Pm���S��3)�l)�q�eӉ���������֢c��1[���A��~=�R��O7!Ш�#����G>���?z>���8�"K��������	z�ͻ�>��q N���]g6��쎒E�� �,ьg� V� �$".p���B�HR��\�7��&d�r������������[��~�D�-��ި�1��;�
h1m�}�`����{1�׏5�!ڳ�����0�h4q�� �]�b&Չ�=K���1,;�� O�K^���#L������*l$�!N:#PK�^����y�F�cYB�
!��K� `���!�K����lZ3D�������Z�'N�t��<����h��N3X�K9��T;ri60�ժ�H�<0~�X������=*��A/�n���(o��]��%D���s���-(�z��*���Y��W��m"X�ᇥ��͌�>�IdL(h��fq�|��7�7>Y��{q�H�f�aZd桰�ę,Z-h*��n����tD�i`�ha)+����À%A
�� �oG6�.n?��Iů�*�|"hD��e@)�#� �Q�|˳�g6JóΪ 5��z-e<���أ����E��4|���ro����Ŏ(�ܒ�B�,��[�v!��;UkBjI���?������?�����x�m��h���������0�i�
���f/N^Uׂ�W:�Y�yF���O
����J��� �!�hIӗU�è�}/+�|qQB��t斚"�� � �0�K)�A�h`_��:�2�i�>�&��E�g�����O~�d��T��؁8R:>�����S�k�r4�tח2D�������_!� ���r�lwJ�X��}�j�Y��%��N�U	�x�ً�؜+TE
��t v-P��`�Yd8٦��f�b8�R��8��IIY*	)eK)�Ry
�O��8<~:!ĉ�݊
Ǐ�o��!B�ב�x�y����vCv��&E��ш�N�����@��Z}UՎ �%Xm��g�v1��H	���t
 �.X�J���L�X!JR�6�B%���T����w}�c6O]�߳4�P����F@�״*�I�X,���I1}�;��Z��~1�<}�N�'RUlxKVm�y
�	�Q4q�E׋�ο!Ó�̌��<�}+ŚAɶD����K�������	\ �.��sȧ�~1��l_��i3ʪM�YA�b�Yc���T1���b/ަ�h׹MPU�����2�Q�T�L-���qxU�#�!��1��eS�Gn�,�L��� ������iK)�5��g[�R�����	�YG��l~��<C˫"� �D
x&�H�����W��pɟ#e@��^kj	���#y1����8e�+)L���ƕL!>D��O��Q�>��{2�:L��dx) $�u|Y���9��j���F�2g�1����!)[
��M-DmӖ��+�EU�y���� ��mlٌT%������ʊ����,�W�C-�N���l��W��(|��=��4�����Z��pq����X/k��i�3r�<�r�t
��e����%@)�9�XwU�����hb���Qir8K���K��*�NH1���]�
�󥺂�p���e#,��$� h&?O�s��ᖬ��*0M�I�]�����!��UEH0�z�S�ī��S�V��36��k���mwb���R��s��L �)��b�B�k�;*Ogxz<=dRP�E"
w,��Ū�
R��e���E�d+\�4F�ÛDМ:%N-�4�ٲ�ұ��ȇ�4u�΁��i�x����YL���s���F�3M���ӓ����H���˯�}���/�"��+�ѧ�̯t�~������}S�p.������_?��w�p�^���o��}�=~�՗���_\�L�	�Nw5���pԮ����� p'�wKTR-���LFG�R!�D��ỵ ~FX�Y�;��n�Fڵh�ߵ�#P�7��������x%�jT�XS�������: q��1�3���bl���TM��gqx4& 6�y�@AxS�85Y}��)#"�r4	��8�z�_
X-���̲�ߐ;7F��Phkh�ӇC��MJ��XR�T�����~1�Ǉ���K��<��[J�ZWe)`	!�E|�Q`MED�d
!-��7���� S��T��!�����9j ����`��|Y~�5��G��[\a���^��#�#����Pw)Ȼ�{����U��f�O}�L�g8�F�3%n�zYy��oo���#&���79+�n�7��2��&�0O�ߤE�\����@��滟e��D3�%�y8N�gwUY�NoY k:�[��G�bx����6�Mc���g�����JXxK���ۀ�:Y��z
��	��h����u�׻�i/۶����4��q�2YR1Y"m��ۻ��qf��"�E��q)%Y��6?��D�.@��j��Ȋ��)�tb)�vui�tb�LGf�Z�@e��@1Ç�=ŗ)6��Z[��A�,4q� K	����i�'����^�ӑm��dq��6W�q�3x���kM���\A-d�,!d�;���<B�MRR�hy_��X�IUx�91�:F:Ȟ�(��)�`����F�	�/�Y���SF#迪`�IJ��Zʫ��}/"
ZX��&$a1-1�Bm��C B-d}�a���W���=MH͐���T�k�rc�	�"^����[2K��&p�
�&��ej)C&.�˅gH��癙qR6� �(�����IybbJu���+��3!Ψi��o�g��0jj���� �T���21k�&�qMIMD�T�S�&�����S�,�Z=�(��و��,�Lܾ(p�Ju�Ї(�]!��+G����)�r&pi��5d4"�G���p3GPwb�c�u�BP7�.nW����`;Y)��2�'���������9^�}�/�w�uQ뿇¬{�ӅШ-[2KY]��,6���3�h&�%�/��h<>�ok\S�Ԝa4U�CXAjv'�xR|"bx-��{�IAL�f˪��H��̵h�v�����@S���4O�Ȑ-kG9<}L 3g��PGA1���9�l�0�
y8��Ǭ�� ZK�b�!����w�kQ��)�m
�e��@�uF����EW<BwBq�wW(�)�&�r� خ����� �,~��I|"5U"`8�²f���R/�p�lɋ�+�d�wn-���Q���-�9�=L
"�&ǅWr��:�ף��Y��U�����B�k��dbR�c�ڑ�)<ԧ=����FAm�E��"H���"�T�0̓cٴ�����G�v������11�M"�8Z��oH��NcH�d)����W�shdy�6�R8~K"���B�H���OvG��|V�u �*k&�6��de��h�    IDATS+��!>Y��(�Nc'L�-T����1��4dHǔ�x-���*%��￞*��v�)C���6.���z�� $&Oa�����$(Ū�0�{��lxZ^Շ��l�Ȑ�l�.����0Y��\\b	�mf�,�|�������#���6�l۬
N�o�4�sB�W�U��m:),���MU�Çw !)W[;8N��c��eL8S
�h��[.�Q�پֱvI!��͆C
�ؕ�w�4Y-%�.��n	�²���$e� �%B������X^9�a<�c� ���ب�U����HT�g�p�*޴���L9rx�U�4�I��x�<�Fe�K1��uٱ+�K��)�*D�#�_��cE�������K�����7
�k�MU O��4�́��=o�~�����<q!l:)8��!X�5�v-kW����1y��kQj�T�`
����R������TS�e�6�,�%Á��$������Tyk�9�<�/�O��a�7&�}x����/^�|x�����������'��۹wo߼��͋��^�<�&��Oj~z��5�F}�	���%?���g����|�B��>zk��/�|���^�T?{�_���|����}b<W��ri�f�����v��"�	��6�ְ���Mq�Kw�e1�@�e��@:O��.@j!�j��K�P�EfU��v�4�@��q�Z �b�8�@YKoV��{ks���F�/�-�l��kK��C�8��֖4"���!�Jz�~i<W�q�� TKʲ}%����dmP����ZK)�4�"��-�����W��W(�����!�){�־��ӎ/%`��C�=���a^��/
�q�d��V�gj����]ѝ��rKd��,)��:BR.%fq
���o)%�jR��2Z�{��5FR�F��uY�-qjQ;�*}tќ�.�LN	{��#$��,Pm�_-�[��7�znH��|
�I�0�:����ޔ���^��'��c>���v�{9C��xk�3a�)U�Ȗ��7�T�@O3�fk�h��<�BL��{�F��j=0��׺��^��I��1��F�,�O8��O�įwhF*��ε��6�Y 7=�Y 0��Y�*#�!F��b-����ѱ�W|��0{��{���0�&�e�D@��m�_�t�4��E�&lB
b &|ʑ�U�H%�]�:aL�BLfi����Z6f�Y	���fcȲ�ꨐ"3:�ŝ�X�@q��!@��+��H���S=e��j�rjC��]t����FY� ֋`{�ݶc4jp%�9������/��QLj5�9:z�J |�����ڠں.&۴�M�!���'\>;�S/�^}>Y�Wmdc:���L��B�H��CI�A��qϋ>�HA�;gH(���0���Q,�k���{{��y�t��Ю
�i<�>1���~�a�7�Sh*A�Y*d�85Y����
�<�n˘jc�����Mk���U�D�tѢy��V@���њV9���0���Љ&��x|1�V�8�eG!��_�NrdSe�#t
�D �u�O��2)�G/�["ǧ�m���nK�#��;��S�,�oI�U(��@��cN�*�l�&�1�ׂ�R�mjd��Ad�����p�*%6�b%�v���ᾲ���{[�S�+��e�*��M�(��<g��*�r��<>Lu���;%�bVa}�;���u�nxK�8�MA��̈���_�������+4Y
�"2/���Z
pf	�-)�)��βk�D#�nTK�)\���Y���,H��~
`ɤ�j/��QGNP�����N���1yLr7����k���BdY嵳�v�W	�v��j�����v�+d�'��!�t�����[@�#��R�N�2�%X��dk�f'ܦFk$�	�j�3��B�M[SS��v����2��gۈ ���]��1qȲ!��e+G��m<x�������0w٪ �e%�4d-����gl|)�
���_���`�U%G+��)��G֋���КBt��HAa��R��Sw��T:uAӑ��S�%�\ܲ�ŘU󗥣N^
'5�h�1eG��b�F�	�T��H@6�l-0�� b���T%e�[6�����
�wf��k!e8B��&��!ĝ�e��å�N`�&`�M%��\a�ݒa6ɂ�N��)�Rōi���m
8q�W8��$�_���ul��o�&��M�]��:L����B�$��a��ъyL�K�<DL�ZMŮ��^����j��R�3jY�o��� �[6��ST+�ߖŐ�*����5M�$@�cj�%�B�X��jlZ3���I5���Ma�`����-�J�J6���WhY����L�T}C�1���iY��6 �1�� �Tk�B���5p"������j-;Pp'G�1R�&BfM`<�5^8�����I���0)t)��0�q�L���zY
X���+�HA��؁�R�=�+�V9�����`��:I��WoƉ�	�	T,+E�����e��q�L��)����@��G�M*#�f"5��b�8��dK�	�Ď[���Ĳ)̠����@z�nIG!������}MgB����/k�Џw޻����崝�[����O����/�������yٙ�N�=��귾z��هw�?�>�g���i�'6�����8�;����B}Y���ˇ����_����[��I���y��O��SM~���+������i����f�,5�}��~��˒��XKL~��S#�|�eᖵӚ`�:o7a�o!�p�l��%��Cш�C���%C����Kd��h	�K�,ނ����]�pf�¤#5R,Z-���)���.�4v۴�$��@	S+�a��K1˼�s��3:��e��Q���v8���H!��u�@�uQ%����I��v�!������\S��"#X"��U�_U8�KP��a�_@��חsN���կVoy$����e��/����H0��p�]xK%
��;3���5Z�l�
�� {�Z����X�y5Aʊ�hΰ��W����7��3c�FQ�)`]GA)�e=@��x���$��D�Jǡ_G�F�,�4�l��2�<���)��"/%�b
�Hd4��6��n-O�ƫ��:2j̯�����Ec;1�.�sz����W�ߨ��>�=�b��{�ك���Z�-Nz{��,G\o�X��b���=ܕ#���%h�z!ؘ�v�ç)���ZK%G�R�/��۲X�PJ`)�V�e��uY�rw�<f:�t�\$A}	��N"��jŬ�HC��\P
Ba������"T��H%�$>�� ��WI�Z)�R1��cn�pL�a�Y�ĩ9I%��M1�M�K
�ƺLɺ���]�_�[����>���兤PIU���<b��O��%p�j-1�!z�z�j䵩�H������@�vTE-S΀�V(�֜�����*�������b�@"^b�P(�#�*�ű��^<���
�,Ŷ������oYV����{��Tɓ� ������oBe�m߁��i�c��ȵN�̄&��T-�ʩ�yʉ#�(@�7�hp�,��Ŭ��'NGߎ�H_��uG!ը��Jxَ1��,S��5q8�3�#���ʛ_,��T�$�Ra�h]��b㩲d6S/&�ר֑)W(�r8�.�.
oi�v'�YY
*����Wb��:���4��5� W.0^- �Qp��:U���S�䍡�Z}U,P�ܜ5�p�a��ƺ+�(LӍj�bӚ������q�m����r|"	R@k<����+�d��!}Q�@G-�$j
���V6B�jGX�
�U��UtDżT�}e!R�r���x1�s+�W��]�������_�@4�D��i���Ny'	O�M���tiZ"@!�[Ƽ2�����{��-�X2)Y��IVP�esbB:�b�$��R���:&RK�1pĂ)@�|׍�N�@�	x��zB2�1��ĵHb	��'6^|�b�s� ��J�W��H��զ�ǧ,��%����|�Y�����Ɠ�)į�]�~��ؾ���R �$�7[U�
�4�r?�tj��&L3��x15V�Z8�<���GS,h)ЋaV��`����]_����f�M(�D΋+�f�4��v<=��nආo�1���Z�u'�kx)̮��Zn#b�Wݣ����f��/��) ���TZ����On��zU������1i 1�8�J�}��.��{@�q9�Z�j
d��a�|�8.����,�&�j��P�H)�u�G|̍dѤ��BG
T����__`�oL8�+�|B.�ǟ���@q�R`�F��6���o˘�b��ZJ%%�d�F��H}��OB��{�^Jy�zm���K`��l��yqd��Đj�L���������Z�V.P�~đW�b;h�h��`'SU%y4�d+/F+kY	Z3$�o0�5�F��
�� �������	�i�&gM�*��+�6-��
!�|V<q`�	�E��pā�;�'S������$�ʟ%�����@�@5�,C��B�j}q���]k)��e�!iJ�Id�fX��J� �y?��!�cٮ��ƣ����БBp��J0���� ��\!�H��  ťHm��Gֲ��|<yL���R�H��Bq����Rh~��Yx)8�k�s7
Bp��oGfJ�!/^��Ι�N�km �s���ߓ��O���K���O-�G���w�޽y������g�oޝ�����k�ߨ}��{o����
a���#�����_�����_|���o������¹�j��l;�l����'������o���BJ�ڴG)KU�� <[�.4�,��u��ù� S��BBo+u���ј- x79N�Fj�l��@�����4��Qx'-B���(�dm�R_]Ȳ�GUf�8�l `��!u�4�vj�F�(��H����)��m��
M�/�d3��R�.f7aH�1��%�A�� H�G�r�����#|�R����L�{I�Nc�_�D�0%t���(n��WH\��녏�K	�+��gw�Ų���<�շ81Ñ����#,�������e)@M><�i�,3KA �p�w��VR��r��E���6�l�1�V(�EܒBfID!S�܋Z�C���^8�Jd�|� %Vk�f��NGL���_�H�p�{��B�@�6���i�u�`���ip���B���3�w'<���������[o���g�W6���s���75�Pc����3je��{`!4MA�1�,���d��#���)kCw�bL�&�����K- hY_Hd�XCR���9J��4I����@����EsR��q 5��u�1�-�%��w!�<@$�-wԘʳR��L��D3� �4e�6ef�b%d!b)3[���HD�ˊ��ф8ʁ�����2D�h�V����� A,pD�Z6yj�1	��|����X� ��7CAY_�Z�f4���_r��b��оy�ag|W�c\#]�ڎT�/���u,t���k�^K�����_Ӌx�A
�F<P��=ڲFۚ@G�^��-�-��D
��~�6��ld�6����u���l�h �z�@�e�j����Q�/��/�a��^w���+E'�R�a��]M�K�T��>�1��	�݁;mC�O��7�R��.&��X�_/x��擒�3�h�&�1����)���:�2~R]5��(kG��
��r%�M"���.������0wE��7@8Z"��Uq�9B�+w�4���2����R�د��0L[�T�![�-8g'�K��^7F۷C����HP,��&���S����3�� �nK1�	J'ۄ�x���@��^��<�UI�k�K�M����*��)8qI��rhH{A3d_��B��^h���za���i��@*�o�R���UI��Wŗ��S�YI��u���)ED�	�8����3������,�#X��,>0�j�)��M��yY��5��Z#�ş�e-�"�\��rS�a��x��/�@<��
�IA���QIL�Ԑ�x������@J�@���	aG�ʊcZ���WoI�ӰT���%fRb
h�<f���:��:���$��Yن���h	^�GafӅ,T�I���a^E��Qk��)�%"�c���vJ�7�I�#T�]�5��$�ǐ�� ���R�h�;���
�����# �+���!f�� 3K"G�T^V� 3��j���TR%�R���\�N���Պ���J�	�.�.�wL��U(�WX��
�� u��Ԛ&�9L��9�=MXLyL2֫T�BVPU4R��F�T
��~ʫ�'K!Y' �u�_��ۣ��D�L�/H\3)��,Eᴹ'����#�R����[4g:q��������m��q݁���Jh�\/`�xw�]|8�L!�$
)�QֲTM-� �jq��WXI�81-�ӒY2A��D����:����
!���K���FA�y������"��&0�tڸe"|"F��H�I�}:U"���]Ϗr�$��Bjm��t8@�Ej��9A��RNs�M�/ţŷ��e����l�l8�5�L�8B�]���@d�+�e��4'��-W[k��qn�Qbg��$��N'�eǞ��Te����>��� �0�j���p�8�u_
XV!M�`�`䥪�l)(�dJF�6U�V�ޮZ��K5}d�@���(�T�l}q�0ٖR�4 �:�	D�����"ďM�x�X�~c[�#CpၺȊ��G�4��Q���q`�'��$���|���|�܃^B�s���޼}|�\�/^�i��ُ��c>�>������5�g�^�e�g��.}�ʼ���ԛ�o����^���7��������=ֳw�������c=G��R��i�v9���3<cێ��8?�v��:8�� ��-�]��i��kH�k�����e%�g�U�H*&��h��e���vݓ���	<"x�'A��.Z��2~��|B@?���J�3K�R�&eZLY�[6 O����w�%Y&EǒU������!��T[UR8Λ�.��M�����ë&�)`�]&4����e1-7�ւd-�LS�� Mmg�R�S��8�J�Rb�8��S�4��E ���i�q�T�����њ�g1�*�$��څ��g�-�OJ���l6L4��ˍ��
B��f;�./�iRPI�r��@ kS���!�w�� �����m|Ϣ/&��n�����|�=��N����[uh����ĠC��S�D20�c��CBP�`=) 0gJU�l�|1߲��6�CT��u�%�`p��^5�Y��h/�[~MS�-���$�75�ӟB�z����m�4	r�H��ے�4�!P��*븛��m����$[L|�lȖ���z�̲I�u��BC�Խr93��A��!+ V�\��x���+�À����WP/B
��i
ֽ�8Z4�B7�%Y|�|Y�r�#�%B���T��%���Ѵ3 N[�R%"����!ƨ]�R� (�$��}����Y�d�H�d1<���s��
yǛ�=� _����eC�G@n�j�iG�
�)#���8�E�����
{�1��Ȗ.��m\�X;%�����т�ȶ�W�}���dm�Q����Ъ�T��f[��*�I� ���x�ji��[*Q�B�Ub��V"��c ��Ǥ� ��vS���8�������6}��÷n���7�B� Ba�B`[�2!�R`�}~�����>���$�oN4:M�8�TZ�Dдv�!��������ALd��G��FK� Df����4���k��"�l�LP���� S`�)��B��(���ly���@y��d&oY;{��d��j�C���E�H�hU5d���W��f ��IjD� <M]v�� �|O@�!��3����f�5j�'��.��5���h�Fڜ雤׋�~�Jt1��U�h��B�Xm��D��+P.��7���o;dᲝv��L��8����:��y3pZ�&2��    IDAT�R�W[*D��pd �	�#�_-��BP����)Pc�$�Z�TA�5C"-��Ȗ+Y����B�}9����d]�n]K&�>�\��2M]*��R�����ğ�ZGG'���pA��ilF�-���w�J	������T��۲�J5gA
�V�uo�FU��	��z?��#PKP*q���NKq�B��C:�d��T��P;%#�/�d�Ť��+y��@g��)(M�8���8�RkqLA���g��֥���I�<��\Lx�����L����j�� �_�ǧAH�O��gxX�"Yq�@��k�T��V*�t��:�*�W��R��'2�JH�2y}�e�m	�P�Dx�,>��Џ�N��Z�,��2LHA����!����7�^
�8P;LxU�8
Yd����%+��<�A`@�V�$n���w	�6�%K�/H�ɵ��,�x�����-�1C"j!�7�%��ز6� ��I��5�?���G�2Sug�udbzd�ǲ��iAD�eY%��MP,�T�8)��� #'��l���ӧ����Ôet
���A���f
�."���]P	M!��-���}�Z��4�Ȗ����7	��e�-13�E9����Q�r�h_I� ��Yd�H�m�b%L-+nxK��W�ע�,��iv�1����/�ڞ3��[a� �j�K���X�o[p�i6�Z^@���]"��"���.pRL_`:-���R)�Y2A��|�<2[ �DK0��0D !	��ބMt�xDT_�E:��5��T����M��Ch<�f`�eݕS3����F�/��8���Y
�W�Dj�MP���O��Y	q���u��%��A����$f1�;K���oC>��$~+.>c���7)��>|�O]���e��|�;�}����"���g���ϛo�����z��o���P����_���ߗu������&y���wo����o~��/��W�y�͛g�}𾨿v�����<�K�����O�kx��K?�[�Ӯ�)v�����;�
Ų��(��R|C+�[ꥩ���)+O�~_��
𽓀�m=�-�c
���-AFB�:Y�uD�c�8��M��<��<qRyx3X��duo��kQG����(dp`/f�L���qq34�eU��F�H�=>C�d-Ϳ%>pKR��f�̢%%n��j���ڑ���'�)DGXY��m�(�,�M��BA"��ǩQ�aR�c�Z�f:��ZR�G���h�5g���W���T1H8R�3���@N"���N�m�^UA�8�r�eR��oNȽ0Y`�~{�����@�ۈG�����p���ݝ*d��6CyT�<�h�Շ�y x5%�D��D�o(lB�%��HaO* &��L��,�x��F6d}�{��ZӤд����U(�ɋ)�u���L����?�S���������g?��_���ޗ�$E��6����$��C�~���Ah�m�V�2(Y�)��/���Qn�l@�+��M�1a��,�)�Ϫ��_�.�h�LӒ���n ���!��tJ�DӕQED,��6���I��}�4�}L4F�)_�zc*�5S�r٤ 	4��r}-KY��@%��e�Č`(@�i9�k�h��p�hJ���_�&�d�y`]"�vP����*=MS����	7�%Yg��%ٺPhf ��i�^i�/NWS �]ȟ��&�Յ���9ɒ�)�Y��mA��G��?��B�?@P�c�|�v��2�J3�9e�t,���J�7@&/�05^���C G�WG�͉�Q�-Mfl4s��e���O�yt79���R�]�4)�O3����hh̐��k�Ra��Z��5��Y�Wo���?��?��?���k-�;��gԴc�(_#ʲ�%� _��8��t,�t�����"˶/
�w�o#L^A�]"Z�j�J�8|ݵHa^J��c���U��<�	���f�K	X:� S^G�e"�ũ��(��!L�J�u�NI���-�	��B;�^���FSʽ-���8��B�������_3�����$t�@�~4V9)"�<�F�&)�c(�ݗr�%�A/F 2��.U�rxY���Ju���6 O�����S�0��N# oY f�Y�d�y��݀P�FyK"��)���H%좗�,ڙ��	&�2~�q��p��D��G���.CN-&_��x�J�u���ˣ]���w�A��d��j��U(h��CP"�jG]/UN��1�0�T�"U͜º�Y#) �)N|-Ԓ��@��Y\ЎxF�EKjUf��
��*�fV�0�Ȃ�'q����I_-�Uqn��X��/���0-+�56�-{���vW;O��ѴK�b4K6}����S@++�V��|�mJ � 7yUu�-���,�ZK�]�L�*�iŁM� ���WR��
M�$�1����v�R��@�g�/�auB�ۗ%<S9�Sy��p��,)7X^j� Z �&�9P��WU9?<�do�@Y{����m��G�,�I�v����Yow>�9�>N"4M����.h�ɥ��lR�3WU��D�1�ډ�e!�w��kM��y爳��c�69}6ZK~���e4�6�.�����K�VwUL
���k'��4��Q�eӏ�'�R�d��kK��p1M>3�Oj����"�gt�*$�����q,�)$�S���ik��e�d�8�-#���c:[h�|}��W��.�}#���?A�i�px48ù�����5�8$��V EٲZ��	�9o�~"�#�v_	���I�oى����^�T�~d��i���N[-KS�ޝ�,�/�Gf@V�@��i����1y����JL��)$x��kS���6�,�]�{���O%�7��x���,�(��吾c�SOY#�F�F���F��l�%��k��"%��vbc0���PPwY�����6���Z�`BX�M"��%</�L���5�#�󡣿%�7#��.���g�|��W_<�E+��goԼ�����={ڪ��3|�O�^���O@�=x���ο���o[�1�/\�L{�,��O/������=�_������_}�����i����_�}�Χ��	p;�����L~}�ؿ�G`��l��Zh�!+h�R;���p�!d5�e�<��z��}խ%�t6���W�U�7��]:����?��!�O�	�I��>����y�W����v�7�mM-Y��f?�KM�{h?�яt1�,|����� 恘d&+F���"L�K8π���C,Sn�;�P����� p�)�D��lG���2�fÝ$NȪ�X|����b�8u��*�o)&� u)��.{"�LM�.��p�����u�����_��3a�	�͓x"!�{������M�L��|�{�t��pH�4k�&H�3o�9����e����3���Q�k���w祺_�r};�8^�W���Ol/s�����T^�J�H��o6���� �с֐OO��5���v5���g&(�|,e#�vE�_
U����K�4� Mw�з;o�zv��X��г��b>S�)�ΗRB�3wrL'Zz$at�LY;4�Ƭ�D��Ɏ�%��A�|�֟^��R�c*��
tF�ʋ�U��K5� �RIً ��Uu�	"�״"-Ýf��P��>��m�gRJ���چ�I͒rݛ�A\6Y4��q�tǁ[�~�f@��lny�{�V�e�r�,Y���b��M�bِR�)��6O��MbYU�:@���t*��;S^s�q�x%�B��������rY��9�O&��5�-5}����O~��G��Fu-�� ʁJ���K�TUqĲ�&3��5��шx��C�^ɺk����x8�n%b!��H�AV_K:4���|x� (�����8OJ�����WR_�ڵ}�@aOp)��6-��Έ˚S� ���L0����uK|Z�G�Rh R������+����w�p�Q���
���'E���C��Kuc�q�z��yx��hF�h6��
1�#tJb�-dj
kDQ[�7�^�R*)�"����/�����:�Y֙(�p:�*o�x8&1� �l�:��,Y��R�Z�&�K�����;�>��ä�q��p�x�;�:J�iU8@4�),P޾�A9>Y1s�-f#�q�Y�b�^���!\SV�*�Ih$�F��BPS��pT�!b�Ԫ��sƙ�	�Te�H���L��*lk�iDk�r}��M���#�,3�,N:�[�@,NY�;.�� ���+,��'�«�9I�f��;f��,�i6g~U�͓߮�ǵ@���H�ā�3�ӄ��+��6��Y���V��T�w��D���v@A]��v���d|s�3��m�6�,C����N�?M^w��Mri�^��bzYyQ�U�U�a�Ey�3�f���TS�ZSH;-h_��4F��l��i�"�i�j�����[�1q�Vo����L6ZK�Z���8h�ᚚA*0}ˤ,�[����3$��)+"�+��,������C��]j�^�EGW�ͩJ�o`|H1�y� ��TbL�^�-m�O�.���1,�i��"4���H��5J$��k��< E@���Ev�+I�Ǭ��m�ǉ  �+�P�%�P,kI_��j����B�y��č��e�eS����m0 ӝ2��
��}������D F�<�#[���oY��ax�򆔅0d1K�^�f
1�mW����%l��W�^�hY�T�{�.��NL>P�0��㙒uCp0�Hʘ�K�Hŷ�����*��'g�(�R��~�b��#����TX�_v;"�I�c
 R�.��%��f�G	��B�j�����3[��,M`�#�]�Z �j�Gn	A`��(2�@��,��-�^���z-H0r��X\!}��I'��Wy���y��I	�L)j�!�'��l3$k)+�y�)Ly����]c�Y�����K��*�d��ZY��-'R�NN��Z�;������4�	ЩJ��.V��I�ʖ������:��m�"��r Ӊَ��q�<�g��ٲa�d�f�*���DK�}�����z�j^�_�g )?���H�!y8�/���'h]���x��W_<�fЯs~�e��6���O��_�s�����y��ό�b��\�/_��4�'�.�O��x<�Ҧ����o��s�S��_��M�|���û�pވ���@�WX|��������5�����d�޸Г�.;���	 t�|W?�.8W��]!��$�F�70d��S�%�*YL���[m@��.P�SL��m���0�x�D��M���|�]��o�&��۝�,5��*a@|�N�����+`V[�|`%D qd��AV��FH�Uǩ����@�5<D UIUp^%�ł��e;3\�3?_;c #@���BФB�"HAd7� 2�K��f�K��j��+4[��J5	�3K�Wq"|�|R��zV�eY��J �i4��k��|`|`/���� �e���≤ 6jq�+�S�EUt[�@-����r��m B�����Z�鵯��������f<dL`�K�K��3ǁ���#�=�b𖵶��H��s��)����@�j�V��<�4��;�|�t��|�@)f�SK����z��ڣ�x{�.���ޜ����=%����>��t����y����?���M��7���ڀ~F1���H4��ƕr�:�脗�)��c�۫7�G�l�hq���N-<�Tj�Z��i`l����Z�#>>,��!��K�
<����'W��a޼�wAϐtl����W_�|������x�����g;�ǿ��0J\�^n����X��"�m�vQ�;.�Y�����j�5q1�YG:��h�|�]0��X6�z�C([ʦ&`��	,#`zIt'�)C���@�ōc�i�]��;>P����,��!L#�}�Z�ܽRv]C���'�z	�S-N���<q��Ne],��E�Z�E�-i�XB�� J��/`����74^�^�5�Z:�<S�c��a�^�^}�ӆ�6k�:�v�=ऐ��Z�E�;M|`��O� �0MރO����-���B}� ��Rm1}1N����t�_|��V�\Uj�LT����ZjĀ��5�:L�څ��og��	;|�]LU�ёUuߝ�i�J�x����-�Tb����&���t�;�j����O@Yf	g�-U���(0����?�0[8���1Bj���S1/�dh"%��cd��[j���ǎ����P� bZWV�OĒ%�C����)˺ե0݇�*%�5�e^58��]@UX��Ĳy8��_nx�jU1�z	�RVkA��=Ad
��.�G�?���}�j�"`
�Ue`/j��W��,�^LU���1��6� �
��X�Fq�!˷,����ĥ�h	/&XY����*�YsJMG,ef�B|�0���)��w�+y�iR�|�+i|�0�#�*AC�����T���]�����t�3�n*H"���
y˺H�8|� R��^���7�<P�%e)E��ʦ�)sh�S���3A|�R*�f�b�1�'nˁ����A��D�i��]�(!�d�D�W�P9N����B6�NH��R�8 �aڹ�1��{l%�8S�o|��^���q,\=/e�@b6�%�Z=�o�5���d#���{I K��,f�#)c������){Q�D3�`R)�WU�&��~qT�ԥ�p긾݊���5���)4Cq�q�(T�^	��@S�ȶM%�3)����]�;�d�J���^�׋�T�vV���%��*�D���Ť�$�{�.BT�Jx]�kZ$;�,���uA�["��z� +���O�X��
�ϣ)G�ע�80�lR��]	��)�ׂ���Vn�W��T����qh
�����(\��T�עLJ*�B�4��*����PHYVydAq;��M���@���kGM;�|�?&�%y�E?o'�_٘z��#�����i�4�#[0�S�U��.���J�3�<ܒ���$��8p���WM���O�ز.��1���!
�^��h�D��������M���Jg��dYO*�@�}E�/��lgkI6�oi��"�Y�||A�I������e��|��|3�
Rn���H	"h�R�ɫmTk^#L�@+���!�t�_��#�d�{���U��M���1�	9N�17����M�~yH��PI&�I�A�8OwWu���}�W��,��k?�Y�Z{�.�������Ou���R��M
e~���ϙ��4�P
��4eB2ZB����<��=���UW�֛~�L5�t�/��
R�^��;���U,�H��5��`� D`҇��JAF0fpL�n��9l|4��ce��5�r*-e�*-K!c8�t�Q��16s�w*׫-��M��sN㹆�w��������x��<��޶���<�8�:��ޝ���=���f�W�/���I�����;�~�OY�����:���}ؽ�QN��g;�i}}u�����/_~����o�_�n�vǋW��1�Yϵ"l��o��y���3>����G}d�}p��F�3)�Z���_��i{�>�������XV�Ry��IY�ϝ�y�Ɯfjy<�sQ�M����O�9?!=�"�BF8e)zп�t�u�qu�d��!BM?���B�]8ZbR�r��R(�9�B����4M��7:�D�V"~%8��t0�
����8[pUG��KouȘ���E�(T�p`��V������A�4_�c�c�h�V
�1�D`�hE�K,�XS"�h�
��N�h��:�yQ&��[�s��,)���i[f'b�@�[N"F��D��[�Jlz�+�>&��f�F�E�Hk2�E�*2`�)���|R��������4u�{L��B��#�B���(˕��gp�=������˿t����?|������6!Y�
��O8x#�O��O}+�B��IIW�k�{��	1u��㐅��������S��s�4O��|��ͧ��޽�U����BG��������D�I]}���R�_�Ԋ4�i*iZ��բ(����O�o��e�J��P�7����    IDAT"0N��z�6}���?m��[�N�ԈC(�Xϕ}��韣>zm^�y	>;�������]'���+���w_�׋��a�޸�[uǕ���Y/[���������p�_�t��ۿ��~����:���.�������j���i�U���V���t[]����VH���^��$�i�$BV���$�ĭ[�eU�H��qL��D)��V� 5֏��+��(�Á����*KИ3d�6NSn= T�&E�0�c:�*�_T.�R�|�Bp��FO��.0P�8�Sم�"NH��9�c#�l���X�Q��g��CЌ:A��m�]���-�#�p�f��D�F<#�G�Z�p|��tn�8fj�����٪ш��\�6Du�f���[��C��dN�M�R�՞(���J�1⸅!��$�
�qL9[M�a@��*}���>9^3�B�m���ψ)�!%�X)�R���
�_!�ԉ��(\�4G��٢������7�)�d�Ɋ�HLs�<� K�AZB�Z���@W���D!L:��c
���$���¯yg|�'QH5"|)�S>ӧP)��(���fR��������<�=�\]mE�����_o[��`L�C��"w��ض�6�9�[!ׅ;O�f���Jw��^)ʋ�9��J��v�keQ#�d����
�DGP:��������V��t-��$�Z�)qY�&M�l� �Lz�B�!iZ�������L�Z͟tĺjՖVii�p��[�hS=T7fǺ(}L��1��7&�MȀwu!���Íu;�8Q)Lc�
Bk�#�"�\b����˅���o��X'�E�J��72
��ptޑJ�,��"SV�ɭ��!�Qm�p
EK�8|��Zf
��ސI���R���~5�_S�M�+d���h�ib2K�U`2���Ӗi*����pL�"��L'ehsu��6ل�ą�U��X��-]��[_���!�ڋP��,�E��r�0�X1�Ș�����|��12�E9-�BH�h�VA�	u��RWr�!�5ʍSb��Y"��m�B�)�9E������}��h���v�`�i�7��|)mo���5ӘE��*Z#0�,�d���K�,>?�5:�?%�c��#��ϯ�\%p𦕨ωƩ%4"���S����R0��)&ĈP��G9BS�L+��Z>�S2K�Pm'�� �锨�\)8�nkr�0��I��0H7��L�H
��e7bʚU�J�V�tF_�M���$��7����DH<�O�����Pmg-8#�j]��	m[m2J1J1��K�i�p6�׼10���9%��&����T�t꭬���0j9�;�WN:����*Bp"�F~w	� ��f����U�y'�h��
� Ĕ�4_K!����&����.�!�3Y���Gd+�d
�|QY5�瘶L=��5X��
�ˁp�l�Ȧҍ�q�D`�9
e�Q>bʯ
��G�1�є5ռL�~K����(��\�ݤh��	���w�F�~���V���r��X
�#?C�Z98��H�n�+d$R�������/TzL�calo��*����F{�t����=;������{���g������̩泙�GoW�}s���+����lw~���w�/_]{Nzs���ݵ�V^���Lև���Y����|G˦�������.�e��_�����͝w�^�x���o�[����~��_����b����
�����m��~���g|��:�ۖ�mam�N���F{�b� T�=ǔB����u"y��/Ԧ1�(��t-�Υ-�o�~����=��� +��)�Q�h|Q������1��)��dR����G޲�AT.�S4:h�JԪ#T�A	`k7b4OA?�Dk�;?Kć���7�h����+�<��08S.�X�D��8A�%�͈&a:�fN4��T�8���ʷE�R�ZRR6�Y�����v�F\<���8�8��a�z�n�߲�^J�)iR筅�Dբ �i�_�h�z Z�h��M�J7��CAn���)n�D�~D�W7S��� ���G<_R?�Ʋ�#�3?q �էi�)�g?����+ݵ�"u�v���>Yk���'�����������G�n}�`�ɟ��?n����;�؍^���u��O�RKLi!�!�i�P�B����V N��ʨ]%�τ��X�����|
J�f�����?�m�'Ӱ�?�Q9�ޯ՘(�_�����_�է�~*k�3����X�82*��DPR��mq:���P���JG3�-�J4�K�Z@F_"AQ��v�D!�R3BJD���u߁ YMnǩ�w�4���Ϭ����?�������h�sf�� �Δ\��\M"k�^m����������������{..1w�m�h�����Q��f���L��	2;�Y8Ӱ5��ݦkh���Id�ji�4:���b�]�ٲ�.��k��e9L�!��*�	5B�hF����o-�;�a҅le 2�%=D�� �F����r�,=��$�fiUAc�@8�	�$�]!�M�B>g���7jn+.�ޑ�Q9�������5 �L|p<�P�/�;���J�T�\M��4�Zܚ�UUj�m��萈�`K��U�&���NLY�F�tȔ0ʂ`��A�ճi�#]筢�eE	�P0��S>���Y�p;��{��k��XE!�]	�l��_K���FU��ˉ)���u�gۥ� �d�u��L9�8L��2�Bth!pG�b?�8��U������5�)�RZ`>���)q0K1Z�����4�ҊN.���WQz��:�d�2Y��N��I�oi�r�'$��r���6�9!|Lj%"���5j�S�"��V�:Nu�VM_"�)$ZES�8)���p�l��2v1�r�A������[����.�A�����Q�e�z�ՉJV��4#����� 9�v�Uh nD勺��I��3=��T�J��P�1G�����2-q�l{^�M�f���yS=�1j��:Fk]s�r��Rk��LK�׃qhSR	��z�~:�G��j�.$q��|��B�K���)��Y��A���O�T�\!��F��Me����@!|�V�)�N
S�#QhjJ4�O�k
�3��ᄴ�)�c8�*&�4|F��E�kE�˥o9��0�,#��mB�)�U�3�ZE*��6��BiVȺ��)Z��`<e��j��O
_���4ၫ��Y�����#._.��T�;"RX�ȝ$�F��t �8�m�(�*Q.G"��BD8@���8�@ph�T�N���V���[�񔀓B�Q烛�%�/��Uf����ګ
~4#�i�X!�MS��aNKȗ�u�BL���y���z6V�i����"}hd��3���1�m������T�_
��D�Z-Dh6A(c ��:^���r��*]?��Ҫ��5�[Wu���b/ʉ@�o���aSQ�t�,b�8K���l#��Ѫ�H�􀀯hRU�L4H�FV!8�ϔ�Z�q�|�Fց����,������3>d���euh*�V�zƔř=7m����H�r��A�܈�S"'��EX'�R���)YL��X��͆�"Ҕ36�֡HG��z%"�_3���B�����\h�j��A��Q�J�63����"�NS���@��M�Ȓ�BRF�@j��ʂ��4�x��g!�)�BH��y�8�8%V�~�)��8�l��OEZ{8��銛%"�T��9]����ژZ8��M�}�<��#����x�\���[鐦|U]�F��f�@@�(d�r������hq�2�$�ojČ��Ҝ������Ȋ�`)B@>�S?�� e��6YB�����B;�O|RSEd������7�ݭ��=��ͳ����8w����۝'�����wǽ/Γ���ҷѺ\�.��.���'��ͫ34�����]�{��]{��O�\�?����� �Y�?�.��t�,�3�?��?й75��7�~뱄�ngHi�Y䤊i�"��݈�I���m4�h��8�EU!�/��q$�e���Q�a�\|YY����RZ�r!@���|J�Ƕ<:�y�����{!For�bEuhT�%г�6�[JM�*ц���b��dN#Gb�p"G�[>5!>p�*1�*�HS�B����ؚ!�V=G8���QȈ&�6J4_2�|&�=AC�L!>r�hd�l�=��F�?=����K�	1M\�NA(++�8�.B�3�^�ą@S.�2}S~!8S�I��'�,����š �hl?Kq>@f]Mi�v�ˢ�ΐ�(�d�U��
���S(�hL�ҍLh���P��`)�u%�Ǳ���x�B=��A�Dd�eݣ���U��m�N$����~�������x�r�~��Ǥ<yCp�S�w-S��N���Gu��@$�����(�dx+��k��3Y�N?Y�vN�S�@��
Y�J8�@!�uh�2j�;���+�������j�%���ۜ�����B��h��q�Ր�F�LT�G�hB�
aj�!)�|�DBe��Z��m�S�4-E"���t% �!��>�B ۋ��\z���!�&�����/;�>�y����0ߍp{����6]ݥ���\�l�[��U��h�߽�^�׌s񎎗�y#�R� ��)8��[)�hG�9
�̖�j�R�BE�%ʲ�A"��,��,��2#>Z�Vs�����1�5i*ė�C�RLȖ�xA�N|`d��5�ƄLE�	L*��,�)���[O��l�)r���Ӏ��o*7)j���mg�z� "ʤ��1Չ����nk0���1�D�Q�&r����>l���3�����:��dQ� 
�L���g�$N��D)z6%�w��H���Ib��0�d�~�r?B�#4֤���o��m+ ,�s��"��R�~*MD��G��V�b��!^��F�p�%U-RW!)B8�md-!�_.�j��5V��nc��N!#d#S"�Ij�|��aG'���_Q:Q�J~>�@��)�P�r_�*�!FL�3�7�,�NL��J������ϐ+gt�ь8�}"c
)��C�e5�gC�"�?�Ԍ&��@=��!mJ���R��%���=��&��7�k��c�	���v�NKEki�@�(�+��,��&�Rj�)+�\������|4?'�O�v�F!�|Ӆ����Yj�F��S��$��S���cZ<D��X#?���Z����7�V��Ħ�J�7j�����C(=��A��K/��P:��e�����r�J4B*�f|Qc�1k��-��M�ǔRN�8��.�p��'�T������4����֎S���5Ja�4
����4�k���i��I_�u�ƙ�(>�1��ڛJ1�ᔫ�)T�8.%���Z��E �F��r
%V�,�9L4qN��U�@���(����q�n���͔�`����0͔bD�:N���.EPݔδ.� �KR�?r!~�Ƒ�O_n�1CD!|����S�X.B>�MWIA$"p�@S�4�s�LӉW�(����7�	��(0��FR���e�fbʚ*50��D�6==݇!s*a��L�1r�t�`L��)j�o9��)�+;'�U]��"e�2����t��m~}�ct�e��c<��O�~�FP��!PC�����P?�<=@��8��W%�!�i-e�f$���eʨM'!�4����8���5��k��-+5�����)�Oh,wv@(�J�g��N�L��h���>�x�7Ef�YqL�s��*�V�D),�Ib����-j���.��:p�8	�̜(����T�W�N��	�l2O��N�ժ>�M�kX"�Z�+g�2���_�V�ə��4�+����}��8UL���F8��M|���8!q�t�f�`�I)�FJ�~���U�!���4�8g��IG瑍�0}Ә�!6�B��ą3��HA�a3?�-�4@��2�$ׯ�~�is$vV�"$��$���MT��"q�E�A��Jg��K7�"0��§Pz~Ѥ�3%��>�9Sz�B��e��-J�&Mk �1>�i��8�lmiz@�ٖ���@�,gӖ���v�9{��X_6�_���t77��~q{s�͟����Y�����f=�ܯ?�=����<��㙎ӕ/����c^�WL2����{���o�_<�~���'9/._\(q��i=���v���[�ƙc�ɮg�V���-�y�(�.#�����&��UȺ��%�i�J����oJʘl{�H�#R3�����<�"�.�[2�8?ĊV����0Lof|�����?�3������� �t�����$)q�hL
בt�	QRϵA._���F`!�����g�����ij�V�t4�M%&M�A8F=�!GK��C�K��A���:���W�#'X�`��q>G
�q��W��43ā �%�Q�Y�Z�`�'�����h:�k��&��Id��F� ��ӏ~I
_.�ƤaBX�u�)'���\LV.A�	�O��h:�	q��p�ڥ@�RX͐E+ķ�D�e&>��6��)L���BE�^�k�U�£���׀ꦭ��w4��/���O?�k\�KRY�����w�x�&
�����g_��C�ڀ�˿���{��>�S�n��*�ӟ���-\{�k��N��m#)Sr��ګԐ�
#�,jLǪE!��BM��G�D�z0�Z�F�L��R�&-�H�.y#ӻ����]���
�?��?X��ե�p�KN��ҁi����Za���۔c�#@g%�Y�M��T&΁[�,!>� �BF8� ���w".��%�I�����K��%����������^��k�_�O�U�^��V8����9u/��}�ʟ�5���p����vGx���gAo�����_�<�T�a�pv~8�:����9��\�n&F���&ub�l��Zw`������P�r0���Hi�����[*5�i[�G>�'�-�-�1�<��m
��P"�~���0�� �� ��h|>\?��������l8)(7ՁȐ��2�Wwka�p��B�4!5YP�p� 7M���)E�I�*�۱�9��Z]�P�Z3�1�%Q�4�A#N�͛7�^�����g�r�X�P�D���s��`��|��&UԀ�,ܔՒ%(WW����Ft8���0�z�:]ݝ�\���B�30S��ƺ4#����z�"djTN	�RL)������?�2��C��SЧQ���
eۅ�m|�ʂ����dr����K��+�c�h���+_d����rm�a�9�p2��鹐��L%���A4�D���O�E#�#JGz˄�ZT�t&�ف�T�i�8�=�g��P�B49��F:h@&J'N>͈_kZ?p���I�$
���(Z�%���,>���C�Z� pF9'Gb���O>㏠�"b�s��� ����ޖkc]Y� �Ag�D4�d[��l۝��ȴɦ���p)�:OG:�8�U�f4��z�4��6pD��/�͔��:Of�8�Ӄ)e6��4[|�������d8K�S�&���A:��0�Lq"����f�P�O�Q���|Yc��Ӣu%�aB�6����Čc���L�������.��s/�g�K���%n��s�8-"�Q�D��'?���,�R����)�T.+��фԉ)c")'a������)�͑�1����,E!r>��$V���ҥĄC��r�sh��)�?|
�;'-��'<��iN:D�Y+�P~Sc��i*!��u���IV{���>0Aj�h:	B��U"M�i>��9����1�-pt$�!pR�d�'�Ogz��|~8��M9�B3�\�B�+�=eVo�����.�(�UQQS!S�J�4d�^�-�Ǵ����d�~z/1D
/�D$W��>
�a��iUV����rj��/E��o�7e�=-:�v��.ħ�tZ�d�q!BU1�EѱVD\o�KX��ˑ�h
��9��(�s&��Mq�M0�B�zn�T�\+eu����'� @u;QsD��R��!BƲh2�h*4��J�	2gD��YR��d3����pY��8�h9�c=�7�&BY�%�z.Z�iB���3v|8�% k�XM�g�-�	Pn� �r���E    IDATT֘��1ª�B`���f�Uy�!��-�� �'�מ���P�G�Q��#~�3�v�4�,>���%8`Rtr"H4�ފ6V��V��Nȗ�)LJ��'�hj��8~Z�Pc�v&������E��}|`;��Y��Ҵ�e�����ʩ+�m*�� Q'�N�
�P]��W1#5SR�������p��O?5��+���~M� �����LT���f����Ӣ��ފ���$f9���p�g)�TQ
r�D���7J$��)_n�B�Z��a#�_z�_Cj��t��A8��e���"�kf����\_z�qq�:�ӽ��w��������~���W/_�������/��{�9{�裙�Z{�D���;?��
;�f{�]�7>Dbg�����fY�(t��IN/�������?���Ϯ��6Ws�E�n���~#h���0������>�qp�E�^��/���v{��р;��=��]b�8m��&a#�-mۍԀ50R��	A�K�����*j�>C0փ�VAD�3��|�;���w9~��A}�k�T�R�.Cg~ʢ�H�0�������4��v�|��Y �k�#�Qf:u�E��B0]��5E+$
�#T�U�B��
~���<�K�V��M��jC�:*Z���T�Ң�)G-L�ƪp4&%�(&����#�DY��h��m�:�T�$���AYm��!f-�?ʲ�ˏ �u����lG�,D�м��WzV=��t��hJ�C[a�W��\Qc)̊r�K�5Nz�t�Ɵ������jV��%P3��Y] ��]��2��ܸhzQ���=��я~�dRFvQc2O��Mi=���YǝSE�r��"Ru|� !D�zh�� ��Ս�(�q���gָ��wN]Eho�&�Nu	z���J�h�c�؁6ұ��������`u�!���^�u{��$l�FURF+HzU���șl���.&��br:Z���[�t���	�K�h��ڝD�*�1�rnO�D�hz��qh������z�����޻����c�_�~�O\/���_S���U�v._��8?�x�㜾B����˯���}�s�z�vg���������3�����%O��n-�&��&[�ג՝�+$v8�Ý"��7W/n|��}q:�� Q��5"P�6� �D��S�ȫ�fme�ms��,�NJJ����J��|SxF���sx��㴃'�Iy9B��[�K-������t�Y��r��)
�P5�Y��q�Ӆt]�k�cW���U#�ru��
Y�6�CM�M)pں�ג1B��O'��@-�\�\���(K�&�O��P���E�t]հZJK�9��Sjڶ4�������'nĖ�^�=�@Yp�v��d%�c�jÊ�`��jY����K��Z�����������%ˡG��h�:'%�b�Z����iw��3u+�`	���+DJ�����BFE�-G��U^|S�D�EO� ���(G�t�˪�D�ސ�UA��� g��ll��B6��-M�Ѭ�V�و̦s4|S _?,0��`䳚!>��z ����"0 �ԏ�KoL�('{��	%ʕ�@Д9� h8��Q�n���t:���@��g��4�М����&�@�K�2:^��4���/0��)$�ա,H}BLe�r�&T�i��K9�\Y9�tcjJd����'�[�ش�� Z�*�1K��`�*�k&S8���B��9U�0�5�j�U7���)'�%@b!�O���%���?��QÏ�`����p��m	d�)Ch9߈o�5&s��i~)|���(��-j�s�5�V��5ͧ��Whv2u����@"�s��'�R�(��c:��z��fgJe�8c6!Y#��cR@��N{e�ҤwݥS�%H$\J���F�ڢR�,��4����t���X���!�(ʢq |f-�� ����VΘT!�6�hY���B����4��qJ�&�A���9����,>�xdc�4+��Ԩ���#�[Q�V�)˭74�U����66šP9H�7� �T�4!l�lB#��%��S�iu��unl�JY��NL�فPB�\<��| N��%���^��5Y�t����U��g��pH���tR�lm�&X{���D �`魮�Q"�h����,��	e�?�LWᥧ�?:�i�TD�68r�!�=m#e!N~���D��!^��*�O_�D
lrO�IV�ܚϗ�U��R�Z�$9�i���4�,��)��E�F��S5�����"��#i����k��Ж�M�SnU������r��Rn�iȖ�N��F��8J ���r�B�~R巽B���8�(�B�q*a��ڴ~�q𥯎��T�U�(=M-Yl����#H��HO�� ��8M�A���dRZHS�M����O�,?�tgQ�4�G0%"K�:��8h���tSH���©M?C��٦G��/��y�B4 �A������-A~f����������E��Q�j���&Rc|4.u�9��$R�1�Fk*Ā�)ڹ����D��%��O�C]Q��QB�F]	U��W�i:��*�\H
��!f��o:#������+-�/�fW�7ԝ����:G����_.���_=�[]��ݙO��?vq�kh=��:_�Oi�_��;��)�{q�]������ �zw��޽����ί�����w��K_�h�_����݅߅}�O�hɓ��Ю:�>ä+*�����
��aj�=�i]�1q�)�#�(��n��!���8���|8�U��j%p�m4��_3�Ј�v���b�C�'r}�ѧ�~����+�-b��ތ�t讘 �4����-ͳk�C����W%������1�SSט8�f�7m�LG����	jL��"Ph�E�e�)�#D"2fk�H	�p�M'�M��q�ir�e%��(o�	ҙEQ@�pRP���YK8@fJ�M����n�O��рUQ����-єZ����R��v�-��`j���0!�
��)kh�ɵ*Z��;���>�h���ƭ�5�(l�	�ֹQ'�I8)L�T%��"ǈPƘ��ۢ]#��#xF���7��Pj	�N�o��R��C�z�,׃>�d�Qd��_�c+�f���M8��M�T-L���F�������ފ�J���D�4�r�q��*�>9FQ��\Y�W�H�T�4�rղu�׆Ȋ����Jٗ�:ml���3��}�{��}���|��2Ҫu�)���4��������V�Ķ��N�
���DR�C�L��ENs�2��������/�@��!��`U�_Y����3�E�Nޟ\� ��mI7�럡���V�;���߽ݹ�	�E��?w�*���l�^_�|�틋����]��y�e��2m7\�k'��'x�p{��}�����%y�>_�������z�����y�y�;rWd�[ۅ`���bu@l#2�G��i�;�ar��B�u+=�4�TJ`:���u���%�q0��!����U/d��FUZr|�/�_�̙h):��Ζ6��_�,?!f��ћZm��9��鉋�����:ܴ��
���Q�k�U�_E��@,G�(�qΧ��ֳ�#�>u%J�U#H�F
M�iw^��>�c���.��:�+�o�~�HK��"�
�.G]E��s�Ʌ�Ja�+�B��@�r�A
S�9BVo�k���8ܿ@P!�,R�KDӀ&��'��"�骞U��bǄ�C
���PE��Bk1��R|-�0���|N>�&���/�hr�hL`����8)��H3<Z{(T�B�K�:Y&d��*����>k�8,����Z~NYm�f���k2��t�Ʀ\�n�)Ӊc��Ympf]�RQcu�4�B'&d���+��*V(��i�B�v���3�Y���@?�Q	������:�C���omb�;&#���!�%2!�ASA?���̪����"j���#H�\��	[�r��6��J�1Ji���'���I'�ߔ_�M�E��	��Cp�ڰ��@�OMn�F����_]8��#R��[�8���W�*� s��D!5c�O�6��J�0��3�"R���ApX�HϨ���B�	r��nx|"�JT.2��ρ��X���lK�=͂�*t�NՆ�V
) ����?�B�\:���Mf�����G��?�ÉV�p#q�l�t
��Buk�TSQ�,qQ4㤋B��n�6����cdf�����8)�jZn�t�mG�n�����G��"Ǥ�J�Ĝ��B#(���3m�F�#^�[��*�Y�8f�V1�p�V��t����_��F`�:L�[E>��v�rYS4#D��Cw�D�B�d���'���g�+�y��j��	�'h�(���ʄ:R�s��q�5�g5�0��7*g���3ߴr�pX��ȩAL��k0M0>�C
�u�D���"LbuK	���OHt�pHQ��c���#�eB8S!��VT�i�`�$[|��A�1e�������!F>�f���\��xK+j�DG3Y`���<��j	�)g�%~˄Wt��N��5)�=�h��G�s�p:'r����/�(9�9�J�(��1�LS
C���D�����mi�%�����#�woi�)w"єkOʚt�|!L�6���D�2�5R�ƙ�j%�l|�Z8��0���CH%�G2Z���2Ī+�?-�9~�B�4�g4���Ж (��5��Jco1jU[�ڴJlj��j��ٵk��ګ�F�jS������~{�����|Ϲι��'�c�I�E�J�Qy|=�h�L�)<+�l�X�,�R�W��d��lv?���R=�S_��:�C�ꓻ^�h,2$+�����r5I����M)`(R8֛({��������ujd�<~�5SQ��Ŵ#�EpVmF�	|�Dr*��n�D�&0�%KB�'�1{���t��R��V�1��4�?�j�n��_�f��Ŝ��/�39��"�H�mﶛ3ƛ���<"q#C;��F0g�	�7~��3-�����,6�P=�����A�ꑧn�'�Զ?v>��?zp�}�,s�[S.����Uϋ�Ŏ��!�a�L_�F9kY�f�V���7��X��x5��f��Z{S��P��ٜ�����β�uk$ԉ6��Y"L#�}��z�C�XxH�n��%ʣ�N��{��j�:��ȵ/}?h��JCK��[E�)jG:ZR�6�eq�����Ucx4���C��`��?e`>,��T�ϐ�e��g�;�t�?
/�4���Y��[M���R�^�W���Z�T< ���#����u���E���M$?���e�
���D�>�8Ūc^�
���}.)kW�����<�'<��S/�6�L.�+�-����R>B�?��
e��/�&��f28B��w20�W[�Q&�#���T����/gy�>��$%d�v5����I��<�  i׾�ǜ��v,v���[	44EwN��Y����?�k�h�/��L�t�k�N��b�da���?��w1\c�D��7��2���,8Z�S���A6ORć/��)Z�+'�1p��U�C,���鋷�*�'�u���q�a@�d�1A�z�B�&��3|߹gZ�F�(/hq����I��fM!�};�%�ힷǏ�/Z*�mʠ��%"!K��8]��tw��9v�J�4|Z�(��.�f��j�D�<�t�v΢�~
���+������^�>�~.wZ��]x]�q���ż���+?͊�E�րʟu��_�y��ss��4�(^��$�;�����u�F~�8c$܆ʽh�=�;�+��Y�N�jk���䙅�bѻ�`s�W�Zإ�E�����V�������Y9?����k�z�~�����}��X���/�`��%=+�c�;�}��g��`w�/�?>���9%�ؚ���5�R��FOG�D�Y�M��_R��lKdK���Ik���;�<Wq.��M�,0�iDEN�*e�N�@�An n�ӧ�Ɯ?mg2�J7��j��mg��B�9�͜"?��%��;�^�v��gǒ��3|֭q����� w���܃���	���F��2�*��	B��Lw`Rd�(�{�����a�P�1�Ԥ����8������[��J<��&�(%��x�$2"Z��;�B�pk�k�' ��6lh�\b�^��9��o2>hRh2X41�LOyb^���G>�w���o�o>�W���,q$-��ڃ�R�6�~�1	Ʉ��_.� �(��������a�t@���I ,Q[�#���b	A�V�׊��+�vB�+�%�$�0�ZXr�#ժ@�Z�&�y���Ci\�F1�?pgw���PZ������W�c*N����+?^Uߎ{���P���͡&ՑPu�_�^Q*�T�T]`v�Wx\������GG
=��ՖJU� q�_�������F�ة@���#�F!�}��U
]wh`��v>�
�_N�M�f�I�����a*�=�A:�O���C��C5�Y�M<�]�h��1p�	~��9���Ё2��@Mn�<��Æ��5^O��Xx~TPJR��#`�z�{VEF�B�h庰� Eha�a7�ǵ(��z��͂�%��u���Tok���n��Oe>��$��l�[�8�M�?���{"8-�`/�H�E��/IG�3P�|�Ēt��p<sE'�G�
�x�B�W����x�T����[:��Ϳ&�q����G�������f6��cxe��G��
o�i�k�[��	q%�h�Z� �'<3��M%Pj?��s��A��V1h�V��;3�n��Z�k���Æ�.%x]����gs�^���h�p�=QV/�x��H�  _E�R�N����S��VթtQ�P��0v}��к2B�C�GY9��h�9Gq?�m}�^*
p�G�^f��c3K�a�h�6﯈\���xɡY覾��ݢ}��Q!����$vQ�j���>p������B}*�Q)�+%k�H���f���m�K�|����A&r���Yw�{nJ���6&.�=i�.'d����^�%a�70"�z����8?E�����&���^ʆ7 �l8�t8~�|2���G��\�|!u|�ޟ�$�_̯�6tHs��c�����]����S�P;�Dn�������������LaɋY~��вG�g��Lw]���i�jx�S�r�M���}�'w�"w}}ҹ˘z�����$_P�.���X�$%�<��Q9�7:��<�t������G��3}�+C9�Isi,��&r �FF�h��p��K�8����Y8��M��
GTy�do��8��H�q��sJ;;u��-���ӓ����U�W;]r^�?�~%�M�}�z�����m�n�m�{��<��T��o� !�s��8y�o�i^���-w�䶛;�˗���oE�L�������ᠽ�� k��Z?1�$�!��WSm�zS���?�J
L6��a!�(��@���'���!��D���l���'w�}	y���mh4e��ػ�n�X峼�
��y56�BX�T܆��&8I,�q.^9������_ٽ����`�p�ە'���V
�s��n��>[�v��v*�w^�~Rc���Ε�]�Z�6���M��y��H�AeJ���͇LEI)EXZC��� �J�qKL��$*6݊ ����Ԉ���DC[��h9��Wި�'��P��R('�g� ��{�CEQB-D,�,�z�kh�lM��nO�S��1�⺲8S:����l9���/�$��%�,@��NK�v���'#7Q���15W(�r��&�@{SNI����=s>����6Ҷj�t5BN	�ܯJ����@aN��pU/��9Va�>�}�W��c�+�FZ��dt$�Aǧ64ɗ1V�����O��9�
bMoM,,$�aK��^l��+d:deL�Y�KQ�Ų��cS�F�bR�ӠBrЧ8)剎�o�ס:����ް{�APq���2�F"����[����~r8ǔf����+��,��w4��@��}[%��u4�X�gdd^�g;��$����u�k�]����y�+�ujxr����"�=�������G����[���<���$�䢤J[Jv�J|�g���E�B�Q��魕T�5�w�~�WE�Wgc�<E-�9�/��:Zn��~~��|��U�<��͡��5���3��8�Dh!�}���e�r����z���_���X�z
-淫-Ng�,�+1b���ܸ��^�����̨����O���r9ˣ�w}�+��:�7o.�t�lu�M�yx��޹�t}�x��,�zk�ݿ�����Ny���Ή*�1������ūnÜj6�?\�l�����7���h#���G>%�q��F;��@�ʞ=��_g�:���<�:[��x��T�P�]ѓPU�~Wʟ~l��G��붔^�*`����4.�{�_% C��|Կ8f��\(o!�Pz0��?��ɳ���=��mO�i4�\u\e���B�wN�]C�<���u���T��x�
EA�^?�u�Lki)X}���K��+G���7�)�,m�e
����z-'���r3��&/%����*���g�s��j�VC�K�?�>�-;Y~�P�&蛣�����&M���Y^4F��=��E�N8������E���Yy�:*E'�3N�	H�R�AY���U%��X�skv�I�7Zi���'L2��9�����
 99�%��}Mu踏��v3�l}&I�g0g�n
l�դ;.�X�ZQ4�C���t�����k1�8�Lf��F2��1}�*&+�G�Ĳ���lq��>잏��e��ϣR��ZuAn���؆"p����yTFڨ�&�_�˼3��O���2�')7#׭JN�\���ܭ��>tZ1�r`2����G4��0OEi�n�5eG0��8>�}V�	h�j�X�<��v��}O,��S�j�3���oiݡ�ih쿇�����h5�X�^}�H2�J�f[�������K�h�f���d�
6��[c��ڠ��d��K-�*���vA��J�	������Mq�#�~�8Q��]8��P�=ls�Z���9��{���`�**���`K+d䠢��a�+�i���G��ā2�r�z�c���߯ۜ-1w�@<�6T�(1As�T��M�&TaN���Kn'�LQs!o/|x�ֲBP8i�EFMLd_�H�id�:�����\���;��Cz�T�̸�#-�H$������,��δ�L�8Gϓd�zP��{p��%��5c��=$$~M�����꟡O���G@2���4踨��jq�
8�F��[|��5�$��&>�D�����l��2c���l3����H��}�d������q��c�*�x��M��b�8Z�T��1�i/у��C�}�V����XM���v1�8��6���Hd�(�FI���J���R���gL�;���Ve� K��1{��V�Ŗ�����C繵.�8{ s���ա�`~�Pe�����ךX�dp'��w�?XYj��[N{�:,�����5����!�Ծ�p�	�������L>���C�l���ɘ	hF��1�0x�Pg��%�b�U)���I�B��co�܍i�Q�Խ��)�dc�q|��f+vE%s9�Tʩ�u�\�^�fda�2����Y�C�k\ӝ����R�;g�T:;/�f������]�J���uZ���4U�[v�����_w�r8�g�A{�7�fC���F|��M�����V���6����M�kW��i\�%����g�>��&-?�%v2g�#|}wF���Շ����(���L�D]�n�[�񉵹����q�ܾ�����r�ܽ6D����������ֽ�	�'���3��ٲ��?,�wn���^�\��'$��dl.+�ߢ��vg��d����Ӡ�kG7iE8�lRض�c4i=�D++w!��]���Ŕ��J���暩�w������õ����7&�Sܼ��j�"iZ,ր*��W}�=���6q|����'��͕d��a��|�P2�?%���g�d���>��I
S2I����!ҽ2�+��2�kj��"�J5sZ+7�]`��b��&=��1H��q�<�S�#R�a���e�=U&��"��v�e,����Ҷj�

2(�5�8�˞���QT�!Z���0K�A�\Z򕝲!�y��i�qϾ,Z>I5\���CS�\�P+Ue4�.S�=�T���3Шk$��njJIPl|Ȏd�dW��cN�D�V��e�;x�̤�+�L����6�!b����A�4����'�������x]���lĠ/=�jTyY�Q�fهL&TY@k�"(�)���n�-�����\�:�R�42כ������ZN���@���Jd��C�6N	设��D���#E��>v`a� �)\�v��'n6S���x���S�߉��=7\3"{���|�S�^���xv��SjLW˙���G4tN}Iï���m�rp_�
cO�.���c�`j�D%��9�
�(�Ƥ;���v�|ޝ�S_\w\.���P���hg܈E.f�w{�9���.g	[�LJ�=��v<8���N�\fU�ps=s]/�|���U���q�Ǽ�~��X-4��u���z�w�yE\<�v���]V��^.�.6c�M[O��$׍v}OF�kd	���G��������ߞ���m�4[��Ԭ��7[��lT�'M7�M����˃��W_;�8���O�$�ݜ���^ɐ��:��U�tb��_�j�뗆�1^7﬘��\;k���O��.���o�+��*w�5u��a�.�e�Q��R���)��yF�i��kB�1����j�V�pMK-��}��@����J���K�1�lX�������mҵo��c&�I��M���OUt��4!Z�<C>9�`�j��#�m��
5��.��a]�	�>p�K�%8��YF6��U��V�>�ci�o 8��M�F�9��T�����7���z��e^�.�L�e��o�t�y��(��@����(W���a�Hl�t��"oa	��Y�Bko"�^�3��֑ݕ[n�đ3�7C�Å�Op�6w	�4}�>���еY��=nӖ1O��J�s�����h�D#��KIB�����a	����U\������m�`�(G/���ߛ�O4�fc�.����X��^�	MB.�H��v�'����d�Dꯇ��}�N�Y��4LLhAx�.j��|���<����tf��T�N=hCG�(�d'�{����+�r�Wn����\D������^� L���7�b	X^�P��TZ*��z��f8�N
ތ
,LbϝxAQ�[�����C�}���!ղ����X����U"T��{�F�b����u�%�*���}�c�'_gZV��(Ø�Mt�M���d�Ts�w�m���)D�p�����U����-��k���Y��{�2m��U��x�?N�p��������ׅb,>܁
���>��&L>��Bo	�2{�.�~���YAJK1�[�Ĕ�+��RKȵ�uC2leR��H{�NՐ���=&k�x^R�Mo���Z(|�i�3.�BW���Ʉ�&�Q8�s����z�6�Cz��]�2����&6)ٹ�;ZxV���q��W��G���~��>g�HZM�r����/c��N�_�����i(����mή���N���/?��sn�|�ec�#V� ��*m�5��F�ԃg��@)�	Bҵ2�Eo� ����hT�E�L���!������P6T�Flb����t�3|Q<ȵ�H��O6��C���]GEKEw�<6�"���5�=Y`�P�Jf�}x��1��6�Fzv�~�.FQ���T�!֞r*��?�.r����Iv�K�Fl�J^X2m��A�'����c�K��rF0��ڑ��P���A���ur�Wt��KT�,�Z1N����
��ke���4�~�?[Y!^�) �c���L�F���Pʔ[t/��7�1<�>�r]=��Y��Xb��)D�o�;�ǲ5�!�l��D�̳�l ����Ԅzϸ���7�g�k<6�f��!��(.`�FD1軾���gu�1���ۭ��KA�R�L�Ւ�)ͪ�n����Jf͝�dR{(.Q�#���J�Z��VА���y�Sk�2�6(�yU��q�����ؗ����8��i@���%�s���-7aϓi��:{ЉFL�|�Ar�F�Z����Ie	ej(4��ML:
d)�+��M�h��ީ�mi�I�
QV�8
Rc�G�1+GN}�qv��t���- W�ee���n�����q?׉��m�$n��$�u��z�D�0�	4�U[����*�7{8zQ�u�C��YjSb7����c�l����ܲ��f_(��<��l�x�u;���짥��'^Q_�m_�~�4o�p����RR�&�Ƶ�+�a���x���S�Z�9 �*4��	2,�%y>V��I$�G���qyB�"��B>M�7�@ԽoY&�f�����O�n��˫�5s25��� ��������1=C}6&[����NJ�1b���1�4;��"�Vhʃ\�J>qEM7���� NP ���zϭZt_���ȹ�A�h�5Gr���;�O�~�**SO�� E��y൦$���t�9�9��B9�D��Tb��K+�De�SB��qX;U���Hq:���@��;�/�E���e�
�������oN�=�u�KKe1��0��RI]�ؒ]rP�ۂa�?�	�=Z�	?kg�>�������?��*���,o���U��̒�Q�g1+���fd;6�_�ߐ�|������ڧ-%���՞|!�5du����������~ŔF"�A�?��� �8���f:Ҍ�|�PA��ץۓ�O\{�+��U>졖[�V��gxt9�d��VA�+�O+8~��z�J|eJ�(�\"�D���xr�i11	ə6�<\����R��J�������o;U��F]�g��y|-&8׈5r�3�Z�Y�;l2��W��R���u�u����y�4�c[o�ɹxXW%��i�
�����W�������_��˵�;�iҖ=�{��wS��o�T����\S��'��u6�����FSj~I�e�n[�r8.���I��ԙGg^e�L�����#ጶW�,�\�{��/·,Ϣ�2O�:)�]�\��y��|����b$'����A��;`�|s�ڏ��6�r�����5۬���F�'�/�!�2v_fN��7�i��F�J?,y﯍G�l{z�����>�%��dݚ�v4�&��Ov�wd���dQ�:�)�(�Ԑ�4�Jk�R>MOF���"!�^Ӌ
&�𭪬�d��4S�D�E�j_3�A���7eQ	W�Q>a7�7�_:�� Ov#;gv@��Hpե���U~"dC��<"�:�Y�' �3"QVv1jÛ&��d��Ϝr��4OiR�b��ʼ�ua�hx��k�K�\��:zY���mհi�bB�6x`eD�@��0��$���vىkt�>�^'_AÄ�^��$N5�p>� �̍�;U"*J������N�8�S�D
xD�b`iw�3众�P	ρ�f�Q��>���
����1	���$�.�x�6�7�j\�A	v��u�n�:��mݗX4R��&��-�e+��Cc܇�[A�dUVqj\af�5αH��*��rU�V�q����5��L��I+U%��3@����8��� �	�K_�N�e�˂�U��VY�����{(J?�$��}L(�^ ������{/F�����GkMGje`w�^����S���m$��>����K�����18��h�u�)j�^�M]�E`8�h{�v}�)56��BT4��1`M�X�#�����s/�=(��3Dk*���ڥ_2��J���s7捫�
e�F�q�Y2�ʝ%��q��v՜�gS�.���R)`2��c�E���N�W4ආ�j[Zf#T��m�	ֶƔ�,��ù\g)�u�TX^Ŧ<��D�Tjd��/��*�O�_�����o�pr3"�(�-�������Um���w����0����W�p�rxaR�'P����o|�� ��4K
��9��I�R��U�+�����3�eX�(���[�X��q,.fD�?� 9=�U�I�_fE��D>�p/�w��8���a��mI�Ӱv8i�D���-�Β����!b,r�%��Tl���������j�X�%d|Z�a�G5�'\Q�����}K�t2�^����i�� �>�Š�ǜI� ���F��w�Rv�$��>���&B D���N����c%:�
�V���U���K"�}灍+_����'���۸T ?����hW#Ծ�#4U�5��n��(�K;�,V�E53�fbS=���oS��Gpl/�!a|���>���"SG�yE��T��#$�Q��U��ɤ!*����D>@o�>��ޡ@Ih�mj&2=��Y���Sr����"��rr�q�H٧$bs����HoW@x�DQ�!������ʡ���mF�S��L��˗�b�M@�H�E�����z͟��_G��-sa��D�?8O�~������ ���eo���Hfk:t\1����ͽ�k�/c`�wi������� .+yρ� V�Pp����"pP�1�%���Mϡ�n�ZQeuY���+;P�Y���^�&�	a���!S��]/��#.YY��o(N3e0��[}���5�ċ�k��]���S�l-��u��V<���W�,n�O�P֥�1�<���?&/v���z�x�������m�]�#��W������4�Tc�4�R��m)�@���z��h�i�y5h���TJ��$R/K�a�Ǝ��O�m��e����s\Ir:��G��������OrS~7IIԪ�t/hϐ�s�������-E���,���<ߙ�����J��4|�%��~����c���*�B(�� �^d
	����Hd��զ�|��,��k�t�fi�g�_����P]��QO1�Ro/2"U�!��n!�(Q�YR�P
n���V?��?9�ET�eѮ��Y�	�W��|�242�Ѥn������S�tP9�#O1m,�N��!�p�7,Z�id�yG��z����w��*�*4C-˯ #�ylC��q:�=�G����Ȑ�Ҩ�������st��Zw ��q,L��z������H =K�����
�5�m��TV�ͨ�D���}��a���S�&yw��Č�U9������?!�Ⱥ�4���3��-�8�����6�,������K��o7���m����҅���̑ ZF���V\C��^[5D|��(t���5�?����D��|��s���v�����6�}������C?��<�lP�����C��19/���vb:޹�쩔�����3���e��_r������O'Z�3�i���K=l�����Z�07�r�oVcwr��Wz�f;����<#���#9�O�{�r�Է��n��\^Uk��Q���k�12l�j޻I��i�;���K}�S�`��*w��Kt�_�����`i�0�;]O��x��GY��d��!C�<��6��{͡���ex�)y�������ש_��&f�r���y�4�3�e��-�>x�b�0ee]�MO�_���7Zz}��P]b���� ���4���Щd�݁��PhK�+�;sy0���f�Ɩ�OiI\�;��4�opϿh ���`DF{Aoe�qf��4�ϝW����UT�J-װ_s���M�rR�!��@�����QŲ�n��',�a{�g�OoA=�����~��Ǐ�	
�PEEk�2�$����(��z��[�+��ַ۞T9q� ��tF��O���_V2�0���)POQAg ��9^�f�A�A�z��jɕ��&�@"��A��\$�����a�Rx��8P��9������.�c�8��uk��j�F݃��p��c=�G�I�EE�H��")-n�b�ʤ��W �fd��&.@(@I�^b99�e;���n᥶�����CI�iB��J�+�#����j�O=k�2��ϰ)3Xޟ�A�X���j0��o>I�|���\���CL"���6�Ő��\4\Wl��4?��ՁY�T��2ؚK<����9?�+�mV�R�9�#�KW�vJ�!�_����N<���P��/������S�
Q��Bv$N��8Z�q�f6&u��h@U9�\��ILN^B	9�F�d1V�p׫&�Q�����jL�UBY���1��激�������4�-ý~�d,Ƌ�+▨!��5z�Z;(�V8�����.�bQ����S�=@`n�ўJ��G�6D��!�0�c�3�Xt�Fr�����Y��
GK�.S-�Wl7P	�F�Z�8�����<�%��.�@S)O�a�ڔOemLE5�߻bМ$π�������h�5�@ �'�9�(md�2Jlb'Dh`~���ڸa@�X( F��r�9(��j����|�&�`|tӨ�S�fכqH��z�X�D�;p;lV��' ��6�A1�,[��|������_\�!%5G�&����m���eq�:/����VGɶ.�b�OA[b�tƭab�>��!�C�hfށ��2p��{R�$S��	���}��F�|t.�Cm�N��+y������-�yʟK�:��6��p5)(-qR*�	�8��`T0�@����~���l���<*��#�}@�¹�,��4>2�L(+؍�EI���ě�*T�O�.��W���o�ļ����/m��^�E��@*��*������2x�-�-�������X�7Pg>�n�G����G�2�l}8���,L^��is<�[��vJ4]~/���I^�>��X�f!�^��1�I��[/q��_���7W�t�!�CY�y�<�G�ҥ�݊��i�0��,����z�Rz^���/d�D��ҝ�������( �L˞wv=�rh�L��;p3JP��~�NGT��3��bU�E	ke!���B�Pv�[�az"��_�k.M�k�p-?x� �1� �f$L'κ��K��9@k,w����š�%[a!�̶�:o�"J����䪊1�5?uUYbF�Ou��j��GH�7���߅��-�&!?�g�[�����/ZC��?�8SQk�}��6(S��|�~k�{��0&9�sMHc�_Ⱥ@̿�<I�����4��n+����@Uy��J|`_+�K���[�4M�	)��[(��"�%��6��,�u��S��SL���zD���6!���@��?h%������׻��94~��<wBQ
E��gc���`�w�#=yz���!��22�%�mX��P ����%7�lp�_��(VͶګ����`G�����m��8�'�j~2�G��-?��-�-���.��_��qa:2]Ӏ1L���4:X�:q�Z6�|�(�}���@ ��q��ifo�27��_��y\����
Z���>�`&g����9�KsH�{3G�ˆǓ�a�{B"����	kZ�&��r�)�68�ҊW�0�P�����bGJ���'\[��W�Fy�!�����C����}O4���'��TD��z`q�eVc+\,�����P�4�,�}`�>+��w+�%�cupŎg䟍
-ԏ�0P�x��'�����&U�S��rDw��i�UW��^{YN�{�8�ٹ70��b�8�����1e6�]�$���;�����e���'��*��[�)MO����vUM��º�F����r{-�yQ4��ꊋ����]}���?g����'�C��'�;�'�[�������F� �us������q�v�$cG�q�95�{���wJ%����we/	��ܛ�O�.�풝����~/��7��?{�y���VuUNn���S��b�r���!O\CE�'o���q�_�.ɋ���^��7G]�Ҁz���z5V��J�*���2�;�Ơ�7N�
�Ov�0���s����g]们�~]_���;��.�#���C�Ӟ�������?��6�����	՟�.����c�a�F�s4���|�,���1�h�����w��Ӯ���MS����y�1�WR���S���2�ºC�D �8��=��j�cVW�z����k�d�Ň�����f*^.G�ܮq�K�@��*H$y��֎��D�.{�i���WJN��C�)��/|���;�l���ьKp��ѱ��_�����s)�p�a��Gn[������u&�Jˣ�~}�*T��-�C���5�7�uB���0��[u<�-)J]��ݧy����v�ӯiW�� ��3�K雵wo��ыOi|������SP3@Aݰ�Ǟ�����1l�a����|�e+UG�@����1��LxL�P�G��lI�5q ��=�@�F2']������K�#��#l$������_�?�����)�`���y/�A�3��ɖ_f<�0���[�@B����{ʡ��^��ד�Y�)�h����%��i�̫/���+\'t�^���(Y4!!����Oc5�fV��Z����S�va�{=Ź����V����R���*oG������U�K��?�p�@Q�,KNM�]��J�v1)3V�B�VٿO+�$=�Q�y�@�� G{}bp�b�E��̗�Y`�՘�/��|wRMS�Z:�O#�]��@j8Ҥ�B��"v��ѭ��ԱjIP���p��@� �SyY�5��_-�ɠ��(�	#��2�4V�f�τ���BQ��f�k[�m���TjYNՆ�\GL�)�xa�W����D�2>B��R'/Q��`� �=���+��>�ۼ������Xm�f夢���N��I�v_��K�#(+n{�LT���`+����y��k�R��ǅe�~Y��$��GKs�Yj,�t�Rk;@Yu�ӏշ�4Z���
�:ޕZ����g�U&{�X�]�x9�*~&��M��dt�u� �C�4&����-���	��2��
���{�,�Ͼw|��tG���1�@3�.}�I�j֍�N^����F�K�d�z�K@�[�ND[F}y������7���	=E3��?�W���Di���X�j��Mo��"-��f;%o�8�����0�(��vD/�{�|�h�d���[�w(��Q�!�7��1w��lX#q��t�%��;�ѵ�k��]x�F�3�0�X��l5%{��̤��N)T�U�o���l�e���{0J�������[&��,6�}��KE��i��I=y��su���STf����Ք�ѓ�}N:�(b:��F��xĽ�ScʹB:� U�D��2g�Ju�WmpY-���z��f�%!?���������z���<6|E�zs:"��UU*A�^'[��ĵ���5_�`phЫ�(_�k�e���f�4�r�O�c�+�!�J���Q=G[7�������v?�S����f�fT�$y���,��E����1�ё��8k">��g����s�-L���sw�第��;�eO%U��~�z�WW� |6��f�m��=v�n�t�O�[�����ji��zn�X�8�{c�k$�I��������y?�iS��9���1At�,�jq��9m�]#-|�������G�Es�����Y�c��4��P����F�D�����6ݪV�|�AqK	�bߪ�[�.��,��pQ_?7��j����D�>�T�쫜��-K=<�ɼ�]l�V����z]!�Z]
+�	����@��q+لj�L9�3-
v�P�^F=s�5+
q�L��ܛ�D`r���L+YB��@����s%���� )_��Z`��z����RW�Zf�̫��G��IZ�p&��f��j>'�:YG�@TJ	*� ��|6�k��@�3 쮨,r��/?O1k��)5�<Ч���G����1�s9=N��_�)��Sr�����7�*3�ڄ+/�8䞦��v�G��<�R�Jl:5jIE�-a�J<�6�Qw�U2� P���X�$�Y�������Sw!�\�Z}�����d��uxG�xoA��{�v�϶�qᬾ�p�.`�-&�I�K���D��]�#���{�F�����v^���&�$<��e�#��rT�b������Ԅ�q���� ��J� ����:ֆ�������֩��}�,l2{,�'���'�m�^�]��_/�Zt.7/��&����R']5.��*o�տ0�<� ��vL�u^����x���۾�~u��������γ���@����.z�k߶sn<W���5f�C�e�ry۶�fޑ:/�p]-Ŵ���T�W�aۏ�o�Ź�Ʊ���6����ꢗq���0û@.##*s�{�0����'�\����MJ��	��hÔW�7'��n�K�zvo��ͼmN���W�;���� ���Ԙ�z���ִ*����C�����
q~[?}����2mj�XO�n�q��G�a�Y�k&�?�ܩXb��/� �?N�b]�i�K,}�(���t)F�K��C�����#�
��5f��-�Ԝ�B��ueAC!���tR�C��	�~OR�*su���yt/�{ �F>�HV74U��Fh�Y=�ɂ��3�h��Ƴq��g|%��*���za��c�S��_�Ǒs����0e'��-b�tf�F��ƞ�,��'��#E#2uԩ�G����)��.t�`r�dw�%;Sw'F'z�2:4Gb��1�=����Z2�t��k����a��2:<bFS�4��u=���h�� �	ϥH��.��>����97D'b$�ȥ���h �3a�L�
��.���9R$e,#T�6���U�M��I!�-�j��L֡�-����H!�l�+�3P�0p��TݣE�;8���H��3܇JvE_��d\��)x�M�C�Xگ�֨-;7�'�����V�h���hS����s�����ʠ�0ްTz�"����l�\$��[���:U�_�75-��}|���ST���~�0ȅ��f�Ç�(��K<2JmF���ۜs)P�TRvq�p����~�jx�'Ϸ;O,�v��J.�2��U�~���#�����lPDH�&{��\&����,@ӿ�zn	����iF_T��U���PT?���� �4E�f�1ů�B�U�,SN������"��Z�)LEY��rYj�[�!󅒭I4���/ʩ�	
Q��E�C�=`#e��uk�a����?r8�N:=8�����F��΁W�/$��h�4wuR�o�5�0F������.D��8dc2ҏo,%Y����]�P��B����d�6S�~��1Ť�V l�w�\bK��I�1)�$&I<}Q���q��U4�����)�IL���5��	��e�������8�B�� �D�OV�����8�Z��p��S+��{��-���JC��t:4�D�7m붦֔�N�]��Z��.ǔ!0�t#<����$U�8��OVTu�1��d�rX�r(���t�7��9uB<�sj&���E���h$X�53�Ę|�Q�F�(��0˪ρ����}m�┒_]��|����45c&H�25"p`�:�:?�j��jں�"[>�8��Iq���l	�jG�`�2єE9�
R�JO��� ���r�6S���J��,�֑
r�ZJ'r��l�8= �3Pnd�Z�)]z%�B3�d���Z8���N���45�g����&ŔI6ů��\h��#+3�0���rX��X>��9��a�.����'ht�k`J@�@�'J����?�)_�.�XS��M���7B� ���Z�*�J�Kho�M�d�(��4�@gJsX!�$pkg!������l�p�Т�9醦���&g�}R�-S�x��j��ynC�h��Fߦ緾.��N�֭����>1r�t�nrz����<}���[�:$�n~�}�k������{�>>����/�����[������~�{rn��+���&Z��ѹ�t�h��wЬ�-rNT� ��4��s�FY�����A> �!��lG��+dY�r�hd�S#�ھ��Se����ߨ:>G-W�(~�yܱ� �-v�'��c�1�QPEY0�itM��.�U>w���j���g���!�Zj�S8��6edc��ɭ��!"|��C��M'�߼
u��&�U�С�(�ĥwY�0B�V�^!{�#JY.B���q���j��6>NU�l����D%'bZLk�	d]q$4��jѩ��-��cd�P��ɇ��~�4EKncM%�UAB5�ҵ\�-�n5shR���6�O�?�z������ @L-J3��G��^x�'����hi"0~���0�����7i_0�V|ב��B�O�hzk�d#N��?P.YU�J?��(�k��������G!>�*�$��H�B�P�1�'�D�pk������������z�-�x��g5=���@zd�oG�*������jOguc��ek�-�G�����������P3B(���pbn;u�� �õ�2=�l��X�6v;�~�������f�������{\��y���=�{�~��I�G��������������+O��:=���~����ٟ?�λ�^�?8���x���O�~��=r����~ݻ=�wx{t����S�T�����nO�X�����*�wx�w{�V) _4k�|K�ړu�NN�������we��@o�}��FuKpR]������3���'?o����&�Ǖ�g�?�=�E��nW3����7w���������w���{���O?��}���O?�[�|~z�_�j̞��9����C�=#
i�q��M'����/�	g٦IA�#Α�A5�I�N8%� 8��"G��������V��"�r��7&�uUQ��FQj��3!��7��*@�4]��pl��ҿ��#�h�M7Z&ʊ`�昺�;�����y4���k�?p+�K��:GcP���r��T-�����1�)�)ԧ%���ѐ[�Q'h8Bv@�yP��ɪ���#��h=�@�=U���)|}"p6�zؕ����7#ޢJ�`j���%�Ƅ(�L�=N��(��n��R35��(�B8��r�g��1�-k6a�ɕ�Y�h�|�FL�h��q�Ǉ�\�J��,jƶAJ����%�!|�rӉ�3���aBE��!R��#��+dB�+�z!�5FR	2��� HD�8���1�3!�����Kta�qL��)��W�v��B�yZ�OS��'{K��m;̗[��M
��ْ�ʯ̔u%��"��I�ţr�)�"ҌDK�����b6�Ԥܔ�[����M�@�6�
p�\1M���c+2�=����ъD����*Ǒ%ŉ'�t:�u
!�x��ku
)���q����J�(�SQ"���,Rє	IW4�*�S�Y��(�,�im�{�嗾�/}��ZR���t#&��G+ǓH~K�D/*Q�SȔ_!2|������mYR��y ��D`���Z~!QR�Ϻ�A�M���t̮:�1;�qzM����NB)F#��pDJ�w���J�o�$�h�d	�~O�B�h�"�d|�B8U�>�|��9�r[W!k�-�� �p)C�W�9�I��>��8��0&�����p�RJ82���lw�R�M$�y(AN�!ĉ_?F"�f6��ŴZ86���^\�� �1Ӈ �!� �$lEtphZD9�1��t���q*������KQ�3���g�VV��)NjƘ!t�ɂ��k8��*�(fQc`��c��쿊��l{.=�m�����4q8��哕Hߘ�Ϟ���*�I�J��%��/�So�끏��8dR��8�6&E��r��B�|�8@|cLxGP�%���h"��j�)�&:U�R��A�e�b�qL�(_�F��k�;ą0ME����;ibՀSxR��L�\������eCŷ��6��.jl�R0���9?˝f�^*�`"�9��a��3B�6�.������~�z�+�Q|��q��T�)ZV��-��vw�V�R�[N�1e:B�z�ɦ�cGAn�$����y�VQ�RpX}6b2�q������L���u��2V���ԺL�g�"Tw�L�U1��E�P���*���k�� >&�n����P9U�¡ ��7
q<�"G3�U�#W4�,Y!��k�Ҧv�f뒫��᫒�*3g�b$�VSQ�F�`�u��R|����B�g��?f�7!����b�'���C�E�7y��1� 
|�;���;�k~��O}��*:oN�0�3=^x��n�w�M?�{n�V���7=�P������֦?�����\���m����lȁo~�����@���V���x���;�JX�����p��;����^��Z�T�:S��؆����E�n��Ç�U9dY@
�q"$��"�����g�R���E�R0��������u���m����-�^�cJA��ɺv��d�n��!A"8D8���(�T:�,��4�N4f��Bl    IDAT��_	�&�"r��R�k�*FQ+���h|���p�2
I�.Dajq,6d����9��Äs*TES=$/d$�rmP��V�������Tz��x�S���q"�UC�:�ϑ�<��Hc����J��'U
q ~Τ �8�D��K�b�8RJ'(����.D����S����2>m��3�[޺/
G�(7����8��(�P�Iu!B�9F����R�[��1���7��M��q=��P���p�j�h��R*��էl�?�Ԟ�ՏQ���4����i��ґ˂s�W�g�,���hR0zl������
�h,�YLH�� o^�rY�7� �=#x���k�.�c���5�}k��tD	Q�VOZ�OT���tӒp��T�h��:!�ҁ��`ʝt��6ي8��vܿ�Y��gO{��}q|	���e�ώ�7�3����w����ڈk?Oy�M�+�mpe۴�h^\<9�;xpz���֛��:ʾ��G��o�����������l]=�^�㯿����cݿ!��|��f�$�oZ�f�'����w��\�y�]�W�{/�;�ۋs+�½�<?�^�7]O��=y�?gb���E��YO��۳�Oh\޺���>�':|)����]ք75�^Pi�#����g_�==����oN<���k���_q��+_y���o=�����/������ӳ���ۯ�>q�qz�F^���(�s��˂N>8�a����"��6�tp9w����݋���eE9s�HT(Yj�9!Vh����w"�KRE�S�4Lx�4ME-��Tc�:ėn'�c:R(���:�X�QY��O��r�:竈�K�ɢ���A��HEsu�m�\
�5u�=�B�(��nD�F�f<iH����">|ՙN 	N�-�>��\�\��pY���S�_c������p
|�\; ��V�LY�Y��Q��������,�G�闎�_G�/�� �L!p)�
�R�!Xu �,�P�T��ZBQ�����'���Aj�ϱ	�D��*|!�V�-V
�%U�\L'���b�%��lL�NH�������v�V(f�ݬ���12
�$�p�-S�S���ř,d�3��d��kO(9Z����LSם��3�?K��F�	��4�.��呿m�_��|� ���(��T�5�#�7�=bxU��:�[��$���H�g����I��`-�jjġ�p:3S�_��cm������k�TW���iOUZj(�{�BS��c�%�dS"h�L�i������J�[���mH|u�LK�?�<5|RrS�C��rHQ�>��%ȡ�����&Pu�H�����"]�t|G�!�o�8���� ;cZ�LG�3�*}�%R&��,%r"cr�Fm�f� \�%��C-r���R���g4|Q����Z�B�'\������,2Y-�;��T!!-AX}r��
U2U�eQ�W�2f��6D[H�I����q,�&�hC�#�LR#��
��T�%bJ�_�DNGǢ�"�>f���W���1ф-������ۢ(�,����i"ۊ��� �NS4K��l�4�@!"�(ה��t�4���V�Z�p�"[�r) ��I����O�)��*�aN �Цt��	drc�{P-��B�[�:$�I���*�aƑ���.�48|u�B�e����ILPir�4�C&T��Y)Swd��Ʃ��v���B���RV7eM�'�n��&(��\]��rE����k��ʹB
����z��8�!�d՘N�o8���c:�,��mg�(�:ϩ�!c6����˜M��m�`��Bp8hm��1��d�e��R�R�B�B���ɾ��.2S�U��aŬ#Z�|���E�ޅ�4��6�uD�pQ��,#�AvO���|N��N�U>)�lc��gh�%1m�F:S�%Y�U��
���r��X�CO9�-�-��z-�-E)w�d���d2!)�pBG?��i�s��,M�g������!.%���j1�5`O�Fnj��_bcj�Uxۢ�FQ���Z;��*j��	������P@�����T�e�[�3�r�8S}���]j�\��Ԍ�3A����FN������Z)!�F�@L������Q��]µW9.�+od{���(�Z�S	�U]�N &����rE��e��_i���nzֵ���\����_�ꛇ��O�8�7��έR7�v�ޏ<<���7'�G��F��ݭ�{�}Kg�Os�fo<8�`����W�z[t�������?���O�k}{������k/����T�����qK�.�����=w�D�鶱�?+� _�i����40v}Y���uz�ьd�U�l�_�߶ehF"(Hm���6�� �Q�PUwc��9��BY�!8�@u��D"�I���?8J#�� ���@S�t�ɷ���b�5��g|W�\�(��VnQ�]�\��Mc
�6D�h�uE�P��Euk��E�?妁�uh�4ߨ���0MKD㳤*�"daF�d�
*Q{k:Q��B0��_��L�ZSejE���K�8��	M�ɍ0�����2���.`E�4M3j��r���t\�Zr��4��=##���Ӊ��5�J"�B���iF�(�Pj��B��"f#C�9k1�S?��~����V�3��_�ҝy�@���<�J'n�]�����̧O����㳢U��Z-W�_3!ӤPu��3���ݙ��߆p\���F��BU���^��*ڨ��s��%���N�Ep�����1�{n@y����O��{��O��O�#�<�w~�TU�������i�m�, �բΨ�0�X$N-J�GT��|����f��J�����i�Ӧ��K�K����zw���O֍��Ǉ#�������ߤ>�9�qKv�=�w�.���{7��~�ß������~�ӓ7��I���������?|q�����'~�Z�O��u<��}�]�1��奝���1JGa��������G-.u��M�l����W�j�?yrFy��m&���ީ�v�zu�x{ԗ��YP3��꾷R��ozC�z=4<z{��ÔN<�;�
���������ϟ<{�3�ׯ�郛��G��G����wο�އO���;o�����/߹}�����gg�aԓ��l��:#���E�n'9(�]5�xr�tg��h2:�N���if!�>�sKA�t��e�'2'	�ϊ6%�A����w�dʌ�[g��ƩU�(�s��eE��>u޺R��k�
g��&�>|��S�
�6M��rHI䐲�vU
���D��!8t$
��tdYAˑ¤t.�}�[>�E�:G�u_�C�Ç
[�Ǒ�FYu�:�>5� �M�pSU��9_
k����KiF�lYF)��Wf�8@F�,�0�&u^�\>B#G]���B[�#^.���@d�S�r9�L�Ժ���^�+W�ȩQ�@�)כD �(�k@z
�56�rd�Ҁ�G�BM�N!�1�_"�ϐ;�����
!��|��Y�UT�V�s��qF!�)���Ukl��E��hWM�(+\d&�o���4N8G����V�4B��A�U1ʭ��0���\�D�D#Onw	�.T�'0�b���ȷ��B�{r�F"�Δ?R�Ί૿�K��u����|��+Ż�RLEM�����B-#^�i���pX�)N}�W-|DFت�AJǈ�\��wwJ#xԊ&ʡc	����=��Uik��Q���2���};+��5fJP�Ad%�E9p~��#.8GH�"��#��o�|:����@"9UdhJ@�|d#q!�9+����R6�U��IQ��Ɣ� M���#�#��CL���q�W�*j���2��M�6��z�u�IV�CB�q�1!�t�����i7�k���NV¶9-_3�"�6q�oi�@�����%lK��h��t��@QF.������Zd�GE��r����a�M�2FF��X"��Q�-��ԤhS|4
h4�CkC�p ̬,����Bh:��c7r�B��G�s(C�Hap
EKojdp�p�\	`jRM!{"J�c��c����G�`��"7}��i[K����s����`�ũ���De�k�TӲL�,��n�'�����(��j�(� 25�)>A%l>�-���` (����ڣ W��5��e����[���M��-Ĕ&DH"���H%(
gd�zb�#����eEkE�"�F�� g���VѨs�{xa>?��0�IL����6�q�G�4j�_�8S>>\"�耳9�f�/�Z|G���P�LY�Ȗ�		W�od�d#2�ض9	��ܔ>X!N����,r%LKO�i]���3r!m �@#�A"*
��0�����J~�ڌ>��sF� I	! ���O��G�X'B��Vᲀ��9B8�c	�IIP0_:���D0� ���Mo���Ei�����RL�T�X'5�ﱫ�	Q:�\6�E�#R����
�q�8��)��iȌ����R��B� �2�Y�u���I�pQ���u%n3�$;%�����ӇH	�P���x;FE�9��D�I����D.�֎�I�DLN�먩>!�[����(��Lݦ1[5��pڷq�@���������ᚸ�Jh�VSN�T�Ü�_!#eB���2T��Q�q��c�6StL���8��
qz^�K1_�Gm��|�r�OO�����4�;��rL�/h�B>nyy���'��/�r���Y�l^�\��Ѽ=�;����6�/�[�d<9{���C7S}��>�yz���|��g2/��]�>�ys�͗�������{����_[�|=���뵟���u�v����nz��N���{߾��3�5b�֡�w! 5ә@��ֶؙp+�������m�Q!�(�Sfjt���"��wnȵLcLY|4�T�hʑ�p��J!���dlKj5VW��	F�"q!)8��"�̨�`��@#���F�h��D0���C!Vi�P.+�^u4Eٖ���$�\QU��eq�"$�_{�%���@�	):u���D��P9H"�i�f:j|�F�(sƄ��ft���Q@A�Y���q��5	d���y~E�R�E��2�NW���K9k_�E��ͦ(f�]���Uu>�5r�fu���8)h*�4SV��fcG�n���JdJ���wR!3��F>2�3��S��G0�����PE#�o�.�B@�׹��)C3���U_���aN�
��{U߸�P�V3�#Z�ܲ����v^�|�Hi�I����Q{�ާ&��/��䷛I��&�'�|�O�GH�?��c���o���	�����Q��I�M@Fq��B��ZR�r��uȣ9.~ s�|������
���2���FD��_k�>�����9����YM?(��Y�� �uy��)�0{�9�����#�G>x��x���|�������O~����s���ŗ_��7_���_���y'�=�C?Z�K���^{>�+�N�o�y�yg�J� �_oI�{�����P�ގDs��^כ� ���v��>^���gv�{��G9���}����A��}N�w�nR>xz{s~�k���'�u���n"n���N�ۛ�~���������g���?�=x��7������~�����/>����y���]}����'GǷ2�n��;&z[/q|����W��q :5�9�*���� bG����:��8p"��M�S%��k��s��̤�A��k/��B|L�8��E�X�2|������5# )�XTq��+*d!/���"nڹM!Y�Q���s�E���V˽%84�r]z�H?)m@��8��e���D�1�z@I�M1鋺[�l�H�=LԉMփ��G���JT�&��6�Yw($2���xxB�	� �>���� ��Q��,M���y� �P!R�$rN��i45fu��	)'WV�88t�N�mh��Ki9�1|}Jou�R:'�l����:nLʈ ��p�oԌ�m�7��(�(���� P锍��!�KI�X?�E���� �'�fD'����[{����-��R��9��p�B�U���?����;��*�n�(�"p��GD��Ȋ?Zj�i��k�	1�O��K��a������)��߯�J�.���L�j��"�h�U^g)Y��q����IYT'O~��L!�>��iƬI�(��aL{L����S���6���:��S��W.e)n�$E4�S�
��K�NV�WD���0�Ɩ�aȦ���90�P�5)$=���F��sG���_�J�'�4IDW�Hy��N�6�)����,��*%�En��B�"��5	Af-9g#�A	�����2KgR�f�
Y��hJ���b+82m T�öR���aȔs������#=԰��#����݋gN����|���<w;0+Ԋ*���I�?Scr���À��L�p�W�٪��T�*�gD��	g��p�]/r!�R����g=�*/�t⪘�|���]1>&ȑQ����BЛB)�2Scmp�(W?=�u�0KB&h����R'�6A.02GWF��D)p2�,��]�D�Y�$+]"rʢ�`�t�0�����i-^� ���.#B�(s��6A9��l8dS�m	8�lr�7�O>5����D�LW�,��D���r3�ʅۍ^�I��?�9d\]4�W���@��mG�*�!dwߊ���
��5F�(DnG�%��:�8�u������K������BxШ�tb�,K.ДS��GP�m}Nj��-�.)�pd�J�'�&&И>r-�&.�N]��O��d�p��i�t�|x-�F��(�fLPJ�K�I��W��+4#D�1re�+]�td�[��q�r�қh[]"�nQQv��!�Y:����q
U��8�D9N�l��KVLF�q"�)o�ڢ�G��J/�vq��J(�D��0U� �su)�rf���y���N��Sј8��#9>�TQ�tc
IN:Y+����0����p�L��i`:Gf�����T���B�Q�,�RŘN��q�XLј�yWG�LkCJ�M���e�X'U��/:Nm���0�ii�()�:#�i�rmhՔo̧S?r���	��a�?x���W��-2�%��LS'���f���aj3L~!��pG���Ə��֥��ĶKE|fJJ
$_.G�ɪ=���*
GpL�M�X��G�s�ʷ�8C�X�syu���[����xW���e|����B7>�aβ�g��oΗ�_��ɼ9J��op�1N�D�zpq~qr���wʝ=���N�//��y��k�4��={��ٳ'z��m/����<E*���5��/&f�N�Ķ��.��2�Id'&Gh7˔�I�,�\H�ND(qx�ɚJ�:��S���VJǗ_VG����½�2jC?�p!j�8S��a����u�'Bui��R#�J�j��L��T�V.K(�"4%^:L8�@~�F\�fz�����h���r�7��T�BL#��-r>|�^��pfs��0/��uLߔ���h>��RR��-}8�:��Z��$N.�vM��FH�>{I�&��t�e4�Lவ|"NN�ȝ�mW)�v�A�2B�jw� 5_(��~Z��\�(��0�:��QKr�c!p�F!N�8����h���.���]I��U�V]��#_�lӸۖt Z2�EP�F!d#�ьP]����4�-����f��d��ЦC�D������Ѻ�����b����5Խ���[ �;�n���7���mˇ~HB�)G>]VI��_���Y�������}���.HƔ�!�c��*�����[��G�*�y��1`��BG�rtn���\߽m%�xj�����s�ի����홬Vꬣ��#j�C��~�֢ӁDL 嶀϶x�#�����k\ώ��.��"��D�<>��o�lv�>b�7n^������/��;��5	7������������Κ�'ϟ|����>��g��+�s��_֝EUn�o�|�^z>���U���+}����N/�}���ğ� �*���F;g����au����7�^�[6��6�{���Eͧ9���޸�q}��̰���C�Ba���aC�w��$�����y�c���^\?����8��£�|����ٽ>�����W^{�o|�����S�L    IDAT��Ǜ룟��o=~���������ӛ��u>m��S���޾N�@��ߙ�8�@���S�s�A7E��-3Ċ�<N	Y=��l�Ā�J�9�OS�\
�Nn�|]I�;i���h��tZ�hu9RHq0�F�������h�T�	)d����B���q����T$2:h|/�q8E-�c55"@�
8�$M!��r�z�`�����=5L��d�k"�)Ga���O��Ap�PBu>G
m�,>AK�h�M�!���m�����j�mSj���PFPW�Z
euR�1���J8qw�d��i��ۦB�a��*
lQ8L��
�.D�`
�Ҟ�4���ե�K�e����E5c��m�-�@ԊP�*��\:�1&��r�3ܨ�1M̢�(�*7`��Z��������OA��W�5&ďYn�R ��nM��.��b�~Q���a�p��rY��L��f�O��\:��i���ScF�g5>��RW�)=4D��z���d!�[rK B��H���H���ݤ����;iK'N�K)�m�L���r��� �n�éI4�~l�tc�C�T�/��R4�T�a�8�6��	�����Ҝ��Ebj���`�4Bpt��jD�[�U�r�F�����kj[R�$��(_zG�(&ı��D�D�|�ќ6�S!E?KG���i2>�T���	�P6���E��MK�4���-8uHmS]�o�u�O͔�dh91��-�J͘cRh�fڶ�i^�kk�Z���tN������9������ӐϭzXy���a�y-Ŝ���8Vǀ�g���f�o��`�����xT���;|�UQ�舸@�Ѩխ�ï(B�,�S-R,Y��t��@�u�&Ժ�v��e�J1�ρ�`�g|}*!���!B��7F�U!F֔��@�d�@m����^�Rf|�(�U{e�4�����o��������d��W�1M+A��-��L��4�H�n�LSc^�������!�K'��x[Y��OM��"Y��I�jg��(<��\x!YSYH9c���rj�S"Z�jAte!���)W(����k�',�BPnS�׉1Y��\��x���k�
Vif�5�f:)��uqlf���QOy���DeY��"�d�� �v�2YtZB�3"&�05&Et��]?ۨBJW]b���KL�c-q���LGȞ��q��Șօ�"7��Q��_�)PTR��|�9�ӏ)}d��ڔ��z���iK�L[EYF�ҕ*1��� !�2�_'�Y��|�X��R�O��H�Ko�����0�@<ґ�gR�<j:j�@�䚦o'9�.���؄eUWV�֒㗋�"@�a�pcu	Z�i!S"M��b�2�:ߌ��"pDS3�.�JޮB�R�8h���Ι��8�p&W]�!��t�r(�̎E�UW.��KoQjn+�Z��j]�2Y�^�:1�z�� 5Sπ|{w40��8lj|�����J�N��w`��k��SV4 r"���L��U���2��"�!�����@���M34�0x��I�9�i{�Y��b�.��.Յ�ƬR��V�z������;)��$w}a�ŕ���9��w��.u��]��4���N��ϊ��b�Ovz;��3�:���o(�9�Bͷٹqy���c�豏���������_|�Oz�Wׂٚ]�|/�=E�ƶ��+���q����0��%K�n�z1n��>D�lۓ�V)t |��L��+a�	��_�F������� g��4!8L��v�o��Ŝ��LkIu�t)mE�G�V��j&�3YJu�pDzUrZ?�d���FM���c�@��SK��EYH����o�V_:>���JT�t�hL;� 
a�	A�m��1���d8x�Oٴ�:�	�	O��M�?��"ę}H3�̱��_h�l��3'sMj�*�.����i�1Gs���|K9B�֒�]��qf
�nʑ�1٦5��T�b2�qD�-�)َ��Ԏ���C��S)�e�j#�(řL��!9�%�#�a@&����:����	! �(�e��m���9��zz�5�%"�~R9@!�ik��X]�h����E�J�F�)2����Z���o~�_��7.����g�g�|��?��Ϗ~��_y
����w�}�Uu�x���:[B
�v�
n%�"���6�iU!hl���z��9w�(�������_����!V�a�6�Ӟ��Ã�}�\������ӣu����ց�T�)�{�.���sF:�ׯ�����������|��^�\?=��Ӈ����O�/���ﶠ5������������.|�q�N�k���m���������`!�Z�^"����(��.~�s}ԋ�sS%3w9��p�U�=�Ud{�W��w��F���	�uh�9��'��Ce�ZX\�[�p���2����>�xv��ѧg/�~������>8>�{�W�>��񣇿������=z�ٗ�?��S���Z���[-�>�v�-Ku�N�F4g�p�3�ܶ�k�����IIS�tN�i �����8����<�@N�?��BH�H\��8�a��n-�L�:o�A6"3��THTJ��B�"�4�n7R�@?'ૡ-�[��ɪ�CV�|��=v,t"�㑏#�����+W31�SP�6������J�(ܵ�z9F�N��8R�T->u�7,�))Ũ��s��5�i&�p�u[Ð��Xf�V��CΩg��:��0���`n�B��vO�)��_G��� �**ݾ��>Rz#n���(DV�1>S
B4Á8��jfj�L3_↭3��)��82#��,4=h#�Q"M�h��!��!���Z_J
��bVB�`��<�qHq��K��BJ'e�x��Th:���8��&�,8&�V�:j�Y�V�2%��U|���5R= !8|L�N]��S���ܪtR�R����§��t��V�%���Mȧ��nu&�UH��q�-��#�C
��m3��w�j��f�V%��a�D�i�R8F��,��Ar�Lm#�~LG?@"Ȕ>�BD�|NK3���T�B�@���
-�X�Uf�t�rk "}���5�&��� ~}�1Uij	i"8��� �R�(^�BRK��I<�������s��0����mN[�C�W=d��|�L��qN>���M3ʢ\	E9�d��i��.�Z;fR����D�����4�
�ʣσ���,�h�Vg�,w��i+��nK0Ŝ���6g�>-��A9'�1�!�q	W"�%{m��8����'��J#!����tK�od�mB�]�8�i��&r��j���~����#bQ%�-_:�h����
\���D�ƚvF�I5�!reu4����xq���f�ISQ�֘,����Z��ht���e�� �+!������V�*zM�F�(Ħ�o��b��fV�>)˂��Q>�N )|#��`�rD{�h���m�ir�B����Ә�i�D0�^��r�v�ʶU�����f���*�����E��!��i�ρ3E1�Ooq�"��7/�#xfw�'+5����r���4VBH��׉�#ԧ�����8�W+Y>b����
h�v�6B�t�����2�/W��U9�f���uP6���S
!qY�����p��6����$ed���d�*��浔x�+aL�9P�N	!ӡIǁp�̘>�B�0+d�tU �2�ja24ȴ�IV�C AҪ�bڄ*Ƈ���a*�q:�q�� Xi�s�(=)8ed�f�MS�č�D*T����L!d��Br���{��F��^=�9,�i�D#_V�2�"�c�W�D8GK��U�o���ʵ��	����@�j��*Wt6�)���S�ϐ��"�t�n@z��%�1t�a���.S�.��i��V���AO"*�GA�U�ԉR�G�"�5JDp�T�«g��UT"B_�h@�X	!�p�!Ԍ���B�?�R�������#)�>X�\��%���!E�['KlC�x�Tօ7<E����m���7պ�����~���h�{w�ۦ����8�������	P"�N��;����������I��j�.�[��y^�c{S��O؟��ç��g��H���:����c�Y;[����ӣ�1n��Gmj]m�!�mn���Ur�vKB���qd>�rI�?�B�H�pT��`ę��4�.D���V�J�ɢ	�7J��_(�����)'MN�}��#$%T	`4
B�F�6�1�k!ddM92K|h+%"�%�V�R�pL&m�~"s���5�ˍ�r���Lc�qL��F���ᵭDN퉶^��)��.Mn�V!�rYc�
Fj!�뿆Kn�W�+!:�i�H�r9��eA|}���G�LK�BFHk�7��~;���O�h�r��4w�_]EK7E6��O�)�����U׈��?R��N4�)#.�>_�.����8959͔^�Qh��=QκhB���\H dZ�/M�A��aV� ��
��{^��/~�_���K^O����BP»���q}�ȟ��w�'	��Q�
	�*��n�y�Z(Z	CC��ҍj BL��TQV�D�~9s���'H{�Iφ��ڽ�ח���w�":m�N]%��=����Խ�Ã��8��No�^~��{��E{���/��ɏ~���~�����	�ӏ>�Ⓩ�>�mO�>p��[�v '@ؿX'��|��=,Ǉ#q���Z���GW���W�3��xշ���x���H�,1��״�(Zk�:'��w��y��q*o��<��L�}s-u���ﶵ��#�b{��p^_9�<�h��#��<�|m���s7U}�ΗA��)�&�����'��'ϟ}� �^|p����ۿ��ӏ~�~�����{����|�/�8�~���k��W�ud;���m;�ޑ��+H4'D�?p�s#�&�.�M+An���A�1 ��t�6�z$��XV:uB���Z�9,ҙY9�^		U����-'�0�;K "d��-�C�ZRF��u�מ�^
E�<:z�����x�"ݣն0)Z���Jc���=69�%��1���_EL_W����(��)��V)�J�TS4�%�U��h	EM-_"�Z)�)׹�M��Dpd�@8?qH��5��3L�tB�>pL[BYY��y)��`�0MLM����|d4#_�Z�\�D�S�_�B�B�M	җ�zqY����[�Ddq�f*�A�FF���VN4S魷uUb��ȚEQRCk[�^�tpL-�6�Y����Dp��Q##���� 4���1��wG|�I�3
�R*d�Fq�n1�N>#�i��w����m��م��/��N���Yi+��nϭθ�o�+����8<4����N"`�*:�8�V��VWFR���BM+=�@Q�|ʥ@Z��491�=T!V��(��y��A�6��E�[�Ʃ%K�Dn]�5y��"X�-�(MVQ����T��R�_c���#q����(�a)�@��2NB�@�C�t�hM�B��"�`v��-��Q��VW@�h�&2+2��@4N� s䲔�I�	-Ŕ�tHgv"!(���a�����Xȩs~�)��%�|��ۣ��P���M�<�c&�P�)�I�Sz���\>���s�阶^N�+�Qu�������m}�2�r���4!m��A��䰲�¯�HG�i�����O!>�3R��6&+1����/E9���զǑ���	�{�B�52`�F���(|�s{�d�� "���?��D(3�'��:�̙ff�G �JL4|!��QF�1��(�W�ӫe�'�K���7�k2dm�}���iK�%���Iy�i�Ƥ$��r홪k,7�c	
)��N��/4�*���d5�
}T(�T��b��d#Yi
B�Dc�ɵ����-2����C�%��M�핐i/tR�O���`d��
� ���P���J�-�ʵ�H�(���L���$J�;F4��N�ޓ�JP畓a�ơ�1��ʝM��L��ȐY���ل� �\V��j!��Va���PSȴ*BD�8��p ��@|�Cci��`�_Tc�T1M�D#ZQ~�(�f8*�E��:��L���DpZQˑ��S(Zjp&W��T�N,GHʬK�_8���2��.ȇ��k�n�l/�� �'2B�k�qFMz'v�B,���
�h���3N��k/�t�"�)�Q��Vm�٢�LC�8
q�8d%0q��օ��|%��6�����R>�;g*Q�Y���&d$��5%�M~�wB�Rn��ԕ<���w��0LW�-�]��r
qf9��4E6�jC��)�n��q"p �6s��,�A�KG.�(G��j/>�h�
�%�ȋy��.�{�ױ�G(��Dj>���Q��f��Ѭ�մwC��y��u�>����CQ���'���Ϸ?�Y��^�^9���'W~1Loh~����^�)��ý�Ϯ\���<��\�ޞV�����up[Z��9��2�q���tpm�o�5u:�3K���+�{��kaw��S"�P���"����|ۅdIiIQS��fn�G�dM��`!�A^�ͩmd��E�C��>ќ �A0��ZJM�6)���ĥ���e��E� �M�|��ʅ��#�� J�c$��TH�U�2�3���U�j�D�zxS>+%��lo��i����qD�U��]Յpf��8���43�U7�ȒbC�7�ߊ��dw�ۧ��)G�O�1�Z{n:�I4�F��?R�TI5JY~�,�<�e�ɯI����0&�.X
��ե���>wS�ZN�z�kʗ�FAi�#d,���Q����c��Nc�J�d�2_!���v	�fd�Y���EKW�3��O9�Vd�:��M������ �~���TT�}���e�ڽi�1"��?�����f������K(�|��_��m	w71�n��ڔVn�咖zz2�P�����������e�>�{����������{k�s���M�����:��oL:�>�y�yx`y2��ϟ��]>8�>��8=�{�����7�|��?~��?z��o����}��/?�䳇y��7�n$����ݑ�<[����tt;�ʗ��5죛�?|}y���|�l��Y��=�ۀu����'m�p�+r�¦������%��ܞ]\H�.˰	K��g����K��F��������	V���A��0�Ow���}/8�sI��Y�`}Iģ/���������ų��c(�txsv����qt���/<x�O����/}|�����}7K?~�����7�*zu�-��{-���ft��������[�!�;gMS�R�,��m��,���4%��5e�^}R��|U��*��^�B@��=B��q23o���W�AL�&���o|�c	����(i�C�C�~o���nmFV��Dj[<�5$�Җ&+���`B8��(�'��jO��6�M�����A�+���?h������>�)�qD�XW�Ն)}#�Fd̢�M�l]�Wf�-ʪ1)-��d ��ʗ��ZT}J�5euB!�>7�퓇6\!m�#+���b)�J�M�Y&<A�m5~�a*-k�t���v�b�`���kiR�R��g4��S!�rtNE����0�9mN� Ui�*�Y�8��Rxd ��v�*h�1��8@QSݶަ�b���Yk�᧖S9d&j:HdG"�i�ik�TF�����,L�1r��9�Ff�@��R�p!����z˟#QH�ۺ9�.J�N�v�_-�qj8@���K�ҍ@Q�d:eķ	��.����1��b+ѾYf�YS���s�I�B@>�u�1�z尖f�B��~�&(%��OJ�h _�Q��!9�jTqh��RNJ���� P��'H?AS'�,�,T?�T��i�����2�M���;���J�)�zv�7���O�G"�X�Is�4m�0)����۝�k,�QS.�S?u"��ߴ&M�ijcd�3�@R%%�v�@~g�5�o�b�
OM
�CĈF���.�Z��Eq��1�/88�,�d�8,���M�2�\>G(�ߪM7���-�U�S%�!��L#�����e4m���    IDATr��/©y�1�L.rRU7�����Ɵ���̓`)!8V�Ju��g9B]�٘r�c����t���Q�5̐��3R��i��+Dg�W��g�9��)��䋚zM赢狲_��Ѫ��a�J�R)F
�Mj�|�uƑ"�3S���Mer�,��
'P���mE1E�I���C1v@��E�+���)+�h�����!���]�b)����HI��ɉ� ��IyZ�w,�e���
���4KA0�V9#�B�,Q
��p|9U���m��ޖЍa!�/}m����d;"B��ǔE
M���j�X���ӡő_�M"}jF#<&���D��BY�	42 ��|Ȉ�2���҈I>"����Q@nϧO�
Qk���, 5S#�5Xt�Q�iF�a�_fJ�����;2Bm�9��8u�d!pVi#�q� ���0q�ćb2j)�M��"k��� j`
9��S!��@�*@�:�C\9�,&<#�� qV����?0E�J�cZ"����B��]5~Ew{@6e�L
3��<BmS����B탖(�2Nd�1i΢��
N�jb;�UDf��mcq8�d��|�-�z�U��[H����ա��I�C��td����nE��B���a��[q�X��,��]��B�R�)C�Q��wĪE�G+�l���R�[��[���V�i��}�B�:]���މ��_�懰�R���>=9���������k�;��U�AUZ���)�Պ�ey@a�zoҏ�=�q�8:;�|�cn���{�_>y���֖��6�Μ���� ,�q����߻ޢ��s���<�v[M*Z�Z�V����sL��t 8�|"���]}�V��hm{jdME�`� _W��1���
a�(�($?5���N-3�t(�w����
��G�?S�-B��X"�N��I�>C�c�N��ӳ�C��)�OAh�54e5S��|��2�w�	��B6��mSN���4�5>dQxj� DL�59��!�)��P����U"&��hj�cLc=�ЉSzY�����^��
IǙ�Z�i��X���0�Ƣ��p M)�`d�����kF'qꜯQN����&��"r��3��m�f�)H�Q���S6��B1�Tj�.Pr��\���� NRi�
�On��X�4)Iq��j�y�e��Q�T��A25c/̺\H$.���[0p�����FW{�#�y�Y���{�����<�d���N����y����EugM�T�l=-5�=����Ks�LW%A�sȊ��.=]q֏\�i7O�^�m��Z��C�i��M<���ܽ����?����߹�9����?~�V���U����z�Ñ���}8q}`S	���H��=��$��vGѡpJ������7�Zݻ��	���M�E������F7h}o��	Ԗ�zr^���D���.JV-�/�g}q��O�3��a�on�;��խ����P�^�ĵ��J�?��������}w�����4�q�g�ݷkkm)��{�O�|���K�}��������'���G?��x���_�����������/�>�MO�ᵝ�}�����r���juk!���Z��ѹ��0vċ�Hޖ�6��:t[��P.�gy��,2��%8��S�n�KA����)�i�d�]��-!�NJ�/WV�qS���0PZ:?P	R�s�I��,���H��YQ���DH�'˱R~���h����h�J]A<��p���\;�#�wYP����}���=4U]]�ZUE����H�iU�+�f1�TBTuQ��ǈ�yR�:WZ�>'��bф,�\Rr!V�f�%$�Б���W����_��n������eh�Ԩ����[n:K�'�:@SY��~�R,D�B��PcFRU4�b@&��`|�r��M4A%�->f����T�IdhF�V��6x������k��-��,ZѢ|��i�IV4>�%�G�oL�H�Q�4�Q'v��mAc�D#k�Cp�4C����K9Ļ'�aft�8���&�t�! =p����\ɨ�+ �y���BD	��	��ٸkP׈OGi�����-����d�S̮�B��f�4ʅ��*T�8AK�_�pS>>�@����(-T��8p�E6�k�T�#�9[��I����A(��Ф�t�������"�B�3^���E[)d)��o�p>���X`:�������s�K��[,�\�-�z�+Mz��g�U��O�HN{R.��"�� ��I�B��I�Ȋrʍ��2#�ң�N{�B��
k�c�ѲD��G�Ko�)>)d�v�f��tXQ �T�]
d6J@D��sG��JL{U2��B��F`�pv��׻F!�Kl���߸/�1��pX��j��7��-��	NnUR"B<�MV��������)��|�֒B���jն1�q�Q���F0�KI��4�E�ΛR�D02���� �/�Y�k�U�=�8m<AD��:T"NOD��v�{��qL�uHܴ%�����Q6��o�x:��@�dH��~�e�9��ar�)Tw�ˢ�k	�I1��·�1��egW������g�F֪����@$��Ϧ�U+���`r�7�o�?��dq؜9Ȧ��؇�;#���c������tr m,B{�q��/�9���iƬ�Fі �<�|6EÛs�YdRV:>�>�� 盶j�i@4�P��SۣP����h)�����}V����L4�i�� d��qLe�7����o�ɪ.2>+:m��[�(�MHSH��X� 
����@�
�bԢ���O��ь�K�r�E�O�h�Q̈́(�a�쀺-G(�b�,��ĥ`j[c�t^�	Fd�R0�_�ܝ���.M܊��>�jfpV
��6��q]�)�_'eS>�2�pD��Ԑ�5F :�ۓ�ӯ�Y�S���}馔q�F.QW���J���ӯ:`Q���rk B�8SMÏ��?rR�V�JG�/�R��>K!I�=G���?=X}J�'��=4�Z����5��R�#/q������}��hZ��]��z�ѷ���ҡ�9O)�j���'�g���:7A��n������}�6�=��	��W_y�����1?��Vm۵�9X��j�<�~�m�����.�vɛ��fE�0)l˼�F����^�(�:=�B��&��h��6�k�N��ڏ�RH�Z8pq)�p���r��`i�ȵ!�,+r:�w�j�&?�R28�X���ӄ�p�2N8B��r�e*Ē�GHMJ��˝*��'���)ϊ�9q"4���C2�v�(A4�(_	x�m��Z��p��
�&K�=��i���̪�3"N~' &5SV�|cR)��rƦO�M�H�5~�����n��P��hUl���>�mr�q�zh��7�e��,��D#ڀ5�v���T��>x���QN�(Q�q�)���C3����r���PE�c�I5%��\��R���D���C��h�6!Cu��~jeM���
!�������z�)��i��DE�����
�ֽ��]�/�����?�������_������Z�鮆�a��mz%�j���^Y4M̻�D�j}w%Ȧ���5�X{��>A_���gAm<��Iϒ7ǧ�/���{x���prvt����=Ox{7���y����8����ko��W?��_��w^����Ͽx����O�/�\��t_�}����W���gWo믐���vM�>�y|�?�_��Õ��������;~=�[��񵯛_9u�8��������ӺS�VӃ���uN�cy�wp���*{�_wWE;��m�����b����;]�`ݮ\_��h��x��g��s������}A�3�'qx|�����o}x�<=z�F�ן_}�h��[L�/���7�x���k�\���?|�W-o~���O=zr��h��i��ݎ�S�)��n�ejҡ�"�q24{q�9�k�;���C�Ji2�FQ#�u�u�v��+��w@c:Lʊz��G���:?���un�L1!�п�@�3�]����G�8�0Ω.J�Q2J15�[E�:��m)���[�-Ao�5��\ʤ*�Cʨ"��2�&}��2�Ҍ�(�NJ���b�F������Ҍ�^�kcB_i)m Su?�T�o�מ����-�B�Rh�]�Lݤ�h����D��,���Wo�m�"����ˀ�oxsXɚ� &��֘lUd��"�J�l�7��&u!�C��t%$E�&M"�,�tN��0_
���`�L�@YR�����h���K�+��u"���UN\c9)��+D9���D�;KƉ��NL?Ô/,���'��U�Xh@S
E��|Q��	_-��g�$�ޮ�i�1��9��&�l��1��5��2[��z�t)s�1Z�������[A��p�.S�p!��yb��J�b���%;��
����+THpN d�8:Dӌ���o��:���O�,�!��S�\4g�t~{E�)�%�i8�LÉ���T����Ĕ��FJ�i#��шU�T��,���
��A��}E��� ہp:p~gzk9�!��	GH�F����a�2e�d�R�R���*1&�}�����.��TJ%J�Af�M˂�Dn��mo�J�*���$6F0��M���Α�gv�i�Hi���k��=���%�1�Jph�1�2�Uw5($��w�cvLcW[-_�)]n���G�d�͈�զ���|Q
J)�V�A"�HD�)�D�)Z:r9�*���)]���Ihhӭ(���bl-��RP�æ��F~S~��"O�i��q{�Ʃ
�p8fu��r �*sģU�7�u���0�����#|��Ӂ�t�B��<����8�J���H"gm���+�T"�4��������gʩ��*g9*��*p8��pa���m:@�Qc�V���F���.��@�%�B!��𦏠Oje�B��p��Y���C��q%��6�s�%jJ�v�UBA�À�S�Asp�1U���f����D���t^|4���(�qD�(�jҘ&�C�?�J�`
������_�I�%cU8�L���[B����8�5\c���5gh@�ԄHIq"O9:!���T�T"0L�;�G�8NէnYF���s(��ܮ�Ǒ��A"Ĵ�|)�!`�|`�Bh-6�r�DN���A.��∲�"��V�� ��1�P?�#�����tj-���@# ��|uw	p`���Si�#X]��<�9�q蔂���o*ġc��ȉ�����7�O*�Ji�HQ��4q~L1���w����A��O���:M��qVZE#2�:�������K"}R�,"*��S��魺�X-~�*ڃ�WN�&R]Js��Ek�̚rj�(J��-
�[�ڐ��1&�g2��A$z;��r�(zt�i�p����D_�&�O;�����vכ������e�^�>���L����˫�c�7��{��.�֟=��{�����pz��n����/�	���,9?:�]q�Wod�@s�~��B�g�m�}s,zX	9vFQo[9����?��?�xE�^��lO�Vh�#;�l��峎rӲ��dQ���=�*2�G'b)-�#�?H�������9mE����S�W��H�������6ńתt��`m�7��
��,�l�0)@T�����#$^���j�p"EY��M��F3�0)�p�6�(!�7�5�rDY�h�C���n.�RhJ��߈�������J�L���i2 |+x�.��6u�w񬐱��M���Z�O3p�bH�љiΉ�6����+�O3�Cc� G�Ɵr����m��v��M�iJ�r��2|S�5&�l��!B��kO��-����y<ҟ��躤�(�y)*�Zu��i���'E�6ЪbD���?�߉1�.P��Gc.k�N'YD� L>��(���,>mڃ���c��ɦY��X�7�E5���ܧ��$c�(��A�����kY�Gy����2Ria�:��U펍0[���Q��z��u���j�wϬ��9	����F�}�S����'&�N��;����=x�x����I���{W~ Ӆ�����ީ����w��'��o�����c_���'�>���Ǜ���#w��3��j�߶t��Ojn��ufx�V���c��E\_�~�폍֯[{:ﰻ/Iv��R��$�:7������7�.��c/֒m������ȟ0]^<=>8�ϭ����}�߹��V��W6�yq�3�|��kf�u�����g�C9�Gr�K?�m��!��J�$���\����'��}ӭ�#:ڿ8����׏}���k{��o������?��|듗~����?~���HL3�x�u�����]sws�b�r�۴N;��z� l���m'L&�vx3~����Sa���9m�Qa��O"{K]@E���p�9eQ�e�s;5��iC�+_:���S�HїkiNljґѶ�]Wnٷ���تg�+�T�lkj]�L����-Q!ˑҊ8]��$
�i��5	�	n���UZJ%諘�ǖǾ]Ҟ5ү�Po]%�Od�Q�^wE�c�4"-�ԝKե�c�v�{��S(������6�>�$�e�"P�4m���cm�T���ј�tvIg|%�e��Yx�J̉$�&��J��B|=���jt;E�P]�¡i���?E$��-���-�^�G�4D-I��	'"K���;4�e�Ő�@!S�D}r��̡��h��I��pR��ݔS3Δ�p�T"5~���Ǭ%|�>�R��dS��Ԥ@F���Y8~�5R�K�Z%���K/�ȯtK�\!)!;������cc�N?M�,���1�9!M���o~���=F��+ ��ȗtV��	�Q 2#5dݚ
��C>�G �N����0��l�bz�K'R3��
5F��blR��\�듲RG�2��#K$�R�duel	�`Z,h����s��9'+���z�VuQ:p��ө���Ѐ��) �8�'�w�������J���\�h`S�z�p�N�?H�S'�v����GV�M9�c
�[�>eA&7c�D�΍M�*-�/W(ߔ�"�1����S��M'�R0�'D����"��%NVE�\]��ȍȉC�ӈ��NE~Sc�3�H��IR����S�5�%���4�d��iHj��VB�(�]�8:u"'<e�^5��!>��pb��T�YѾQ���.K!|V���r`~4�����ޢ%�H!D'�
U�tmtD"���E�6�d��<B���J'D�eA��d�Uc�r�RYi6�.+�i9) ��F!xf�4�@�+!$+��޴��OVW9jzn�$��e�Lz�F]ͨ(��O����vF��}�O�.��5/�#�)��V�nu!Hc�舶:A8���å����7H�8�(�V�G��[��|�Q�I�H�i��hL(��@��a`c��n:�i��L	� P�T��#�	E�!`�F��?c���L'����*��r�U�pV+;�|Yru>:k���_Km�֕D�*��F�
MV���b�,��{ TBh�W%��WK:�3 ��
!T�J`����6�i�VK�:'R��L����f� ���X��cN� $��>���HW���n��ٵ�,�`
�Bګ��5,Z{�� �A�T.e���4�4���M�,`������s�I!��ᖜS��\>~��#8
^%n�h6����_�˧�����C߿��n�L�xD�g�B����4VW4E+7��2���'��`¬���*��#T�h�
ŬP�B�"�G�-��;���^������NA��Σ�~\���w��d�8� ��^Z��K������w�/�ܼ���t7�~������/��9vs�G�����=��^�O�x���������U�XW7/��-��Ꮫ�g'�}����.�p�]��;x����_��HWdB���Zo'ߢ��� 
�:���?�����b���K�'YB6�ٮ6v�@0q�+�T�� L(��V�/)p�V!k����R��*�_�(pd��A��o��T4�f960Yd K�C�fKƑk��vt;�F��`dqZ��H̍���rG�D��&��l�k)OTQ�8�?�z�8L�++�>!p��ZH=��    IDATSVV���eQp� B��N��?���hL���9S�h�#�S?B���B��>��/$�*յpd@�c��2��y\�")��4�nl!!|�l���b�>�]�u��o�1��Z)&�^�{p��F�u�X�*�r��(Y{�#I�����ҭ�:0�Sz��P@ 
�a���G��"����L�%�K�ơ\(���\�E�'&�~8U����=�]M�8]s,�����S�?^�Ŭ§6��M����J֫4��8�����	�k8Մ��/�d��p �Z&r��<�n���(�3-4���/�
Ǘ��c�}7-��a��ى;%����'�/�����xG��_<;��K<x�O���O�����{oY����������hG�ط�D���Vw�[��� ��>8׽;��t�tᴱ2��}�t��ַ4����/�1s���H��[��z`b~�y��b�-�n���s7Y}����r=����b�ӟ|e����U�>hiK.�.��:&�UՉ���=����'ۍF�W���̋��q{�%�^���f(?��%�ק�>9>{ॉ�����������O=<=8�z���F�.|�Y�2����������z���)뤺=��S�(�й��s;���6_���^�s4����̱K�i� �K�o}�[�$%��:�9��O_��Jd�"x�m�t��򢇂N���;�@����{��rg(\�|@��L��[�������c�9���M5�z�!B��y$z����9�(��IPT:�Z
��?MW�n�
�)YS�^Z8�ls��2|�v	�ÄQ�%�iI�R�,Z�h� ��l8}�B�%�c*�3Ev��7�pc�J>L��3S�Ȝ�X5S�BF�\E����Wۮ����b
�l�J�CI"�IMԨ[���R�aQ����%XH�=׆��0�������(W�8���7��F߯b$�~�Q�Q?�꽎��W-J{>��PBTȪ�������I�o4m]Ui��@�Oc�#��Ώ�A�b�DY��|:Ek A4Su�,�RLE�E4Z�p�bi����"Yr[�Ȝh��z�<K5M�O'����t��d�4F���_ic�0Jqho1�u%�;�Fmw}sF!P�������֮&N�E�9z�Ѻ�����媥t!���BU'hQ�|Km�+MӔ	U1VN��)q"91W����kl�B�2Q
+gA� dE��JK���s,�tS~�ɗ�z1���4Sh�T�����L�d�
i���tSYΐM�M���#3N�w|�"�&�)Z7��8�s���MCf-�J k��\�@QS`��c��li!d㌲���(���
&��h�9��XN�v	��Y������(�~�_�ic꒲i�8��C�JԳQ.J�]��aYj�R�[dM�1�R��r���������hڈƩgj��L�8p|ej*Nz�Ф��=A��`YF�>�h���?�9��� dhKh#Ho�Bm�n��WC�Ҍ�g	���O��C�X9L�Ԋ��B�:��G��YQ�
%�xa���w�w��J.A�P:9Ü&� )Z'�Y4�����h�OM:��Df=7:������:�C�d�Tu�BMʪ!f�|N`H)q�R��V�Jv��2���H����pRH��(,��[��Ȏ_Q8'��4:ܞ}�z� ��_��Js�fQUL9AY�ҭt�cDC�b���S�c�I$�R��z���T=�nK!#nʗ�!ޘxk�OX��h���đ��ճ�����j�4�>E-DK+y��fL4ӥr�hZ�BL������m0ec�Yt�N�����JSnNg����C�\m�?K3�'R�,Q~MV�Xb}��#������*4Y|R���9:7
��!��Z��(�I�R#� Z��U	�s�"?+�cJg�j��L���\&3�hfU)
!�?|��?��(G�cZ4�i 씃�a;�9r!-%�8�8�#�����~8��,Q΀)��Ւ�;��ʿk�c���$2�`� �|��,�o�G7����Vt�� Ha�Mm�qN���@�ۮU~�Ą��_h|�c����e�JX��M����z�p)xK�Wr�N��mܵ��x��ErG�7׾���2{�޹����]��������7>�qF�ۛ�D`��T�+���������������v���J�NϾ����~�����Q>��SIggN��wW���yϵ��~}��K���W�I�&x��F�����,���6N����hODm]�m����إo� ��3�O�ܙ֌�����׌N��Ǵ6�SNV�_�q Y��$��&��8@[�GK3�6 ��,�*xS#�hU8�������B3Z�h��5�� �c�z���3-Qʤ��'=�i��M��ʴZ�Z8�B!����:�3����
`�J�d�'�����S��KvF�4�hFB��4�/��t�n�BƜNc���&� �q����pLSN�	��.+A~�������	brR��紨rC�z0����@�����B�d;�k	�{l&+��m�ϐ�E)G6-d*�*����R׫���2�T(M���I�Ƿ�z��U4%V�#�#�IM�e���KĬ!�H����
�g%g�ەƇPN��N	����>Ho���Rz#s�(#I�k�7@�C
���D$�jE�P�u=Ֆ�>�"&S�V}{ƥ��^z�n�t�d����ۺ����sO�K����G�{��E�ź�a�:��u�~������珎��O����ܻr|�V}Y���������7�����/}F���n�/�t�F��]k����˫�"��s���߫����}k7��Z���4u��:W/<<���[�:�Le����W+}�^_�_��=�R�]�H���<q��|�<R­B�"��\n�:�>��,m��w7:}�����7�^������+6��.^��{jW��~}m��3)�߾�o�����
\����پu��?��98������o��?y�k/����G�����韼�����w��Kon_^{��'��ġ�R�Z�$F{b�u�-�k��]_r�M��Σ¹a-��rGQ%����N��|�;Ntg��sX��z�~�@6U��!Bc�v�1�y*�r��C���:3��A���V!4~�pUH�9+�	��x ���%7��:'��{5���)^�rݯ�v�h5�t�Դ�e��|4S�1Z���LY�(g�w��O��8��[~uE�+!���)_��!*����SQ:�4)�b]��y8Ј�jؔN��'�`,%5>�ç1jJ�P��曎2_�=���������*�פmA��J����֞3Ӫ�_!��Jm]n�;����r9�jX"�������'���+l!�U���Y
P	��d��uRQ���)�+��kEpN��B��\:Ӳ8���M�6��R:pB�L��F^]"�RF�N"��L�6(p<N����p)|�)��R�/�(D���Wujc��WW�S�U���=�*ȪH��F���
�_h.k�yS�E�\#�w�M)vÅ���q�8ę\)�@��4�[�F�)��(���03�e��
�Zn��8�B���S|
0͗Ωa����L�t)n��糤�U�TY�4��I��� �7�q��S-=X;ܦ1Ζ�N0N:��c3MH!�|�C)�|Njj�B�MEY� ���8����F��0�)���i��)�
�&�N�DЦϑ��^�Z���&(A�\�)�� (�[K�h��J�	�D�D(��o$�f#�M����dh�ֻ�6p�B�8�5�~��"��"#˲@���h�S�i���%n�W��"��'R�H�i�h��^nS�83Mx���*��-e�����,d������4�ۈ�!�[��r���3����B�M�4��8�Bh�hRΏ��3E�k��Q
����B"��?��� 8��!� |�u"���i��D�F>���7�1NE��H�2��BS��]�M�\:��*=r�t�9ˁ#Tw�Y���5��R"�E˕��Q��DY�?>�L����/��LYR��M98��ojC��l*Z��� �ȏfl�r���/�Yn��+!��Xk�I/�(� ?��=IM:�͊R�s�M)����{F�,f�iZ	>'��f*�2���.H]AF0�"8�rR@؝V.�VdU�	D`]u9�����I�+��rWe�|��=�h��	o,j�\NM���A!f���R��1�n�f��J�3H}Y4x͠���&f��*4��N1M��Ƒ�:��/Yw�#[V�w�߻�� N��m�0$�cl�8���)�u~�"[�b�"4/3bf�KwWwW>�|�.J�[�=k?�Y�Z{�}��ӧ�l(/;�(yLG�rx�XdCHH�(.�UR=p��H$�ʃ��L���%Y��E�A8�\!B���[/`�6��3:�z-r^:��3"ْ��ˁ�N=W�§��<�^�ʢ����e$�	�/�=�l�J'аmq�m���G��R�	��ŁҌÈS�Y`r!�M\S�t��%$����+�� ��,h����M"8Kw����ٵ��r=v}����=�<;�=���*⳧�\��PD,��x���W�z��J�k�?vr�~̿y�/s"���9���|v��x��{z�������{���7~�k]�tu���<��O�J��Wc+&Dk%���5����vaʵk�z����>"��P
�cH�0���b+�rQZ��S@H��l�E�r�T�'*�U	C,#�r|d�q 5@ʿ$*���pm�m��V���5M6��2��U�SCH�,@�N�zd.�@F�t4�򆧆YO�kh�'$!f��'8�lQ�,pp�i�bj\�E�����g�ń�iֳ&���Ș(!Ș%��M�>�>&W�N!z�C��Ǉ{M>D8��8����oX�؁�(C�D�����I�@�����i���¢%�'�I����r�[gUsp"X��������D���ec2�*�v��d�
���Y8�H
�Oaڤ�/�+PxC�@�h�S�!��e�Ķ��ɫN������*�7�pl2&�q�waW)]{gK$i�� �.�z=w�ulov��k�ॶ�͒�I@�@\.��7�4ͳ�����KN�M���R�^�Lq�~R�%���1K��*P����	������ν��;�V��?\��}{�z���~���}�����/��[����ԯn~��^=�t=��o�L��#��W�/~�������WH*�\����|���pj����;��������E�mq�V�5�kl�'�-��V�k�w;䕔�%Z�b���Y����ᾮ�/y���z_\��ո�F8�H��I�{�+��]���:+<*�Ý�]_�k!������k+�b���a}�QP���)?�������,�o�����G	zy����[>��Ͽ|��_��oy���w����[>�����|�v3Z�k2��9����Pa[����Vɶ7���e�9�����!&kh�5�� �Pvg���=�i���n���ۨ?��υh>�!+ɲ�ew}�,Aۉ��>���9ɝ��t�'��|��N��5d}�lv�+D�ch�
S��н+ʆd�tb㨄f�
@ַ,8*$���q9���I'4�\�^#D�ݸ�}�l���d�ͦ��*�m<|j	�Kڡ�KA�� ,�����j��U�y9|nj�F�j#S#�ϥ��+�@dn��^(}u�
ŊB+D^/�U��5��I�ג¥P��f,)A���x�����&��5q�Z�oe
ԛ�{�5���b0�N��կ��2�!N
��<o'թ5H-�[%�4Y�8f�Ԡ�CY_�CfP�q�2�5��#��ihpØ���<6�j��NB!Y8��O:������WIᐤ�l�ӷ��KG?QG!D�8\Z����WO��F��⨊�p:�3�w82/�~�r�o���?���؎i��>u�*ƐK3dSF��0�k=&D��<'���*�4����gh���e7#6����p48) �8I!�+�I�i����PC3����ϕ�^������@6>��}KDN�W^ف��V'[�'�I�r3�0�� �i�z�!G�L� ���АR�ly'0W��|X9�2�Z!�q����\lL�D�[H=A�g���jy1I54}��&D��E(������fP+#;��C>rC}��r��M������,ld4Τ�4���p�����>NI��zRŊ*�^�J�\�
N�2ʂ#WŰ��Ӹؼb�i�r��gĬ�\���*Q��b���j�d���n�0!p�ɋ���M-��Ȇن(<;�!��.�7C���N�fa�Y�jt���,�z^4�pƈl�U��p���Hs���������;������V�c/���d$8����UCI��z�n��!���܌J�[�0KQ����ҕ���^�&�,��6�%ȅ��:'v�i�ไW@ƨ�rU|U�zwQk#A�B}���dKZ�o��2�wd.C!����F�������Ғ��k���9�D4<THS �ݐ�ߐ�����S�+)$��rRXr�`e�� 2:e� ��>�����D��⒑c�N�4��h��l���i��4d^-&��{�?e��=�5%����1j���[�U6CA��0�a�އx�	̕o�
@ �!��bcB؉�Ak��5`I�U�@>�D+�HMR�)
�����[w
�!fe�R���y,ˬ�!��Gn�!W���ٌ\� C&$W`) �D���-,N5pQ3)14
��M��R���V5g
c���V>\���a냱�׫e~�������oÄ��gH'��F�[���mg4;W9��^�⥠�d�*���٬�'gW�G����+��v�;}�74O��Į���g�eų������NG`�pq�2꺝)��M�3W}1���ݪ��ݭȅ�'Q��?�������+;���V��"�O..ϯ<t��i�7���N�_ϑ�<�R�B��ě�!�?�U���+��y�+Uo)���(=�b��oyK�]C��D���*�W6��S�t��P��!�X�ò#�\\c7�kR�5�B���n+����FN�pimS����KG��@KgJb@x�ةB�����! ���ؤ�)[CH-B��+~+ �X!§�Mc�@���J�
s\��*|�L�^?�lZ��r����V�d+���˫�j�lu�I��8C�Уѷ m�d��/��=}
�\�q'��A4:ldYR!�)5���D "�8{�y���MP��{R����i֗�/q
��^F}��\�S`K��a(�����\�V���o
G�hJ�8ԏ�#���H�t���a�� �-*��"�K��aOa�5
�d+�D��B��l^�h*��D����C-#YR.�z��;�'|����v&����^h��-����}M��;�&�!9���*����CK }U��2�f��g��'��H�wN�펝�؎�d�'2o�7[�<./>w��w��zxe�/�5�n���u��w֮�����o���|��{绻�O?���Ono���;��g���I�}���"�ݙ���Tm_/��pr�xz�rչm�U��^ߺ௙<j.��<=��d����g�����Z��y�(��{��[7.}���C��{������nA�=I�nGk����zj���"���wz��w̮;
kC����b��0�7/��z��kٺC�2���5������;K��@�����^e����p�c�^�&wg�Ƣ�������W�{���>}���ˋ����ۇ?�����G������W�����;�y����P%�f}\�@�V��	���T����g�׶���x�')��BS���d1���./��l����}�u��Ci���GH'��L�'	2�,��y'�=$�����'X�z^4=���
�)���DT�c�K���zQ�`��J|c#v���G4Qt����+���BxEq!�_�p6��3��2)}�$��Ƿf������\��x�g
��{
�UH��&��5�bP=��^�,���R���\�z�y-Y=5�o���%������#T�\nj��W�
.#C�V��Y>>v�HRgπ�    IDATk������5�*�O��Z:{Ux�ڽ6MKꮪo
%�i^R�m��Ph
�x`�«BRM�a������+POD�N�v��^�"�R�lQ�ۼ�>O\v6PO�U2����B4Ma��)V:E�O��;�R�!-)0=��)�h� JK����b��+K^}Q��]�ʰ���&��T�#*Y�B6���
�K`
��fȢx�)��.�����B^.��[��\v\J��6S0��*��,q�B2�d	r1I�s�)�r�V�z�
���gcR`#�;mE�e���%�����4dC03*I,�f%�V�!CTKT1���Z���� �E��9:ɦ��N�-��v��q*�,\�f�����ek�A����\M$8��@��	�e1�k��x����4<�y���O�w��J�	�� R!	��O'�VC��1Z���D�P�~�[���l�o��T�!�v�6E
ኟ��C���0gÔ��Bd���\B̑�ώ|腈�RE�G���05X.x^�
�����m��95�'8�@�M!��iB\��G��s�3���e�{��z"Z�Ra�Q���f�8�S�Z��ǛQT|&���8�P.mR���Efh!z�!ۤdao��P_�K�@SCI��T?-���	��̈S�'XvC:q��(��(�+N�R�!/WV�h���kc�!��.q����B�p�~)ℌ�y���h#�I��afW�W����&P=U��D�+���ȋψ���0��pv�W�Q�k����*�#d�-����Ĺ*F`|+1Dc�Èg�P��U��A��e�5,Q8N���h�yH`WU ;NQ%�Zx�ꏯ�����٩����J��g�\�*ah8Ir�!��}���
.o:�N�����UXI@F.��6>DC���g���[7���k��U�U��eg�K�@cHD�k��U�����4SF�׬b^}
!�z�����9��qJM_K�=����(x����&��|�)&o%ES')m�2�Ό���g�m���R�t�@���X�a�Ȓ��FU%���R�B��6� �#۲�]F!��V��i�&�(�2�a��6�\� ����.�ha����yE���m�?��@↉����Ҁm�*'����腘x����JGS�~���G���JBL}:�hK���e
%��M,re�秏�R�&����T=��/m1W�Ο���˧���N?Suq�����]4�3X�~ ��ٺ����uCr|~�n�v:�}��k��[�S�[�ח��^��~��_�=9������ݭ�7nw.�zBåSS�W�O?�L�VO�Un
l}S3/+�6w������*�}sYe�N�f��!���0�!�ͳN�r!��؎q d���(�Ӹ�r�fF�I�X}3�~
Q}r%VL^�ʘ�RpIWR.UI��t��)��J�Z��p��Z�l�20'W��R.X�Q)  ���,ZvF��I|��z�\6��o�Kekq��e83�f��$x�J�	��Tف�Y_O�#��6[4�_/���X�UU����a$�T|=}�c4�đ����\��+UU^���F����[^!�酛�����!��Ŕ�ѿU�,�B�&�[a�W5v����w����Bd?��K�Rg��ov3̥o�t�L��~�0U���ƀH�%�]�hգ
��ݼ�0���N�S��	)�!(P��KT���
�Bc���y=���4���o��G?��L�O!���J�(�I�D�� �ف�ȧ��7�[�~�i��w�d�qQVs(<d�����qM��)�w�+w.݈|���{����_�<9�����p��s�����~������>�մ�<���7��<��b�����s��d�a=�w)�~5s= ��؎4�ݭ��ܾ=��\+���ȴݝ4Z}d�;`�n�qg����5Pi4�R�?&Z��m���,�Z�Mk��(��}e�ʹ����s�G'��j�N>5\߼�]�W��!⸍�	����� ��Q>��gR�Sg��z��hm#o�r�?��Z��y~�������W���:�ݿZ��_��%�"�|��+Wן~t��_}�KטN�,=:y�۽�!פ��A��mW��o[�tp��� ��� �۵l{�a�ث�`���@"p=�O�l�ˈ�|���y�έzn~�� ��⢼��tz��=�nku�!���M�nݡ�&M�HW�CG�K��V�\D�M�t��B��P�/*\1nĺE�c�3V�jz!�DD$4)E�m5��z�Z��V��D\���nRi��[CR����2,q�NDA��[
�d���y���!�;1pwX�:
�p�}M���$�eʃ������r��2C�F�gR4qO�"���������@/�V�ah�ͨ%rSӖph���UR��ck-������71��6Q�u�W�Y��!�eٿ����ZՑR?���zQ�S�!n�ƨ[}8s��ՆOMRU��·~�\����r%���V�\j���e�&63�Ce�ÇD+���
��:G����O�]�>\�4�C�̰yD%bͰ���� �E�\������ڀM3��I9eLٔ���ѯ�G_�M�~��M.��k���=X�h�ZUZ%�'*MC^x{,2��%bT^����j1��\B�	2:L�Bz�|�j8�E/�W�%�A��$/�&J;\�	҉���`3�Ѵrќ��j��p?,��UH�@�	̨ ��K-\S�>M���� ,!�)hq�Nl
z����j�� �U-��K���*CC���A�8�9��ũ*CxQ��\��!�'r"p��pQ;��M���~s�A�LJ�@ⳇ\*ۺq��^/D_y�ԗk����f�bX�$4�dH�7/I�i)���x�+��&�$޹��� \3���� ����(��([`��'�H!d��&�g#3�]�tCȋ\����+�]\���!)��>"M����$6�⧯T�&�f4-}g\��*�v������\t�pE�Wa5�뫇W3,\��A6����B��CG#�V�2�Z!�� c�{<�h�d�� qy�͈�+!��TŰKmH<��h�(@��4+�=:1E�OͰ�)TX��Ŗ�X=D�-*r��#�G��$H$DDK<��d-&��TxKTِ&����Z��E�\�	aL�&J�c�!l�Yg�
+���[�����p�>�lFj�d)���Az�C�āD��e)��PaZ�-Z����ђ�*=2|�2������g#�a'�W�Z�TR���!Ӑ�@`v��u�q�+���%�A�箘s5��d�&�Q���Z�ê�5�6�����zw�VR.jt��&�p�Z����SRvdA��GH�0cz.:vQ����
Ky�g�o�r5)"͝�g"�r��0� 00�d�i�BJ�֔�I����5��zD��&<W6�
ގ8cF>Qe�a344��� NY�}�!��E/�	d˛�>��]�B�8Hᔫ�(�b�!��D�4��V�l-��b(��e�5ʼ�x�џ�����IGU8UR�6'�W�5%I3/�Ow��L�.�j��o��7�m+pq��	xL�Ķ[�g;?����b�����/W#�O\�����=��8Ϸ_�r��ܓ*>��Z��QM������ �`^z��H��w��әG��w�������Mr.�z���ʥ>+�C��n�g�zr��5���6;vK�W��ZX�E4e�4���ￏ)�˿y5G��X}:��t��� [�\��zͲW>����z:�P:�����$�i?�9n�B �7�@%I�|������K��}��£�+�>Pc�U�B��	�ь���a.��:Qz^�U(��ɯ�ӌ_�R+��THv�#�x���[F��Q��`Ȏ�˕N
�(B.�L*�7h��@}q-���[R1�*x��m"h�Ѧ06ܰ��
�����x��+2Dc4���LD��g��Ko�%�@;�y�P-He�h�ƣ���l:h��@(0�8�8��i���Q�=��6��b�R���V�鵦�G.v!$8��ov��!n4婇�{XFd�q�Os��l=&M���T����0���ϐ\loR���*>�mZ/��݋��U������ྦ�ٮ�A@籠�&���3��%����P}%��Z��6lbC{[�t_.���U��T����=��[ozGǗWO�M�3����x�������=�+�>�q�c����'������?��ݒ�͇]���׻��s_��>�e诉v>Ĩw���ܾ%ީ���ѾlV�_��ښ�z���ga�B��s��t�e��%��������}E�lT����hWw��ί��{��/�����#XU�C����Ⱦ�z/��iA������*O��#�/p8�ƽ���{_"����^�������2[Y��j
�d7u�4^�A�Ct��5*8w+�r}���������������ۣ�������s~n�����w��o���/�^��_�����ǯ^|�j=6'�`M�p����M��Co
jFӀ\��8���۹ʘ}�g�pC���E[=�p{�F�i�M7l�nFzZ�y�eӯUۚ;%�ir	�Ԉ�ڽn��%��j�9�svU�(��rߋ����
q���Ճf
�"6�'AQ����5A!R��s^"):�'
G~Kښ����H
ϐEm�5`3b@05F����E�U�%]���>.s!h�\j�|�,�GK_��\,}6Z7���(H�\�˖?���c��(�]�t�@M�T����2�#�������6���KgI�\4�c��;��Z���c
@��c�{�P�p�V���K��I9@�	�����}'�(wM�5i'�%U�����i�� 4 Mx	�R�7DS���fFݙ�l�\�R��k5�z��(l�icp)Ҽ�'X��Udʼ�֤EV!�t�4ނ��/��B��(�z�vH.�,��W����
)��0��6��l�D�e�QC�V�l ;�[�����Wz���i�%��f8��@��F"A���iE�Y0 p�8��'/��T������-��K�GK!��S�3������>~�KD\��,�7ӱ�x����fs�R����/'�X"���F��X����M�z�M��0^F�p6�>���s���hlF6���;=&{�8�J�7D�O�@�0�iF.E��~Ȑ�OaD�fmE	�����9,�&��k��[^����j\�Rh���p��Y,��8��j�(�\3; )4�V$�L
!�r!�7�t*���H��)�Z
�\8l���X�݋����~`L^F.�؆pdC���jh��Z"@4�)�H35���J.;R��V�1U7I����"3��pM@|`�s�!��x|K�l�.HC����oI�r��G`��&�tl^=���{[Cxy#Ёg�X����hZ���e�WO�%�1+�7/�޻�!\�觕ha�
� �����!������pvl��&->ovŰ��A���p�"����7��	�sR��t8ڀj�-,�����\`^tjyٌ����@F�ZxF���0���2�e�x��Mru���5R�j��"�YvҁwB�F'#���҄�ϲ���1�Z8#~���z�bZ.H�O`�5�hf4Yڇ	*�!�)7���zM�H���l��[9�-;�Ry]6�^�,D�^��dgQ >^T���9ӹ�G`3���O3bp��w%�Z|}kU"��D�y�\MAh"��0B%1&3o!��Y�D [#2Y*,\?)pF�}"����͛2MFv����J
�1�C��D����M{&�ȆS&"J��B0��p��m����V6���=�8���2�L"8���B�B�\zQ�H����Kj4���t�2F�!�u�5�C�	o�"@��&�3<�tƥ�����kh�����b�W@��?����?��ˢxv�H��H�zMA��ʘ��h1�B`��bU ��^�����.�� ��]�)���z�ac�'�@.v
�����ѱG&��Y�����*�wۏm{nӊ<�4Oߓ�맯�&&� ף!����.i�'3M���������]���ŭ��v}|��vׯ.��߮���y�֭x��j-�Z��"f"�����Xs��E�o3Z��B^Q.n��fP8Z�Yc�jl|�P����݂wr��,�c4gh|��آֺ�{
N�cA3�߰��g�Z��Y�n�gK$�Y���%\_��f��OG
C`�I1Y
lq�8��R�Iy�׋r5n8�R@çVI��a�V�2��D�ח���3�B�r�7��!#8�=L���dX���Z�e	��s�5�R4䵝"�j�zL�V�^)ޘ�)$3[�DF����dg���ě)N�-;���5�=�����!P�'f��O�)�C
�1�(0��\�!�Wk���+�+Cޤ�e�Z��S��SR=B)���.�P+���_sljhͱ�
 F.�X:L�Qv��[+��Af^\��zC}�f(o��^(���'D=@�ëg��뵋א�p�cz�x��ry%��.]A�������7;��)�/	o�]Я>��N���hϔ0+.kӫ�4��U	QPC�>���d_�k[�?ܻ�q��v^��j��w{s�+i��'�[������j}7�oc��w��G���������ë����8�}�F��N}٬�|���ݢ�[���(h��彵���Io��������������eEy����sɱ�s��gN,�_�=6�8�7�u8|���ns����&E��ًuO�c���x����{�\�?����+��neA��R��nE:�v�����hw�>��8[���቏��G=�3���v����:�YXK��SKcB��j���:����'7���s��N^���sr�;wg�'W�s���W�����Ň���._�z�Ɣ]�r�J:�1�v�չհh�ی?f��pM���4�(��u�}oC���S���^�fC�h�� u��h�ֆ�BRR���v�M��Z�׿�(J%5�sD�݊�5�`�����M��$}���Ϋ�O��!>y;=�S��QU8��(��b(F%�:1��i
api�z�c�b�i�D�h�� ��wt$�qKa�I��05�UK9D::�E�<)�J��JUR /�#��	���l�GΑW
d [Ñ��T��L���G�w��^�z�� �n=�5#�,,e3R����\�y��Y�ݸ��}��e��'?����Gd����fTOw�do:����XYC��*^k�mj�����)eQ^ǔ�(S� �4[3ML����d�B(7̋�Q�zC�20���w2��>wn�2#�����2|(c�̠���`�\,�X���PIR�eG"0/�8@m&HA��0&)8d��&�<�mږ�l�Ͷ�n�9��:v6�XM�[�ҹ/�E��̶8ąU/�\
�2z��a7Y��A�TF;.֎���4#=�t�֓Sa�"ґ�β�
���N3)����&�G(K��'�yq�"n�z=�/	�� ���* HD����8/<r�RI+����Ӥ�\��D��z���֫���mH?B�њ�2�%X���b�IȦ���2ФHv��x��fL^C"�i1�M�8�!\�B4�a���U�-!).E��l�S1l:\
�$W�@=0[x��B��a*�PT�|\�G�Q�BإNʁ4��'�,���K��S��x:!�s�mvZ1�D{H���L��EA
����!��!LMHv��ޞ� ������.oC6Csܣ��*m8�(;ߝ�#U����~rU&����0W%��TUa��e3�~��`v�eǁ� 3��lY
�	A�� �	OJaE���kZ�����![^�d���Dbˢ"$�a�v��c��qS�=)}"
�j�/D,$f�-)>�fd�S_R�^�M���%\ːBKG 3YL
ZQl|S��L���8�+��!CҰ�e����0�C�� ��H�O��Ap2J�WHo��Z�Ü)sm�K${
��xI��Y�f�N��I�����ٹĎr����k����]��Y[�
���F�Wcse ��*5�\�͛+���&i:�e�B�׸&|�E�^�֫=�l� ��    IDATᐎQ�*���Q���j(</�X`
�P�V/6f�
����ɶE+W�1͢!~�t�Gϕ�rV��x�)2Q���p.#�$���>$�z��א��9WW���$�� D`ϢAj���\M�p�𲣙N�C�,Ѭ�@"�z�j@K��_����~eDK.oLF ��L�j�%�a$(P�� �z��ɞإ�Z$!M�}S�B�s�1E��(`��J�oU�D~8�bө fQ�e�H�F�I��\Jd
-H��p}k�K*�a啽�2BF*qC!p�݇gCŐ�$����iv\5j�Z����>Y���%J��_[��ȎI�z\�4XO�ؖ�'����]޹`�.���|=��H�<��\����8�(���R���οȮN|Fx������o�sE���U���ݟ��|z�9]�t���)4\���ߜ���?�����7�WG~�$���P�I5_5��Ѭ��$� MK���Bo:@}����-����,��&f{ Y�M����IQ����X��A90D���A-$N�d;@ǀ�!��蛣�ؒ"�A�>N<�J�H�C&Nx ��r�ڡfN..�M������V0`K�<�@o`�1��N`5���%�W.j� f��#��_�v�V�6v�h����\�0�78
�d �xx��DH|z+0�sQ����I��`�B��γs$�fD�p
�L�H��&�~���PxSx?�L`�e��L>0����GN�`M�㤆��f�㨤q��8j�j:�Dq	�,�m���끤R#˕-�25!@H
��l������YT��!�=M^["Pن���(����2F��"�1�4�p��P��"�{"��"^I�OY�j@�u��7̱=���j#�W~d���#$�?������v�M�O��_�d��ʒ�Q+��_&�LȒ��B�c2Z��g(|"���wC�m$<�������=[yy�����[��̱CP�On/ώ?��;�#w��ٳ��͟��w���['7�?�y�B�l��vݷ�����w%�
�������4ݺ��d������Ե�p\�L�w�7n#6MD���HK���y��h���g}������t��|Q���w(���N*w����ѝ���M��'��K_��v���yI�:Z�뇛��K?�����B�����
l����������b��t�l�T�������1����+q�X�-�?��� �Ą�g+��~�۽U���g��c�n��o��	�'��׻�?�9yry������k����>��׷?��9G�zy�����u��4��˟�ZN:�2����1+io���>?�����1G` �LY��k讌�^,�ܾ�im6{��2I	j�:[�}"�W�D}��s�H�"{Q���S��9Y����ɐK��!4q
Hs'�����s7M`j'휞�M'��n����H..�-�P#�ު2D�&VҧI���.���"���@�B�6�Qp�9
MG.:�Z=4��������+�>SR=���o/0[�j@h�bq����C�a���5���{ϗ��.��R(R2(D�\h�~7`�����Z᳁8��B��ҙˀ�>���'��5�8�&5�̢{��6��Y1�*L1��W���V����A"+�����Pp(�(L���Wͭ0Nk����M� \F��z��-d��NF��m�HQPL��K�>�����2k��::d(�Rp����RH�!�C	�W!�\�V�Pj��d��SY�S_���������ݜ#������mͽO;����i���2��uf��-${�k�y1#�Gy�V�(^C���(\��#�&����lj��l�j�"o������U�&Pa��ddL����Ƌih:i�����fa�b�"ť~=��'�A��1��H!�oQ��E����x�+ �,���đ�+h��(���b��Z|I�p}�����5����Á�� �4�C4�d�"���&JA�k�֚�(\ .�(vL������͝8o��հlL^F=[,�`eG�`m�����A�ZS�r �ڪ�f��Ԋ�۽�b1�U���۷8py'v�ZE2bү�2��pE����&5e��Ϯ LH3���d�z�j��np [_�hh��� Xmh��r3Y��[�c"�B6j��\V��l:�#��n�0(@hB��k@�/�I�=
�CY8�f���ث��Lɶ��j�Tl|5�|=����oO���,֐l"ҥ̈�6|��Q}�t��R��[1 �8E%�&:Z#CZ�ą`Rm� 5�
'2�i٭I:��&�t�R��4���2["��Rc��\LHʣ_l|L�b�o�|^mj(#$��0"���%�/�&�x�FG���3L�Ɏ,#|8i�?���b��
�6�a� ]Qb�0�֜�SlZ�#=�
�E1µ��!2�h��y�!�l6@L��Im�~�����Ҥn���!G�U%��`��!�ҳ����b{��3���<}�0s��>��!������������pIqb���7�Df�5�C�/�:����t��١1�������0v�D؅�!����5�}�3��qf��Ĺ�*I����@=BL�*����o�U�H���!���5d4��;C4���aXr3� �Qx:��`��>��p4ᚡmc�\�l[�D{/(��,5�aI��2M,�/���7}�y��$D�ֳ@:2vL� �j(c���Vm�2�a�a&;�>0�q��8���B��!�����V��D��J��H�M��Y�@�<��KT8~r�v��wG7痞���a����������*���C�i����u����¯f?�:�ݺ�z�st��2���������L��6�O����ͯW�8�{z�eP��	-�tr�{����D���,B�3;����4�2l��\ع\��3ke5� �Pp�,�*`�i1�m��448�-�0��&�X�W��V���8}�)!���R=~�$��\��M6q=�����t�C�hZ�pd-���!M��!�7;2P��x3�ǩ%2kk�&���~k�.렇a����ޑ�B.E"zmb+,���B4^6A
op�Z�GV`R�`�j���^��0'R�e���掦�����q2Ҭ�8�	��sA��E�#$[.��l.}�C$oe+c���U��ˮ0��`X8�J�qn��qʥ>�5o�)l8��m�~��4��jk.�q�^c��g�	�Ƌ�Ձ`c�+�^�8��D���d@4"��ϲH�{�6k�^FpD��F����#��Z��z8J���QӸ����S�S�B�!���IU!�0�5�r}�T),�K�.�"x��P
4�CRl���.�z�󬋛�`P��k��J���a]C$Dݕ֮�z�'�K�`�ݑ��w劖R+��5�B$|8�m7X�U���m?w��|�?�y�r�y���+�,����Q��Q�_�g�/Ϗ\G�^�h�z��{��������ͫ��<7�f���t��Z��$����Q���J`�zl	��F뿂�m��ƵG��4�S�u����o����������YZ�d��3j��]C����=½��������n]��o�3��M�����j��,��3ss�Yf�zft�q}�:��O�+������Y���7�[]Kn��gL�V]Wa|*Y���p�^/�C���������w�j��#_Ck-�3��6���>U<����H�sUa� c�NɇW��~������w>�����/~st�������K7�����n���_�֗�����:�M�՛�m׵UʥA3!�w������e7�G4��u���d�m�^m�?1][wnk�:�f{�\�߻�ɮ*'ĉ���ٹp{�cS6#S�^��g+)�N
���)q NI4W�ewJ�����eFB�Ys���k�4�KGVy��/�[h1Z
��Є{����}"�ͱ�tZۆ\[%���xeh֖2���jD�������0�5���n������t���z�b+@R#P.H!��ޒ�|;��{����&I�xs1��k�1BP!57�*���ݝr!�^f D M���Kq�^�����
N�t�*�)o"�y!��d*Ty�t�$D��|5��[�\�v���ʀ�3���梗+�b��_ofl�pN�(.��V�^Ch��lTIQ:P���a��P�EY�b��� %�&\eQ�ũ
�����e�&֐!��@=���"���Z|M1*������]��ɔUEċ��zo��8|��B75����fӧ��aj)�
*������^���E� ���J�iI�l������������(P�}-��㻕�S.D`
�5��P�R#�24)H���Zj�鋵υ�S��Nӧ�x"�5`��%!��+��q�[7���K�ktx2C�jc�AV$��^C˖(YF��M�)�6���A�A<�p.S�[.�(0�	Z@⥆i���f�Gl�9L��)Ga���Ҥ��8>2��8��r�!�kUA�)�ږa�5Y=��a��S`���Wl�j�[.��m���8�� e��&�0UC��ˌpJ��������2dK$�)Y"�a"L�N�Z��Ů'X13��:}C�~3�hơo�����]��b8�4|��5w8�&۰u� �66�p%�W��BAk��щ#\#[Id�zC�pE�q"0(WF�|=��GЫP�쌦	L��")�
�e�C�>'2Y.|�
�)� @࿗!MA����J!X=�R�Z�B�x[D��!���p�U[OS+K=�J����td��#hZjz^��>P^�lC
�jd���C�)��M�
�yрz�V`��\l$�@!M=pp�r���x�ȁ!�}
MM���*���/��ȉ4q�TF�����6^����(�!�!r�"�1i�V<��W�	�����b�o���Z!!4�1b�@ꛯ�f�k*d�;;�9ҩ�V�d;��Є��&����*U%Z�Y���ʋ��"V���c�ѳ�#���S�N*���oGf� gN_������@4�J dp"��;�)�dR����,D,���	���F#��>zE"T��O.J.F�4�����,5����k��р%��q���o��� '2yq�P@���k8b��eh��\����E-����	�Z�Ʌ�B
C3A:͋�����P����;�Q@��W`4�GO9�@��b"G��f��B�DT�v�2}���8֡�M�}�AR@�
t�����0q���`��*VT�f���R���!dU޿���*�e��zAEPm�>�@n?S�Jw��nN�x��Q���v���bj���o\L]_G�p��
χx��0'��tN���ϯ�o����8��Y�.	���}/��3��=bO�\����$d]T�>�����7�U�83�ّR����[
��֛���4d4�6��`�{�T8��p�֪>}6Cٓ䪰U���ҽ~IdDֳ���K�QR�j���K�4�ȥ-ѭ�Œ� �����b1˲)-)CY�����h��ՠZyD+��5x��!�K�En�@}���;�	��7Ӣ
)ŨEX��F;\ϥ�v�Y /��I����N6�^���G ��Z)�as��U���S��n���/��G'�����I��WC6oG$A�&*evU�hU�pv��6<~�6P�WT!��+�&���v�=<�<[��y�/����VP�TC��;�A,�N�^j���p!l}eg7�7|q\x��_��X �,��l���v�=§~.S�,�������t�-W�������7 �k b�s��,�f�`B����r(ۿ�ŗתvE�l.����^OAyU�Á.t��&J���)¥d�RC��BW[�-DP+[��p�|�kI�7���n��wϾ����{��R:��c���m~<R;��:��n��3w�.��w����������������O~��F������r����j�(�/�#�����ׯP�n�g-anm
X�k�nb���%�t��ĳEl�#�G�'y�niz+e�=mg�;��>8C�l����������[���6�a}>���okZ���#ꮥ:Wپ��_5yq>�X�o����://�.}a����U�	�6Њp?sMӯy���f�:v��޽��em�U����}�#�Ӱo��^�%�f�&�{Jv}��Z����iQ�8
��t&�?9=zzty~v�����_���^\���>��������n~���7QxB�ܗ��^ny�&�-m}��n�DF �j5.���ׁX��
��l��r?��F����ln���]�R �3h���>'a
/Wj�R"�o �.�0�r��"��t��0L^�!�� �M�~6��n0sK��YI��46}|�ދ�I	�,�PQ*1��f�V^^|^���RcK�H:^;��F��ߧ���Ŋ�%Z��@蔧#|�����,���
��y��cڋ>�)����]8��R'%o��px-��1d���h��w�N.��ܑ���%CM���N�##��`k(��$������_���f�P�(���&BJ�Ү�e�{5��O����U%/�nw�����iؔ��4�A��%���S����pD1��f$֝6Q��e���7J-��D Ű �4#j����ՆC\%V�1*�&����d!�z��?���RB�,��b
��/\o�����T3��
賩�I!W-�RT�up�ړ�z;Gj
V["�R{�rt�n�9����<y	*�!M^��=�N
5H��U %5�v5Wu��mT�	aꟹ@H�ZYUK���B���E˕��P��)�m�ĭ D���KGA�m I�í)xe'�Q���4'����B�S`�$��e#0� ������fM�Q=8�1�և��t���rX�_�*d�o"�s��Sf���Pk(6��5�( �D�5;k�Z�{̘-r"����brA��"���@��/W`S�K�`eX1�*�7�MiE�B��q�T q��Q�4�b���x�����5Y�o�O���"^.\���l+����UFʳ�T�\���)dG�r��t�p�z�jS�,W!����Ga)nkB�\
4[7��j�MJ��kl�&BD->M��	2Dy��tj$���lv�/�W��g�1��V��W=�l.�
@�����+�� U	,�(�AM�%b3,,o"2B&�6�A���4F6�p��R�;��)�{i¡�ح<A����u�$o^�Cf�n�E�+c�"����g^�� d3f�R�^��JE����F�)�74}x!q��D#"Sa}�l��W	��fdW�׈�굩_
Q� l���t���+��)�`�r�ҜcZ��"�H�1�|hW���!C
F��5�,5
ZQ|}48�E���kUᕭ�䢐�N ��!�υ`F�h5x꧀�*�2�K��Q.�a5.����r�S:L��e#���Bjl^��К>#����4dpɲQVy��yi�i�p�'��hF�Ԕ��҇J�f�Q5Ȉ�Ɖ@��eh�� }�X�6E��1)W�X Mjh��Sʥ����C�(���X��:��S6W��錗!�K#^�8�&H��zMU��Ze�]�!�[1vU1�Å��VI=�dh���Q�*��FJ1DnF�@d��3,iy�8���c�\��QϦ�n�/�׳5jbyc�e�S���))�2�k�C0[��L��N!�(CM�&����Dd)E��)"E"��e)I��0/��C`�����/\IzC�������-��9z�h4�8�КT	Gߔ�(�����H�LJ�b���!R����`J�9��k>�7Y�f��|k��7���J�7��)}_ض.	�9yi�����':]�]e��:޹8z����c��r�M�zљg=�}՞�BZ_Vk��6��z�����
'q坞�oCg��>�Wڞ�cz�`:�g�z��]E�LG�U��|��Ȫd�?Cv��� ���G�`�pM���0)k@/�r	�#�]:LH!�Қ��i��#�c��%Y��
Ӭ�Z�t�R�aZ�t�i���)CQ\�z�h�뫜�Q�_    IDAT�!�T"_���5�l8f���FY����B2��Ŧ ���qBȶ����Ɏ_���;6cJʨG��f�g���#0�^��!լjU���f�~^��!]��t�U�f�1��B�ؐ�;���'�O��Z�>�I!�M�fe#��@-��i-N)�2��qXO��,�V�5��(��	�Z�*9����[�]
�[א�o��w��^�߼�� ���9g��\�nuR���X=��\���mmպ���)�^��X:lRlY��j+QL`�T	[��b��ˀ$˨R���5�8����MJ�Q��Z�j�ޤ�����my)�o�.�Ș���^"��B%�+�R�������ӵS���w�w�\h=s�@�~��KlB�T�`i*�݊��
4l��C6i�a��(j���Z���Zw�q�.��@pu�:����^5ܖ[�3��TϞ\>9]_�z���������?}�s�w_��v���t��Q#�\���w��׹����!���X�n;�֣��Sc���������r��� �-zv���vGГ���#_��p|��q� �;��7�/�������݋�W�w�
�k_�K��c��_�ܮ���5�I��v��\�����ٳ��=[w8�����/�-ϧ�WOΞ=9������������tOxy~|�~��=�{7$�\XR��@a�Θ��Klv���-�3�m�C���m3�?��Y��������c�ݖIݢ=�E;�x𳧟���������_�`���3��߼R�o���n�Hi2d��T���ٵ�����Wg�?@���#�Ya���خq��ib
��c��DW�;�6W��r�R�@��VCժ�~�T�+���掅��D�N��f�@�lv�������A����Nl�:�;��V^Sp	��DL�m$Z�٦I�"H7�e�\��s!���!raҤS�y	6G^�:1�φ0��H��,l|MRB�I)@�B�e���L��q��v���"�x)M-��e7/��DD+��l8�^y�����4I1��(��¶@��h���b��׿�u7��֦b����L�{�GD�&hF��h\6 �@d�Q��<Kg����G��:�pfF��54G��&Y=�I���",@��~��K��^�7D����&ٜ����"'?��U�������k}�[����p2"�@�c�u�Z⑒i�c
T�A�mU`(���"�.#�!�4�h���g���u�������͐mɠZ�Ǥ4xY��脥�TZ��[o���0n�b�x`����=�q�agZ�}c��4� ͼ��EF�]J:#�#eYX��qGMj1��v�tC>�G��
��'���������#�f
*O�@:I�[����/$�o�����<��j�@�p1�f�]���Ő��������@���_��-%�!XE��UC��0�R�p`J3�� ��.��f�3��);j|�������Q�40��"J�\&�39�4|��q�0<#�9c�h�A���f���,�,˙#�@8�d�^>d0K�A(`����%�>fz�Q�-m��3���ܤ��(�c�����-��	�jN�O0J���4�"uL��5�1�O�UiLY1�O�d�	Bx�hKKJ!8�l��0��6�^�8�0�6�+�QE4�G��k
xg��c�؅����i,�[�LiЄ��!'^ V�Ӱ���~JL��H��	�7X����L�pxu�[��ܠ/4Ge�2����?!��0Y�"�7�;r�JC�
/P�L�	\R���.����ʲΝ�R��Q������k%F�c&�Ӷ�1AjHU�F�ARhs#���fzx��1OS�ic^�3���hif%p)C.��3��̹��;�d�i���'��X'�	���Q�R���0yb`UH��g�H&��d,1�d�̓<|} s!�'�L��Q�,[�*��
��>��2+|T�\�-�4�B"$e�Li	 ����G�Y��!��p�-�!�΁��9eT&��%s��$��E#1�Njx�����$�e`$`�_01�c�A�dI�a���h..����ˣ�<�}��4��A�&�M!ĕ0_QQ�Y�d&s�b�E6H���b�;�=��ni��; 9Zx�����`��F�)�=5�x�VtJ0V<8����`dZ�]tzHI�&���*��h�ʤ��)rȼ���y	��u��������|��Ġd�3�%Slr���%�
d-�tb�d*tQx�'�̲���2�J@b9��o��`��8�s�r�9�el@r_�LҀ�)��	����4h�,�W�b6,�F�  �i2!��X�a� �ѓ����p�,3�dr.R�N�����"1�+0!�@�_4&�\�)�;�4L&Iz���Ne�@..�d�2w�OYΔ�r��VX&��Z�a�#1�=��e�� @W��Le9�WU ����^D3�L���ryˎr|��[�nm���s����S#��,�k�Ob�k92�Z���w|��6����������ocu����Ba��~|�c|5�x!��S�=K#�6b߷����Ϸ����=9�k��$��[�f�S�Рɿz�˔�6��i5 ^����9=!* �fHzr$fs#S�jAH���p�'&Ll% C_�x�J�Ơ	O�РD��e�䘆�3.���Z\$u��r�3!��SQ�5v��Ʌ>���,�/�x(����5e3N9@�6h)���l���۲����8�P��L���l)!K;d�!͵"��k.�e)��"S���@Ec�U�4����,��F�k��H��!�6��%C�Z!L)iB��d�&���h�+!G���ʡ'd�$�1��P�`NYhK#�Em��䒒����w[���&��C)�t��Kk_������$O��Us$���Ny�xɁ{JKz�Y�'SV�]3EK/���:+�-YD3���O]���7�Y�Y-�̻VC��H�BT=}r1��<�� ��3�̕�7���|�'�Ç���%��no����������ġ��ސ��d�d�4E�5y)���s�ZH&��⎝�¾��������s��w�vn|W�B�돽�}�$vo�w�ys�ڼ��?�����;���/Ϟ]��������v�{��6]6�3��j��Y�J؃�8��)�Y�9ѫk͸-
<N�%�q��0���U�ᑜOO�N�T���y�������ϏϞ=���Y��ǹ�8u���@���������xD��X�y���ϐ�H��˗::77�=�}ύ��������v����ݽ՞��^����7H;�=)���S۾�t��|�t�\�|q��7c��g�*帍��������n��{[�ȵT���n��q��En�n�����3OH�W~�K������o7������?����|���
�/��0/_�����rq$�$YnZa�1�4�� ;{	�V��0�,�F�eR�=o�L���o���Y�3B�EDhX7����G^z�#�W�R��).���q	4�ސ �R2�eAE�4��ͥL�ʟɒ�y D�l �V��t�0�J���e��4
�:��8��'��rtX>f�!�K�KL̢=+%�^�r��ILs�/Y���s�FК�����廳)K�(�N�� З*#� �m�.�:�^|�:`�����[z�2[��2�jFNi^��|���� r�[�X���_��Ep���Z[D�1J�"(�QM�^�t������X��NB�
'C$f J.h�`�24P��8>|������&�?WJ*�E|sQ&<��y�����Ȇ�iR�0�rந*�G%w����6���t�N�zk)PG�;�~
�|�����6

#���&�oꞢ>�_�!f�`#G$�j1;��S�!����y�m-$��o�� N�J��a�i���y��
*C��Z���-Y��q�T�c��wqܹ�r8V/��J�` 3Ns} #��F�<�{y�d��LSu��q�եFŶ�  zɘ��'ː_3d�իd0x&3���d�",�`�iY�>p��=���	f#����h0wȊ+
�(C�*#�fBb�%�gBF/=���0e��p�`�@�������@oXv�����A/hq�ۮ�Bc��!?A2�3�i�mT9��Lx5�p��B�eQl��e�`�-+Y �L4� �4���'��� 	X
#%2���(�&�*(}�1�"��'eыK)I佗�d`�F��I��% gK�U�!k<d��g o��
)Uu3�|q*�� ��3dV��a�<i�1`0T&��,[0Bs`A!��V�f�23X���d.�u�l�SdU�!��T��Sn��d�0���.s&[�}���7�*�,=����<; ��&0�)[rV���7X�g�3d�c�y��>M�,��ɗ@c���X7X%��"����\X���Ѡ/nVruq$�󴍆;YKr:v��p���%/��Īf2%!%�g�BiIɄ��9�|��֦�gEh�#�/*Hs���*��1�]
���Qh��%%=eɛ)�3%�T�!��Pt0�L`e&��v2��������ED2�a

I�o<�r�i@�%���WzW��`��)(A�t'��l��Ք-�D� DD�� s��$ai��g�L��(�0bI�z�DF&4FYY��r���UW4.��� 	1�;X�b�++J3^�<W�׊��D�OY��j !���Qy�	��Uܼ�0/HK�����P���E�!<`H���� T�����Dx�I��g�p8GO�F�
9B_VEl9з^��4 ���]+f�r3�`F8�M���^�H�%��`	`�D��+$�	�di�h��0�%��J)KrK݃�J266�*�]��,7��;����� L4L�v�e��� C�:����]nQ�Fcf�g�+�و������i`h:�$��������n�,}���u&#Ct�\Wi��B^` ����@i���
Y��+��/:M-�l���,��cA����ˋےݕ/����6ߖo|۾��{T�/��Ʉ�gz�~|{��Y+�oyovu�\���vt�p�sﵻ>��_}|������׿yos|@�f��Q������j��i���g����|͞�|��۞^=0�Ӧ�W/p���������4 �z�@ÄJhr��p&�⮱��9f ����ftcه�d^e��v�&C�ƕ�>��F� ����1��p�	F�R��e2�0� Jl��`��D曻Y����Bf�X�I)eKYDK0��ӌ��Ȕ@툷���������;9+��Ks�be�^��I���+C�<��BU�|� L� g�����޲v�47�&��Vtf	�+�&*.6�9VKr��� c�if�0�3a�mQBY-�\��)̷��f�� ��%��?��*DyZ�ZΔXeR�d#+Mݰ�e6h&�y�/��N�؄YT�%&�H�C�_n�X�=P`��XH�����ȬL4�"��p�E�3[�3AZ����	�)064H!� 	��rKP2���%+C�!�7(K�KH�z�``�`xBb DE?��۴��@�̓�Ke<�t%�k8R�k��k�]�I�Έ7�=z�����x>��B�ޭ~��7������b���,�Sʆ�Ȗ)��R�T9_�9"�K��_sC��_9B[n�yr���U>����׫�}�����/nV�7[���������k�����哋��-_�f��X�@����s��'NE�J`���]�|³����j�B@)�g��W�z w^Z��w�����r�����d���ӧG'O�O���G��k�����G��7�i>��m�� +N�^=�]�+@�Xdt{�-�^v�����{7=}l���w�ݻ�����ݹ����������Ɲ�-7��������a|^rsuuq��U�s(C��<�v!�f�ۗ�gߜ||��z|���\r~�tuy�+p}O��8��n�o_�=���y�_������wϏ�>:99�����h�ܣ�eؚB��Ӂ /G�h�����3����ySz��m��l��{��Y�����VvV؍Q!�K.qb#��'RJ.F����ᖼ �1�+1/�m{�;bɊ��1񔹏�� ���?�J�
����;nm���M���R\9P�h�gQ�T>�`b�Ţď-Z���їU)�2�Y2@ 7&-A�x�j,�����ױSr�y��W��	}�;�q]bʅ +A	�e[�5h���C�	�dVT��#g%`#�ÀI��!\,��#)J��Q�3.$J���*a�e.�-���@0��~���'�b�guU�(�C���m��V��Puګ�e1#D���� ��fH�?��{���z����*U$�FY�x-'+f7}v��?䨮>�X�j�X��
�=T�^\}��AP`^���K=�;
�t�3���0�ʔ��E���w�u�&w3Z<�4�V$茮.�&=q�4ܣlw���� ���̕�l;�j'��u�����W�;RL�4L� �v�D1rp �u���S���47 �x��m9��ҁ��0�&�0H���:x^��/�(��djix���`��d:���,G� �\`�J����01�	�0�li��-�ǆ��ؖ�s�J�H�d�3+�8|B���OD�aZ����H��dbY�bI��SV�6��	��B���ev�,E$�`p�0��%���-�LFH�ɢ�i)���%��,���&N&`�*���3Zz3M�`ȵ��3���ZA& �ԥ��Jɵ����m$�@H�`���	f�0�FӐ1�Crc�'�2�b�V;A9H�i��܁K�/�$ɔ�������j�Q�Y�w�ӳ��,-� H�,�n�(K��0(���(�f��3^�[r1�ޖKuIg<���E f�4 9VWUT,���s;$=�tGH�� ��4��X���B���ߠ�gIr��4`sJ��4�s4Y���|�WD�#X��#A����O�2	g1,e���ː	�4���v`M�LO�TO�".�����eHf*�8ͨ�����4K�q�Œ���`zN�ds��[]\ ӨN�`�t���Q�d0�%Yn V^VJ!(�қ-Ûo#�i�*�� ��IFU����i�E��^�(���&�R́5*<~�\�eB_��r@YC:��x�"����A�K/=C���R�y	AC���0s�1̥�;6H��d���j�\��E�L(�4� Gˆ.	�� �����iIy���T>�8X��N �eJ[&% m����I.VQh	�Z"'��X�d�t����I����Y\KH	�!9Si��.�#
	��zKzK���FL�����xe��,)a������L`5,s�\{�L�X��@Yi"��Kbd0MS��k8��d0����/=�ہ��A�\\�L��(͠7#,â���o�w9},c�|�m�	F�K$��z�����{�0�AKd�@�|�kB��F�.M¹P C-�|��s�QZ.���F
|.EDE��cE��-1�X`䋙�,�VPʧ��l�s��.��8d%�FE��s<$R�OSh`�KҠ//Vz#�ܝ�j{�����+����4e��%�B?�ʩ� f!�����d	0�ܬ�^�I!�	�����զ���X�	{��+����w��.�uJ:�>�����]��v�g;�����>�u�-D�4v]&|js}5~%�'"��W>[��4�����n�/Ϸ�7/O��{�W�m�koN�/<��Ruh�FJ^�K2�\��2�COYQ�:�j��i�"���&zx�&�*
%!@̖z��)}2$X[b��YK��/��IPlK�it `�k�	�`�B2_xc&�4���MH���)�%3���F-y)�оm�GR�4ɷFZg�o��7X+?؜3�Yg+X�ɧ`h�Pi�V �$���L?Mɬ��&&�a(a����TɁ�-���2��O<=M0������c �8:���f�4��*s�7���V��J���3�[r�}*��)��L_��PDV0�����Гgb�����g�ll^/�bs��nZ    IDAT����h%I&x<̫[H���c`�S����L0Te�1Ȩ�0WE3= �I'f<\0Xz	t�	�La! a8�x��E\��e�r����H��jl�BG�d2�I>%�&��I,B�s�0�`��3��g�=�b0���˙��R��[��=º����&�Po�"�+��ʛ?��� ��EEj@�+���q��lTCl� �qp<���A,�n'��y��5������w���z|���j��w��_��o���ƛ�G㶀{6��:��=P���͝�S�������3���[��й<�����%����H�e�2󭰺�J������
�ы��'ώ^<}~yt�������g^^�-͓����gcg�=t~ �mWwg�������2����m��[~��z<�4�_5�87�V���f���|���ۻ6m�?��;��d��ރ�����۾�`����������{��;�m�K�$��b�7<��Zd]���_E�<�ٸ�<>am�ܒ�h��C6g�؇��3_:�;t5*�5�;�v/v�>��߾������7��������[�'Φ�I��kյMGs��l�-�A/_�Y-˶/U� $#d�y�g��}�{��Q�3�E�0l��J�kP��k�	�����c2=p��&�{�@6X�0c`j$�'Kն_�D�L6�2Q��t+G2 ^W�7�{�B��!%F0��Hz�ș��96��lͬ*�՘	6��,a��A�eR8 �|�"IO���!r^2q��ps� �0Ƹn,� zera5!� 4��K�[�/��O���R��GMH0��QE�L
C��\b�oуu�	0���=L��].l�^�Z���."N�{�����%i��7Yi�� /�$�3d��˗�]�����C��W���܁��˝^���AAy!�^_����`���׍ʧ��W�n�~���� /L�wF�Ff�#�%��V,w+	��/�"�: V�)�h*ͭSw� �0b��%ȸ-�R2Qr78�EQ�L���dCV���P���\V�p���k���	<KH��A����jGk�њ&ŕ�!�����#�&����G��� g��������P�Xvj�m�Z
FVB��k�GS��>`ʗ�Ҥǋl�B��Yn����	w5��1 �M˥�3ф��=_�B$?7!NI��V�Z�Y-1����`#�m�!WӐ X"��ic��l�++B&Cn-�0ظ`��a�^.��]L(��h0����V&H��o!J�@�l�E:3��k_���F��b1�c'y����0��fy���9*���|�G^����Y�5Z�RZ�#q�h|�Q�1C���C��g-�*N#"+f@�M�%��L�Hʍ�0	S�D�?h^��)	�T�\����'�If�� �Đ��DCO&�U�f��k��Ч4K�q4�7�Ֆh���u����2g-yz���̫�I��	-Y���l� "���`�?H���/��-�)<�,��s$h��a%s4s��b�I<y&B�፺�9e��,Jr	|13�)�%Yt�\�u 9k���&�ٰ��lIoH 	/�?@��D.���˱@��S�����R��O�|i��ff�f���adbɚ�U�$c���� �4`'>3+*��k^dS��S���/+��P��@]X`�Ј���ۺx�a���Y	�f^i
ג����a��|�xʟ ��w���4dB�3�_x�%\zeB���2!���!�=�OT1�v���l" � :_>�rr��+3��`|g�dH�9�Y��&G�F ��Tz`BX�|�B���Dcz�a/����^V���㥀��A��	�LȬx�0L��Sxۏ�`-g;���H��FV`�k���>���K�e��#�m��`�%P���5�W�4�c���hd�J ��/+���h`�̼rl��c�NY�炡�0�H���Iǈ�`+��.0G���y^�Y�+A�NUT6��#$;
�B�>k��L3�l�d��2��0�r ^Ry��
̊�AIc��-N��F�R2�lъ�(2��Ґ���f3�{  �3p9�� tݛ��B�)�W���s�X����Ó�w�z��U��1��$�a�����,Zȶ�!4<%�Yuz��nw�sT�p��X��\o�ǃ�7 �Y���J?����[뫵/�uLƧD4||7�_�r������������Ʒ9�l�m��^�wz���t�`�춏lx{vsc��ͭ띍�}?���[Ϡ��O��,C<�)j6��RŎ|�18���u��Vs��|�CI�FRC�'��@�7}��|x,a��-���#�<�d���#7�Ό9��pA^�֖%�����=T���1,K&#ڢwbNe0.���Yh��1H���6y�f`�����d���*Цg"�-Y�gjIoЛokn�s�j�^�)���$K`rƌ�I3@J3�c.1P��g�u{PZ✴��#�)BsM&3/�)�if4񣊟W;����L�%���b2�Ea%��x�E7�P!���3�>~��ɨ�\Z��=�er�K�)3��sT��B~��1
�>@��U�����J�.y����B$�5~|�f|<@�h]8�0ܗ���mL�����!SY���e2��0�!�05F�Ű�@-m	)��d9,!(i��	�Y�@8��@�*|O�)eBO�4�`��k�Ҩ�GM!�`�6LK�7� Y�P#*��Q,���[�����F`�Lo�~��Ge;��{��u�7�AÍ��i�xOs)��+�Y�Ć�Px�z(�)�*�D��C��s���C�}�����v�1�^�K�g÷�zL���ۛ�������o������ų��g��Ƿ \۟��\����5׶�.-ߜ0���ь��=��:��=�I.�U���ù?j�l�[���8�~������=}v���G�<9�aͧǧ�|��a���2]��C��ȕ����,xԾ��]�觿�rS�p+�گt��贾X�R\�o��o�}�q���ڽ\��S{���%g�Ǜ;�GO��p�}px�����v��_��g?��>�9߿�{��H�j����jc�oo��*�@��v�S~���ח7��~��S�3��v.|��?���1�yd�d��Ρ宱�w�����8?�s�p{��7o?�}v�E}��{���l�A_�R�S�ǎ�o�d���pg�#b0���r�r���3�F��G?��GJ;��EfK����-J	�oX�����\ZB��j$�#��B������F 3���ʬe�|U�dt�Gi�,`�ز�*��9��`uJJ�L�H)��L X<hE�.�`�FE�{`����� 4��s���d4���I͉��rU�(�Ʉ~�ۙ�9�;e��d<��J�9��l� �Ʉ.S�by�/I^|���d� ���H��������HF+��h�����@�`=D�X�G��kluUP�Y�H ��Pa�g��@��ڕ�������#1qі<0Z���	0$����htǋ2N��dBY!�(�?3B3_!ܴ��F^>�)%[�L�����yT���U��F�4S�A�͖��Nr��V`���?}p��	��}���&T6zq�����Li�1U������U<�k�	��%���`	|�5N
�]���IG,<6zl�%���K_���cU/��L{I�-%#�:�؟�Ӌ�~0��Ņ����\\�F�����SLs�Lr��]9��pf�/1��+�@>/�6|9��W�����t�1��"��*K�dx ���Mei�#Tx�;=)K�����X���,=z2�VBoO���!k�2�W�|c��4��h*-����ѐ�2i ���@��hY�<\0Ѭv���DO6ʭ��]C�����Ls�W�J�����6�.[ǂ����@�p:G4 ��H���Rz%T�&>��Il0��=�IL�� }��!�E�TH��I�� ��k)�4�2kw�R����J��4�� Ѱ�0��L2Y�׌$�j7s,.�B3j��M"���9�Il��!V<�Z����r��E!w�*8�M�9�Ԝ�0z֊��ِ���i.0>�(������ T020H�F����)&3NJ f&$�>� ��+��i0X�h�J�{��Ɵ#�X� ��#&���ǨF^�z���� ��[�|��	��B��9 /�!���X��L�$P�%#�L/g^ (k��)�*��Ջ���].�=���Ow�.)�4E�	Ƥ3��tRX�B�# �gt�*��$%K���i�L��A��6�!S�fK���2}��fK6�ac%`�� g��eN�>NI��Y\̬d.xd>e�eS�9:����lڲȐLf�j�/%��5i	��fY�j^L2):��,1�4��dQ�|)�3�A)���e���ɮ�����H�f��.0�����+#J���H!��� �7�	A�i���Qf��@ �n��Rz0�3�������(Q\��D���,�ę,DA� �vy��Ā��!H	��������G^��d" �y-�#7K���3=dK�Q�Rʱ�1c�� Cii�NI(�Ґ0���D,��8�9Yc�/D��� Ú 	�'<�@���
d HC8�����U� ���3.r<qr!`�/^|���EV�� }B��U9O<N��X!>|腛� @@��O�O��O��M%1�y�h�G�\b��nPV���ȫ�,i�B�� �	S3��Xj �:Cq嬍��� =	�T��Ճ�Y��(��
�u�$�(����	aQ�%�d���l`FRn3ɣ�FD3_�f��
oiq��rks�U����w��������r��G7�E�g����1}�����{�;WϏ< ��������۸:ؾ��n����m��f�۲�Wg#��N�����í��M?�y�����]ρϽ;��������	d�Ac�Á�`���di��RZڱ�r�W�5Yǘ"��4(i�I�3���F�R�p4��:���� ,�s�4�Rl����:&z�Ҡo�*OV�q�Ao:,Y���S�Z�-���8Z&ch�>c����.C��5�(-mKr^	 -1$�OH�Q(e2�XirL���,�)����XV�z'�ZS.��B25cOH����� �1���6�;�#Li���L�����R\0zV�,��s$Ϡ4d.`ul��6���H��)�L>3�
!0M ���L���F���Zr�_\���%|����>�ys���&�"�on�ln��]�����;����Z�����f<�4�:���,.�r�0��4=%�%�9�̹;�< eAahBb��̑��(M��k!H��r��#�9�y���S{�0|�t�,�K��X�BC��E�\�fʢ7w��Y�$��P��;O <@{���s�n.��O����/[��>��ɨ�P1K�':l2C�創DY=����� ���+i8/���{R�o��}&R=�>H�t���ws�5n��Ƞ�b�.��������������K��w�~r}���ܥ��͏C�^�޵o{��E�[�27|��x��;Ο���[wTEO ��xܫ��xx����j!xց���B－��O�?9����^�~r��ܧ*�}��w̞�^���#�}y��Ru~8����7O> IcyN�p��]wh��E��VLp�uW�$��.<z���{y�c<�p>���9;x~r~zp|��񽧿{��������}ᵃ��6����+�Z���7w��ܝ�M�������j�o��l���x�2�kl��#��#\�
h��ܦ��J��>�m�]�:J'��������;�����^������?>��O~���7[��3������������k��=�3J^M�nn�?���1���Y��r������}o�{3�;U!pq�x$L��pv"Q��Ȑ�l���͌�{�r�̋C�Lzx=��C�&/x��T�����=���_gh9Xr��LO@5s ����l���Y�U3%ӫ�� �X�c��pB��1;L �c-1J�f��>|���YJ�)�;!����m�I; �ޟ1r��jL��%���@6��ې���x��	f�d$L�L�gV�w�{	i`sF���Ph��5J�<<�L4
L���S
)y�C�Aȫ�Z��+�	���ȍ.� K Lb ܅V�X�f�#�2�	��9���$�J�8�7k�|�M�Xj��e0�`S��ɼ��-�����`��"�F<%��\Eo���ל=��F���:f&J����W�2tv8p�%$k��TPl��C#V��C� �R��*�VX����˄Mz�![�����*
�%Y��@o����y������������H������CZ�%�Y 	�b�6���E�3��bX��Y�|9 j�~��G ]�"္{�#�B�!k�
ʒ4�+\˼h!��S��.uL�q�'��a�0�0q�}�O!&��Ysw%���ׇ~��R�E ��2A�@�4U���l���5����1 �UJO��` �k��i�_!�Rj3�Tr:� =}C��J+(ZVBE�6_��������r�"1�+�ނ9�iT���x��[Q��ۖfQ��4A-|!�� �$l=��6��FɊ2C┼<QA��A.����-	�ޤ��Ҥ
/aVT�d�<�@	iI)[C�F�ױ�+�1󄔪!I�5!N�`��!�I���GV���Xf B^�����EB=��������(�,U�0	���r����O/��?hk��e%IA)���B�	���¥����j8�*�XRv��-��x .7�N��?
�(�5:@f�-k�vc�j�FAɳ�K���ǯL�iF��rT��d�*[&z`��$�Y���o.􄢃q7_&�>63MH��H�j�N����9����	�)������ GV��H����<� ���!��MӶ��,��"�0ɬ}� �%B��$��4h��h�Y!�)�%AVK2��0�W{zK�dH�A��J9��I��Ld.�1�0+_B��2L6sCP�s�Y��/F�I���A3�y�cq��; x�LCnfK)�
!�*Zѱ��Bf,�������̀�V�f.:�Df���L���S\ � �y��ѹP209��ǒ `6,�hߢ�o`���YWQ�oe%
�`�C?��ߞ���p�9�-�҃���HІ)`#ڲ�H	I#^�&z�`�# fJx<fzxQ(ͬ��I��0!5����6� ���������X��B^&��F�|��;N�0�Uo%W�ޖ���G���_Q2Y :�D����ʨ|� ��@eNc�G���JI�Xpd������0�E�C#���� �B+`,1�s�N@Ri`�6S�%s	LXu�D��F�G�yQ�	��  ��a�%�0J粧��p�q.i8��"�U��P���H��
G�6�T��5
�կ~�R ���	�=r�d��l�+<%/�4Ģ$H�#:}[+����e��Ō���Y�dzZ�>���Ɍ�_��{yq�-����ϊx[���G6����/��W>|r�'8wo|�a׳�;{~El�����Ʃ�|�v��=�t�
��i��٨s�U��n�����[ߌ����O�d%I�VH�r�c ���O_d-ՍHt^�x��D�s ��v�Qaȷc�4�s)�fK&�����
i)�����)|�f	�"#a�x�Ac�h9���o�����XF	\�`I�#��0;@	L�\nU�i���Ɋ�WVH��d��9�8q������%�𖔼,1�vJ��Dl��c94ӇI�K#�ri��h�Ini�Uz�Hr�/t!̓�*fD0#N=�1S%,���1��O?-��O�/�^��|�jӐ!
ZUDf"�JCni�-XT��`(��`�F��	�>�ʜf����@���"`K���L�&�|u3>?�H����    IDAT����Ss>Vnں�����Ƣ��ܸ��Y�i���j�u��զ���X��������W�.�ח{�x�x%����n6�}��_�s�d�r�R�;��Ct;�GکƷ��${�A�ڌc�Cf�o;<NR򭺎c�(��y�-}�X�'�L�CO�Y�6V,鋘l���`�+M��Dec���s	IY��&����B����&7Vϵ(]�=��aןy���Y\Q��ol{0v����ga :�D�$��IL~L�2#�Ȕ2����e_K������A�7[��k{du�Ú�=ͭ��_�����W�t���f�=>�n�e[/���G���+���U���3�,% s�E��%寍���ʞ^� �����p|	�ŹМ>?>�����gǿ���������'Gg/.��W��­}��`젌C�FAtC�h	5Mxg��R[�eiӀ���+͓�Ѹ 6����Ɩ���q���Ӣ�(_[��ٓOv~�{���_�����������<�>~�sos�z������7�W�z��[�c���]Q�t��l�OwJ�ʟ/�8Fv����X������m���<�8�Yn^�q��f����g_|�����_��W�gn�zf��~�s���>H��4v�w��1F>� ȊHi&�����zK���������،��8��H�$�@�ݎe[�c�N0�F�`�l[�ʡ(�L�����<&gVs�)Ϫ�u�sy��t ���:�����Z�Mtò��j�{xfE0��|����bI�����DܔH(�c���^��i"K��;�Z\�>|�����V�108E�@�d*KJ�� *2��.w�W� t��T1H�@YDz}0s�vzc�`*$�4FTz�QL����m�8�!�oX�C�z�­	�4L V�Gx����@���ki�ɐ��0���.���
Ci@��>pAb'w=���z_4�.9Р"`�!t�:��̓��o��"=���c/H*�{d���e�p�x<��I�UZ�|K���%F\>x����~5�W"v���J���/�4�6ӳ2��	����є�C f�_�"�|�D!uI����j�Q�T�2�R�nٟ�&3�I 9�!���"=w�p�Р��|G�2_��w���W������f\��/��1��虔��Bk�C��eu��3G�:Y7��Nr1$ tWo	��O�BH[�1���o~�`�
����UxH���Ƥ�ު0�����$,yQ"�F��������� �D'�T�J�+(%6T��PbB
��`y/�r2W�pȕi�9dEAd��4�-��b�pK)�r���l��`\j�mhu���p��4�F�K 3�Z�o��¥4ɫW�é�6������GA��
������gAahS�0������~f֫jq6}�+_���^r�>�Dx����� � g�oT��Sw7���nQ�G�_����o����"vR��<���#!`6��R&�׾�5K�j�c�1����҆��!�(�����F��Zm�cH��F��M��`a��dQ�#<���i:�TM��Y	L���r䥫�^��ܥDp�:c�	8L�ڋ�;+%|J	;<.H�� �wJG�����\�=rP�'���
��B@�@���[40�2*igÈ.b���*�\CD���Qu�b�L9 煍�e21$F#.@�$���q��ۿ���2W��Ye��/Yuh-)��rڇ�s���b�&������rj���)� ⎿m#(�X��J���#��'�� ��P�̄P�����������|�����D��J�1�������k6�/g�p�7S�)+ܒ�I��H�2�
J#.�r$���lYJf�Q2�]i�l�Ķ�A�
\�Z�H���'��y� Ȝ{<��`�2-%���d 7��C�5S��F	��|X�K���Ӂ��0��5� ,A�9RKU-��p`F�W�(ؘ�B����vH�L0��	��\��B�"g�,�䁗a���J���Db@ʧ��K1<0��Z�X
�7S��iΝ�@lȜ�Ҽ�}YfG3* U�+Db��x���1"���`���:�<	�B*�FU{0r#�U��K��e"�p�� h.�x �G��%���eII���ir$8X|�ˋ,��$ZQ�	�,͆eH3!���$�@ds�M0Vʘ2hқ��#��� I�q�q*�k��!z�sa2h��I'`m)1 � ,J��lD+[�'p).#�X�4�R���u!�{J	D�������
�?Z1I��,Y!�h�3���s Q�H��3Mz`B��C6�b��\�1�� #4�1�£X��=FR82�<� k�K�W��ַ<�S�>ː����LQ;
f��yj-[z.h�(a ��BS� ���"4/͡�
ܖȋ�p�����B�L���w�{�����L��֗�^\�]��_��B� �D�jo��sxg��i7m�����������{���ܗ���dcu��6�_����z~X���ɴM���G�����҇�.O��ެԢ(�KI	y�K�#RQ\�ZDi�p�@K;��Bu2/��`Eb6,3���5/�5J&�B� �TS9���Ï���`O��0��X%@F+nK�3K��<e�Z:�!s	�di���39}��4(�)K���{��SF����LK��Z�m<%��F�r�<�x(%���<	MI�ڸ����	3�m��S	���S�%%@�rc6
�
�
��Q`h:|�bK �b�+�a9�/@ɷk�aƚ��d�P��L)s�/�����)���ט0r�S`�2J��nr7�V���;�W�Wn+m�n]�$�r�u�ru���������;>g�G�Xr��}ǥ���A���=��N�'�74���>��O6V�mm����L���v⠸^�l�_"�^����;'B,;�T~��A^�������p�d<C�\�+��ЌҬ�m��I	`���K�`` �-��g@9(��f�c#��4X�<֘U@�N�
Fc��ʗ�3Jz�,p&�kO0���wM��ʽҩW�2ﭑ����ð��X�z~��#.F�K�$ �f�3���2*�����Ƥ�j0�lT�@��6~�����y�>;�9[��Ջ���׶�������;�o]?�|�t�b����^V��\���;t�d2R�|y�x�pf����O�|ƘF�2k3�z3�Tn�����s�<?~~t��ώ/���x�������_������J9]ڤ�,z�,߉�4Ŧ�Kc�:�m��Ǒ5Q'��]9Yb/��)4�C��V��?x5�z�W�o�����bӦ��+!�7Ϟ�?���?���/~��_��/��^~fuqg�7���k�ۮm�����K1�������/n�8�U'�e+�7�n5����`g�f�����#�;�?�y��w���o}����^{��������!��X����\_��v�a���*�hS��#������e��7�l�բd������f��s➱!�d切��O��Y�f�9p�!�%�eYMd+6ἆtz&'"$�C�B�@�w��ܶ$�2G��V&H� ���*�裏hz�T.�LF��(t.;�%�T��-	`�	h,G�L"*J�8�hi9��91���v�/V?����q�����2�2�9�;���D�q	��w�1�a�L(sC�\f 2��+4K���6fͯ:e% ��&�p��48�Ŋ���W3B�)$�+�;Ｃ�Z�z�]~��E�WA��"P�.��]����UK	(��iD��΄�Q�Y,HVy���/񐙄c��Œ�	�H�a"W]%[
�XxeJO8^0\X����*���2*^���82� )��(�d�oI/�����x��-
���[ը0���4���p���((0���k�t�$�82��R���GR<�)Y���r��<�����߻ϴ$2&'/�فP����@�W8@M ?~K�Qc	U��R0�Q���_�R�Y�q�!6x���en�mU�������ܘ!�8��������
Q0��ݢ^���n+�{nK�:�n�"G"=2��	��40��Zdei�7�^��� Czxh�bғ|J��:�ȋnFމC����f?�;44�t�ڢ0+N!��d���bY��� )��,1���D��}�.�-�����nxG�I�Z�0I�;ޑ���$	m{��!�6�Ti�y����+%�,���x㍶�#i�}��_G�]�L��>|�f��=x$�E���A7ʁ�c�GVh��G�:&�yiw�U��³�X��K���X�#]7�okq4�M/
ZK�j�c�Im������1l�k*�*BBI�LIp\hK<`CiH  ?=	�U/z��0q
A�PxE�R �8�`�m0<uFO�'Ox$��(r����Q��ud5��3�?h!�VU���
��$�L lf;�V��7�)�n�a�HWE��D�Q�Cfo�bQ ��%8@� 7 YE��_`z�@h�޳ry���{k�MK���x���f�!�c��l�&�rlK�^9�T#I��]J21jۘ3����6�v�rgB.
6$NF(�rh#P�]A/�DN/Pm�<ŌǒUV�v8/9;�Y�H�Ifjx�I�/��-�������l�Lpf	�Ȓ�k���V]���6�n�1����@��R�U+\"�9���Lh�B�EOi'P)����B��H��6�X�v��gL������V�`��F�	h��pB��
K�`46��"/�J O����;r��#��lZ��j��C:JI�g�����VÇg��l;j���o�J�������ȋ� ��L\"���9�����{�C0�u�pJ�0�+� _\TJ&�PTikf��i�2a�R�b�-	�hK�4����K��260ݦ�IÔ�����a	ɔl���T��3�R��ڒ`�!	6!AQ�ek��%G�%6Jcd�wr�2q7��ń�^�-�̍YdQSf50؁���
K)��VK��f,��|;},��G���5��xV�D J�N.���J?s�.+�I�
y:C+�)��k`饗	�v��G�y������s:�s��
&B�Q+�^Q�.�s��y=T����nh��{��Ii<BHChi`�(4%�y��pA!a K[&�4�T��P���0� �PD��l�~��x��y��DN�#7K��W��|���c+�r�B��d�_Vd3�3�e.�)IK0r%�(A�B���
f�����[�d�.2�zGq�t}�70�?���=���­]����ߗ1n�OE�����j�_���ٺs��x����k�/�_����+��Q�y�ޡ�ܿ��7����t�2���������>舫�c�Z<�aB���*�,���.ْg5��8rw�9z����;_j�Q�+�����7��"�l���ղ'i�jc�9X� \�qR�rS�l��,=����W�4�����f8}�1��0���Q�0%+%0���Yc�J`���SH������2�|O~q!�`3[V2J��?%M<��63,��p��c�O�r��~&�K��n�#�Ȗ�TڟJO3�H!�{��
g�1!�J��|J,&��N�1�3%�[��&O$vL�EL�q#�wb��[\r��[N���`�
]�G�WO�x(@������;���>�6>&��3�Y:\��l����?�s?������{+߻��Ћ}OA����뱵��腟 ܻ���޼8�:~��'�ܴ�.� ��۶}Vs��乛'{>׾�"���_\����^����ݭ�FΚ���@�K�>�S���̬2�l?��
'��:`�ю�?�Q1\�k �<@��4��ؘ&r9������,:0Y>�b!����ǒ2�M+��L�˲��2<z��X��\�=Xx�%{� ��O~��ӟ��Ə�c�p�M:H0��D'�Ai�k2�n)����My�_X���;
�����݃������4�����y�ss�Ξm�����w��rg�d����ő/D�IK�F=>&�T�s��w-����g</��jc�8����4�O.���x���oT��Ie���g~���������ON~�ɋ�����}qv�������k?*��Ⱥ�Ɏ���}�̅WII�%- cW2$�0֯����~�}��`�@XX�e��GҐ"%r8���Wu�����s������yN�:���g��a�����V���s<���!\�J1ر�`���)��U��O�������i���Nz_�����_\�jԞ�����ީ������_���ώ�::~��ozK��xy�`g�r����xo{�-�e��d|U�ng��S��y|:����Q1v��cٖ���7N7��o_�q}����ɫ�������t�O�����/\l���g*�<������b�oj� ��,el�Ѵ!����^S=��\�����޵�M�m#�����#�m-$�����?A�k��U��:�j���Ȏ&�@�����n�)�xJiF)nis����`����A��8y��t���'@�T�k\�f�!	�(2�:�!y+�2aX�s"-0L�J�F�	L�F��d3����т����vۮ<��b�� ��I&�%�ڲN 6&C=�pM\�dJ����9Lɔ�>r=�L w�R�`HV^}	�M�M����/MB`�n���!o&���qw��33�f��ѣ�?��@gv�rFbR�9Z��&b���̈�;ο��/����͝�&���%y�Ǌ��ډ%%=� �{�f�D":)��F2v/M%�F��)<���R���+z�d��O�McRӑ�8>{f�-�f���CQ�� �D�g�1JL���4���L>BN���bA��eqQ�5_��@�l��?~��
n��J������*Xh��%ZʖF�[�4�叐I��$)�"�d����U֛T! ɼP�"A�6�����x�.d�n�s�LG\k�xQʪ���X�ULJ��$C�K��d�DY��y�kbRDNo:�@L�2k�hx	��@5 =YC��F��~����J��ъ�Y��J�Ld�H����R��Ȓ�F�D�Cg82�ܴ�����I���<_�h0��'�8��r����,%�h�Angr�!Y�L�]L���Pqll��uݩ�]�4)!���E�����V���G�~�i��O!C��pz���jF��(?�y��J4h4)x%������^�$���'gO��R�'G��X2�կ~��R�j��j(�!�u��B6 ��)id��TmJx�<W�\=Ֆ��d$fĝF/V�ܱѨO$4��\̚���Tt�+��N&���v�<ŵo�17Jr�ce��h�f�<#WR`uK��ʮ竩�f����I�ܥa^�K��aPs�8�zy��Ď������\���Ǧ�WX^��4e"gq	�����}ۉL/yG�����S���g�i������'�z��fьd��κ\�/6T���t"� _�f�&�Y�r���7&;�|$f� ܱU̚R����-%5�3/���sQ$c,�7�(B�$�$XV2�����J�r�I�ʂ�IK)%�Fi�4G�10a���r$S�U��l��Q����k�@J�y�1��Bz6,m����Zr�9�4;����P�&��^/\=A�%�LC�D��+�|X��a�`�5�\�q����	�k��f�?�CTrPO'��X8̅ �p����ѐ ��hl0�W^C�Ųc�5�H�D,�f�o�,$ζY9-/C$��~V#�E�?`ʐBP���&L�7d�J�� z��n�ǣQ��)�|�K�3[.4)��"ϺE����!��F�$�Ӑ	��81��C�JI?M�/�5�	SCz���c��Yng<{�>�4�R�|��l� x�|֘�4J&x��(	e��$JTzz���iʤ!� ]Z��c`����d3w'�x^R,���4�!;�@��s�i��9�c0�/rы˪�Nn2=0�(.��,�)�w0wC�W
Hǔ�-6g6 �L�ih�`�
Q�`:$9j�a*��dV���|��`njܑ �/%=��s��$@9���f���(�0B��    IDAT�d%�%�g�V��0�ipJO��ѣGN�h5V.��@ښ�^n��}7N�u��'�s�Xŝ������	�S/�k�`��s���p�Y�g"�v�mE(��1�6 ��pt�#(/��F�u��������9����y[W[�>����\��9x���]ƃ��OZ�c���m�&��թf:o����H��������t�׫���9~���C���c�-�/��%&aTO���	�e�$si�ٺ�6E�ӛ&̜/�����:~��}ŗ��*Wld�5��TIg�ˤdx:*2��`��S�a�J_���fA�,ج}V��|y�4�4��B�M0��I�,+�|�L��%�Hf�eIN�OS��XMm3"c`�0��Of��1�j{�FHи0MM�z����VѪ$G��jXz��ѐ��j�SCo��r��s$�˦2��-�V�0k2}H+����%��+#}��҈�7,�F�m?��������b��/ޣ��u�3��(+)MMs)"w-60� <����Zk������jzB������n_�yC���wS�[+��˭�;�_}m�����s�)����~X��r������_���+xƋ�����Ѽ8�88�)y��{�t��c �;wv��9w>�y����ܿ\m9�om�sX����������E�n�Y��&��v�	�=,�TV��0�G�'sW�@'1�j�MP�c,b����~Iu�N��M��~n� e�E,<�%	��0��@1�K3^wn^�%���J^��^da�q6/o��7S� �׋q���(
nJ�vS��&��!+�e�/ߕUʒ&�j1pY�6�C��ʹ��)���ZW]˭������w}����o���>x������q�f��L��j��/%/��FY��5>6�S�2q�/Y�X��\Sx��Ū�+T�)� ��l5�;ٞ_�}���O��'O�<>yvz~r�~vtz|�_��������F��C�e�/OX#�[���3�	F`u���W���y�xN���W�������6]v�m�XQ�A��u3"���G�{�W'�;�w��|����o�=}��WG�|�������7_�<�;���o�w���W��A9FJ����/�^zh�B�z|߬��)��~��#{�2v�N�����]��gO����_���7~�í�'G?9<���l�:^{t4�WbȔg;x�^�rJ����	�	Xo��[���0[Jm+���J��8��똮/]"�B�!��ܙDiK�BOn��ա_�zlfH�;d"s/�ސ>�)�4��5�Lz$�U&w�uܝq��]HT0�;�ɢ�\&Д��	|Q1�����\�US��Mt��(���#�S	�=k���A�f�J�#�5/l0�:}�����?��@j|+�!�&�th�ǐ	�- ����hL��V�-Rjh�`�f^�Z0d�3�aH��P)�ka�j��5C�L�i�T3u��M+�l7+�g�[�]�7/e�}[����r���I��z��^<� ��պ#g�Oي[PHo0J��r3x��Op7��A���Qe�`}2!��^��r�@�{&zQ�zqO.%���]P����X��ҁ��85��G!,�{+^�ZG	�T�����!w�[)�@�Jy��! l��	�\�e���	g� z�M[P�y��fG��8
!��.�ܹ!O�ȅ�cs:�-=@z���>��e�P_8��VP��u�*/C̐��*+K9�%p
���J�y&�_%%I���U�RJ���U��-�6s�)���~���X�&ML&=$��4�ӐE$��	r@����+��O0��c�g�G%O�L���^��*���# .1%ZC=�$�1(��'p$� �n.�rf��`{�r�v0�CR놎в2$d*���f&z���K8��.ML�T�S�&&�:/j\:6��p֑,�I�������8���/��>��#���W2������q��D�d��5AC`2~H��#=�C��!���G;�3a��/I2%�qo.	zM VJ����$LܦL�!�ы�3Zy�3���0dn? �h \D!ȶ���������l)��$*9��ʓ����z�ku`�.�,g�nH�+�U1(+B�R��'?����jE�ҫtd�D2��'Z��BȊ>%��(TfD�9]'���?��uG+aE��Yζ�痞w�}��q��I��m	H�zߣ;�qb7w���	"������,��p��`r�D�B.�#W�DJ
�86G}���h��
f���Ti�R����wh\�	�EJ.�,���ŉ#�kGQ�%�1�GbQ��id� 8Q�A�r����oj�K<0������^Ҷ�H�
`�gV�k�����0�H�<���$Y��X*#y$4L�����\t8�\�L �A24ZBJHB���|�i�H�-J)i��	IS��5���w�7;E�-�|�2��.�Ń�/M�lHR��z�&Ά`ťVO�Q:�J[& ����7*&`�EȊ�LSm�4̆ ��4�ݺ�2E?e�4^0�!)��͔^ �\�)�e2�3ش�V�yoǕ|� �c��z^Nz`H=�~8�l�xP��@JBiO��:���\�� L�DDLnv#����ꐯ�6e¤E�����V|:�4_�)�'+G��̄�c��&}U�7+�Lz=�6c��D��VA�Af�����h�'�iq�U`h�g�W/O�O�@\.Ǘҕ=xg]��'B�C��/PkW�^# �;������ar��.�&#G2eG+R2��A�5%W�^�4�;��"��7��?N	��(�h��&.���Pb& ��&���ѐ�eR���P�+Y��E�� �W鼬g�2Z#�G����
45�������Dm�|e.�&SkQJ��<%S���j� �����9�#)h����
Mc�LX�Cp+���mI�H�r�� N�����*�(��m��ϯ��{�|v�p�p<�p-1�Kn{c|5�����t��V]_�^�ݿ��z����7���4����O�z��o���/ͱwp�aÊ)s�IUڔ�QU�4;��i�zV^�dWnTz�V0���j$�MVR`�0��y� �!YϷ�S�g}���ҷ�3SGV�XO�B�3*q'��(�>@S�\,/Md�J��,&�P��!%�4�EI�|�$%B��i��$kA�9�-
/A�i�F{�����C�Aϑ�0��E4�sv%�*� �0����^�?'E�A�a$04L�mŐ���'�\�0s+RjH*��|2ğ�a.H2�4����Xļ��9j4Y��FCo�'�t�79A��6prI���+BV�L���C���dA�D�1|���7.wv7�=I�so�����]�w���:������\��;y�����huy�������bu�C����Lʷ�����Uڪa��78����������y�U_�}p��}�#w��ۗ;��r����}9����zi���׾�l����P%�����<��Uu�8�e��=;S.��4��:ǐW%UCJ�����^�Y2Ǽ���iZ��_,JL��*�����KpBWz���S�̏�+,����>���n���旋Wa�i�ϖ�U�[�o��e ��K3��v�1_Wdl\�қ�,���F~�<T�1��H��?��Ů��X��BӋ��ݽݻ���,��?��o����w/�N���S/��}�_y�3�^[.��^O�D�����Ļ�ar<����z�^9L�W�^�?��:�y�F�8y��O����R��˫�/�ʞ�<b�v�8�/AТ{��Hd9���1r�9�YGb7�kB֩__�*8��)��$�0cC�
P:/���3��x�{���[o\��X����u^��Y_�����˳��j}�O��^}m�ꞧ��c>�^b<?��񭳈̨�A�k�٘��z�+��[���>����jWF��A&�3����A~�w����o�x��ճ���������M0&�����SV:&�:�	A#�iV�򚂃��ѣG��wA�z�%Z�ӥ09�Z�0������ B�D�Pzz8B�&����<�Uڲ�GP&2���sO`"h�&�\����T�?�'�r亞v��{x���,�n`��Fi�G	��Ph��LdQ\Dj����BDg�"6� x�M�<y�7�� ��*Wr'2J$�m������PS�k�����ɇ>~JB������2dYK���"�/�2�sē;���'���Lfh�f� gr�4wCA�GR�3Me���h��N߆�h�"c�<uS'p$��[���`�k�\d<Ӱ�%��&q(�6�x���D�ډU �57�L�I��8�%�b��94�#U�&K6Gi�inh����x�[�����!MĞ��p0 ��rB�sIx�|��T�UVe(1sw�WX�f�@S����r�WzՆ�%
������i�H���O�s{�h%S�Rڎh.��ɒ)`�Ja��Pl�\P�C&��� �Ћh��^��Ұ��n"EW1a�f�a!'KF\C`æCI�B�V��)��LfL`6��\�	�ٔ]���.a� ��+���kT�H#�KfFV��i��@O�`��p��hH�i�C�0|yix��s!`������P�`��X�ҋK�
S��D��������VY�
�FV����Vz� 3C�֚Iby	]�r#���"���i�Z�xP1I���\���s� ���>*�ͅF+���BF.C�� `Ja��G���e`ʹ�r�c8"ݪ�j��LEP�OQDģ��9� ,��)+����Y�8:$�J,_�4 9@ƿ4C�q�KI��L��,��������R`2kQ�͎)*V���ܫ9-$$���������1��s׫Fd&Q��  *8�޾r��So�`��<�[�.ڦ_���xf������"��B�z[�����	�� ��>z��q�G�nnz��ـ�4�ҋA�Ul�=��1�e3�N6���!z�ß������a�S��b(g���V�˟��@�)S�*�Y��b��F�/f=6̓�|r�1��r�e]��@ޠJ����ԜPb�G<":�_&l��3�%hX��DKË;�:��ʄc9�`�I�q��?��|��,�▤!e�DM045Vzq�Rb�ZT�0e�}�?_\���a��K�����}叽$*���� �_��_>|��"��UՐ�!`<�9w�L�R�齆�ճ����_%&I�6z���B3[x� �\$��k$@�,\ixY��!#)�z�"�]���I��%Y�'�^�H5&�	���!N9�	s��4Zl�.���S��ߐ�S�hR��VC�Y�I�N/t�0$�����V&0ZAe?k!	r�w����H�՘̱��"�FB�i(7���a�z^f=�l	�y�R}^�����Y���4 !����(C�ifC&��a�x.EυW)D�`��DUJaș�]O��5�1�&��B8�2	�ut�R�t �;];��?*@���h��-���c�X�qa�RϝK/y�w	h1;�8Z-C��M�	d.mQl�Ӡe��@�PJ�c�4ACx0CB���1b(4f�y3E����&K��  ;ZE�'#�$r ��	�r��>���u�z�������F9�bh.B#�,�k�h����	�D��L$@BU�@.(�0N=��y5֦rj�BJ��P0D���)�F3>g1ض�v} ��tyT��1�,Es�q|������y>u���\�_����7�	��|�Om�_�Z&�Υo;<�w�w�WG�3�5Ƿ�1��5i�r�Q;�&'��b�j� p�0_���>�d	�/�5Lch� �0��!�^�!k�Y�ҳ�)�Rʚ�~Toف�z��ZrqK�U����49b���X���'���)P�'7��c
qF&+æ9��I ��C�ِ&���1dl���3�^2�!L���K��e.��E��@&`�I�R�0�-p�x��{z}<���J.�^k����� #�BR�Z���EB�$`�ȍ�	���0�D�Rd^�x0�c��6��a0�ϱ�h����O�:���O��H�j��H�n�?w��q�筶D����ݺ��;��?���_������ӣ����<�ꅯ�q�t�rFj達s]��r�w���q��M����|��''~��z�#hW�;s��n���/��?������û��⾿�x��=6�}����љG�'���������z{k��Y�˱EC�,f�,��&[���AtJ�'����sG�J��n�!�Yj�_�+%ߐSC��Ǧ���5��hȼ�02�!%����
��Li���@��D�����}��Gy�o��6�8��(�7Bb�I#�i�4eC.���I���֚�L��o����W>�h{;G����Gk~�cC�^w�����#�{?��?����<�:9}��#:����yK?غ�H��nc�{	uMB^�o�����ʗ̊�<ug;E�+ �/�0{�ř�~�����?<yv���WϏ.�N����Û�c�߆���2���DUR��۔E$�YGF7M�o�0NJ͐�3���x�#O�.�О�[�Pr�8��Q˝��������_�p�K�=�X]�a�����������;������ݫW�6}��o�?P��k/���*�o��)L'<�9��3�?/��=�������]�'�ק׾"u�/��}��o������;�q����~�����r�^�T(��N͝��njB�	�(���*xAsQ�K��oe�T7�9R���9b�'��L#K�!@F���e��k!1 � �ǀ�X3"A� �\&�@��ˍ��^�qI-U)�,�Uq��\�yvBI(�gg�x!�l��
RD&�=�U#��炄�_8`l�z�����]�M^��]��n�P��wl��C&ĬG�3�i��C�d` �V�D�0��̑L)�\X�$���6$9�v�戄�X0b�F������z�A� $=B�#Ys��.�� 0zy �'8:������U6;����ư
vZC$M�/��
!%�J/0i�õ����	�a�����]H)O	��r%+�2���|��!�]�##B�Ko{L�K��	�����++Ne�ihF�����`Y!/PBEp�`:^ۍb�e�	|��R5��s�45��W�q���$��*7G����#z��Ͱ��^���I,����*,�X)�\,����HՊ��(_^���l)#��K^�T5���IV��ŝ��p�j͂ t�f(t=����V����yQ��H(2�	F�����=w.��2~B����{kA�.a��	043J$8�.�qR�hHِ���P��ZS�p"�
AC���-:���Uɓ	\ �Xe�$[#��|����R�TG��.	fz��[Jz�;dq� (C,�z�9�-y�/r����J���6�9���0�6�;�HI�E��L�-s�\�Y�R�96}J�l`�����	%\�B#�e��p8Nax���D�L���2��Qd^ �4�S-�H�qg��Ȏt=_��p\Ȕ�L�����,��r0$���gq�@�Z�`���Y��Z����U1$j(%9��)�����u���0N&C2/xMZ�L4��"/Ͱ&��Y�;�{��VWL�8]�1�5h֤4J�;~TŅ1�D�.�G��m�S I��� �2_J}RP�!������fM��O��e��>�U3w	@2!G�,�����Ν\J�������#���RZz<�@�	jBP�=0�|��+=eVM�l"Q1��0S�E�f��5iG"�3�i����2Lи$�j�2��Vt�8����#ˤ4�a���w�\L�����K` �$�jR4�� ��#�@.Z$�m����j���Q��F�w�'���c`�!�U��|�͑@c�E�%@�2)��a�h���}��ڌ
�Fk.��L$%J�̫��a�$rz��'ZC!��	������qg��Zb<㺪7}��9�(����iq

O�i�DG;���2�%4S=��0�@�B.P�&E�{Q�����? ��/a���    IDAT��x40�����ar)Z��4)�������O����D�E�4�ٙ`��05x�B�՗��#�6�0⎙�Ԝ׬ ���Eh ����X�/�d+
�(B���j0�q�Rt�'%r���&O'���Fc��gj�5�`z̊ @�	²�����+f .�e�����;�/+r�BQ�h1S��^E�7w���#Q==���N�*���қI$���Hhi�J*�����B�ɡXŅ	C�o�[-�d��*�8jH�fQ0+ �i�d_J�J_\�2�B���f�� d����<+͒� ��4�zx ��U@�*y����㥡�9M�tÝYw\��;��˭]7���9�vC�SO_�7ll�o�^�j}~��9��}K�e��>�rq�M�=�_)7�g�[k��1���/p�R���4z=_�Us0,mVM���W�2$ �n�R��X��U%�S���R���ox�%�8�e�B��02��F���
r:��YV �Ơg�(X���R�����+�!G-����PF[�C���3l���D���9�Y���ɨ�g���M�W��Bȋ�� ��-�4���@`�R2��l�6�7 �'a&=�Z.��g�"�H�@C��H��c  6�jB�K����JЦ�`���L����P�8�1��(!�8s�+B}eN�L��PD$�(.S�����	�S����<~�o׳L��~J��O�z�=ߦ���~����{�ڣ������OC�zv����j��V] �Ƥ���Άc�_i�Z��tDЁ���/^�x���f�>v��>����g�&������ᓃ��޸{����W.�}�덷|��p���a����3�yv��1����uhw�i���qjM�I��gR���J�Um�%�`dV�&K�˰��aB9�㧧�cӸDB)V���̊��I�7!�E=޹�1}�;W�Xw�J�Ᏻ�{U�6��K��䦶�:�e�_��_��-F�(F��o�4&�l�j�.�e�c�M�Յ��/g���5��lﯯ7����|P�1����t�k��������[�~��?����WϞ_�N<��jz�W�mo�&�-��#F�2��l|=�������^`$~mC� _���y�ڭ/�Y�oT=;z�O_<?����'ϯ>yz��ߜz�飝~t���!�^�=�_�::�<�*K��U"W�Y�0z&��jH����H�Q7�N50��:#{O�1���L��.7��6.|a�:8j6.O<66��;_\��~r�>?[�����ͷ��oܻ��l��t�r��y���.?�)í�4�� ��
>E����������z��^����n��ݺ�yo�}|�����{_���8<���m��q=���R�5��V�4��4C�j�W��S�!D����}�:#�BQ�0�)!���5�՜&$����᫱�S���l�<��1� �G�j"�]gr�_�^^�DP�^J���4ѳ
��4��i���(vˉ�[ �(%iRhK��9�Kp� ��e�� [�ʚ,��[�\ ��W��9����XM��$y��/i@��<f^x�<x����a�I�����������!A50r�䙉��8i ���<�*ݞ2��{�J�8�^c�g��PV�)	�A0#��F\%2���_I*���ޒ	�#k{L�>|�JɊнH��5�=0��s�����N���Y�I��rxI�L�!�%�mv����n�4��8ዢ'��;I6$�v��4f�K�%�ʨw{��rB�����u���z�ɱ	��y�Ig���U�0�L��}���(\`R�2A��O�@�J4���悟^\.L ɳ����i�h\��y̐rc���t,Ø)G��LhK�҄g��J�)UIC��L(�"j2t�R�� (AP&.�!-ʸr�w� /�B0�
X�4E�$��+6���B#CR�X�h��PV�&B [-e���!���Df-s^��L��`T�W��2N^�saʱ<1h8��D�*d�|����Q��	D�K�M�l��@Ⱡ�0��5A��-V�Z�i(5�4`�������  s��W�d&Ò�F9㚸������������z� k�	��CC��ڮ-�F/ʜ�LL��b�i��!4L���a���U������4_��͢�N0T�2!hEF�J@��CbsX9sz7;g0ؖ����Ci�!Z��;�|�d����a��C&�f-[=%B��|�3qO.JCx���h��:��R;�^,�Lތ���I`~�_�g��fF[0���̃1Im.	%O�%GC�	zJ�ӧ,"<G}��Iu�4�4p7�g=i ��T���R\z=LQxPJ�L��7G	�sV2FfA���>g�	�Z��9��!	��K� j�	L��"A/O=<d�^��S" AK T�_�5��f���17w$ r��u��'��)�W=�Yk
�!�����Ā�2�+T��3͠��ۙLm`0TEO���( �Z��R��gO7[}.��-H�����D�l�݊�ٽ.�z�lv��Ǐ��p��=�^������cR2�A_zVr�%���h�q�����M�Kc@�
G�\V?�/�Y[�H�b��fP,{@/: r^Z�X`�� �_C_�d�����1��b�
�
ֱ6��㏊���5Z B r9�6YM�e^�"j�ʜU��Pz�8'�!<|Ac�'=VE֖ �kfHV&����/��IC૯�4�f�'O~$��H@C0s$hx4���2Q��Rt��0�U�'9X�L(=�m6^4\�4���Q�&�e��PO�x���������%!:g��W.9\i�W�U���e^�-
+r��i���Y,r�zM��3wYE�0 L�H� }%☬�J�"�e�q�
@@e���R�A"���/�F)"�Ǳ�h���h�oeJ�]A��L���`#���]>�Y��d0J�&"�&F�5)�X	��y2+�4�%`��ȫ(�a��3�S7���D�<��>9r�u|
e�Gvv�w�ά��sy�n�=�������핑9�n���OC�_���s�n�\��c��kv�7��2��X���'mJ���1����@����.`���H���8�0��M�*$��61x��$9_��җ^ʨ$SD$�5�kp�(0Y	�1Ӥ�Ez�Qb3��!p�T2�@��>rz��G^�&�h�	bUr��d��3���(g�Y�nZG��R����W���I��=�����"��O��Ӈ)O`r����I���zYF�o䷇%�����wV��*��L�aB�3V�@�h��0��QM�i�n��c5�A�>2!kA�bã��V�� ?�%�ƌ�f���5�ՇSz��}����{�ln��������gO��>{~�����3(����y�?~3WG�H���&o�k�=��YyR����׮ˉp|�k$0~�S��p[�bj�Fݮ|,lsuv��Z|����^���|�ݯ����o��f��������KC<<�y�ˍC�G�ߔ�L5�������7YV��P/�z�سz���Υ���k��1��m2�R�/�9�!yQ�x�<	��G�X���'�i�U��+Wd"H�ף`)�j�v��RYD���.+w. ���/Y���.%7�Xl@z���T o`h���ۜ*|��j�×T�\�/�F��~�m�>������>Ri��,7e.w���ÿ��߸�{qt�;�M�{2+��_��ӊc:�mzж���rJ�}�^=��
��9��in�Wa�;���9.!|a�ک��;��ώ^�����''�|q�ٗ�o�|@���i��=�����J�ߛ�їM�Bf"�u[�Yk���Q=%+e�L��	0��fb�x�j��"ZP�������#Ӟh:��ԕ��M��ܧYϮ=�\�_#}곧��_�x����}�N�'���{~ |������X/���74���js5��v|P�_a)�H�pwg|�-�x��ON��X��xo�j���������^�x��\>�#��K�����q�.���R�a;�@e���DP�rM�D�re�J\l9�ĸ���o���%{1��c����W,zAk�E�fH�=�$�K�^��!�R�B<�@�Qϑ�oG�����p�,f�h�	1Q
�񊖗�|�"j�� �c���,SiL9JUt�n[�L����`�5���R�����p��wYnv�3�=<J�;<��������GƐUK��K �l.��`������h�
:��#y��@�� 5S��g⒠J �5���/�����!��?Yb�ϥ	�R���4���^����Lii�s�5������B�42����;f�9*#/ ^��=6JQ�*ysі�16j3���fV��z= �[�H��愬�����^��C�jk�Jf�M�� �w��]C�;��ҨD��j�ėҤ���E .�4�v�y���*JYa�O�R|��	z��T��&��fL��R�&�(����y��;PZ�L�pj(����m�4)V�i�rANhZGʙRCR��V1H�4!)�3=/M-g2ӴJ��dX�9 ��p�ʡ!T��\�0E��l	�אC�����H����	�a.=��j�;k��������'d��
 !f<M�	w�6��7 &T�h�0����J@���fl�&�!�̐#MA����DE�-A��F�x d��P�1�JElv�� j`1`���Ap΁F8�4A��!��zQ"� �kȚR>VG>L�"�0N=k���T=2=��EI@�$J����D���f�g��ʁ/̆�"6�4|���}��^%��?���*PT�af�Q�I�B��zCTzVr�h90SJ@^3Z���!�!_V2N^��0QBjem�z!`�c���o&�ޙx�^+x0|������ߒ=��d� +UiX#�JQ1ɐ�0�F�y��X1����\b�9�ro�L��	��Hn:$�O�s�)1����Xͅ\&� w��gS���	�`Ȅr#keB�_O3�>��ʐL?�%
|T��S�Wnr&�Gg`z0.��>	�99��I�J�X���P�)�����/l�2����9N�� � V�������u�4���d4U��ʷ�w �hMS���0�ᨙ09����-M��Ž��~"ek��L���`�d�jQ�q����5��� �9�Tձ�����*yyS�
rр���{Yt\������'�8��"���O����|TL��`Շ�L�"3i �v��K./���ah�㤁F�����\b�Xl���D��ɼ���EC.a�ZVz.L����\2�2��Y�z5d���O�U[+��ڂ��GR�`��Q�9�|��7c.�wV�vNAg�)�9�Kò
�g-ni��򊐯��(a�0y��4Ԙ��50mx	��8�9�p�Ƚ��3MA��x�K&H��x` �P>���Mѳ�c��k��yՀ���D�9NV)�RL��r��8bj�0h�i�ehX��OH�%��,xoI\��|l�&82^���l��Lћ  9M�eK3](c��0�>�10��G�0��h
;���ԛ&���_��_�(�o�(ׯ~��>~����c���s�N$�m eǎ��Lz���ܼDI�7�ņ�Z����^/�d&4�zB����f("��1��)C6�0N!��C���#���\��跗��4+wq}"B
>@2��CH��Ү��qW�ĵ�ƒ�_&�Ӱ�Lv��Yt^� Pi	SO�A,����wsf�f��[qVl-7_�B3�0���Z ��<s+g�9#&-�v�aT�'sAŋUDC.4���d.�zVH��i���"��҃!1}` <�4���i�˄U��	%��Xd�cHB�Y��+f���n(���C�6�����F����U
��>�Y���D_ny�Uc��@���	�s���7��
�]�1��]�����ri�s)
%��UO�<}˓2���W��K/+Oo��@C�!Y�!i��C�U�X.�%@!_B ���2' ���K��;ݘ�1B�Ɨwn]y�yoߣ�+���ѩ�k5w��֞��=�W3����w����L���«�i�v}�cu>v�x��t�>��:��r���om��/,����>O]�y`�{�3�E�'0��(�<S]��p&�����������o�v��+���;>䵳}��>��<we)�+�_vV;���W��kٵ? �U�W�z��a����J�>t�ɳrI���c-}�4��z^�F��X�y����Pk������C�d�~�Nnd���C�"�w=.)%�V�Db#�����-��m��^(�F�L/%g`��&��af��<����5 �4 d)q��+W�^H������s���=s�u�s�ޖ�.^�-G��e�Fuo�����o�e�<�e����̓�C�g���=�s���ד4�ӓ����j<�3%?��s0�W�%mд)y{:7����'g�g�O�<�������/Ξ<���˯���M_|l7C���WϾ�Pn�nRj�L��aFij���d8e<ɕ:Y�J.��'kCY�κ<�������8��u���(X~���j9�O�����5ɞ{����uo�����h��:~����:���Xky��`�iQǒ�98}㾯���p>A�	�GԾ0�_e�.��y����w��y�֟}��/ׯ����S�0N �/���宿rX9��"bi���L	�}eʚm�o�`�2$�5]������'�i�A�䂳(���7��掍Qݥ�!�P�
C���Y�-�Y&�`z^�x� CvL�O(�xܵ	�P����<x �L��:�0L>m�!q`zw�roM���Aq���� >�6����&'�9S���Y ��^/�Y�ʈ���P�w�)�������0�-�F_>'f���4Cbf�b�$�������o[E2n.c30�oR"1����Pb�B�K�~�Q�L){{O���pS+�ڏ�����RU�-�:;�b�s�4��l��d�4%F���n�{���ok�!E�C7�<l��W��w�eTU����8
�G}��O)f�ܭ�KM����4ˁ��� �IB3�������Ui��ҖG`5'3ac"(O�	��#(�&[ Js���43���������mij�C��d����E�l�O����M*���ʙ\}�0�>�@�N�qb��ηmX�/�ak!�+$�Z�Ec��
��Ļ�
����8W ��'�"B��9RB����'�5��j���G�Ut�9�5Gϰi�`�aᐓ!ee���w�yGJ��\{��)���̋�IŔ��-j.�j�@��r��=GQ$ ەRD<�ʋ���iL_�	�4�%S>E'+&BY�fRr`B�2	`Hd��/($G=�=N��ԍ�腠����L���y��Ԥԁ�Vbș�Tх(��"^�0��Ǭ�������gTjeh:��Z��&mCMqŰi�� 7)�4��U.Hֲ��F& gB+"���j�p.�1��'��V/=X�k3"�
� ����� �B�B-U���3���|�M\o�xx�Q$��&N��'��!ǎ��Α{��^_�`4�v;96xI�)N'
�6��'�}���TD�z��$�ՃI�PDCӧ)��|�Z���K@hC<e���>߹j�Cʶ(L��L��bj��ͷ�V�r"/$ ��k�EO�3j�y�%τ�@��!Y&� ��ː{G[�'�)|�N��f�璵�)��U>0���i x4�_&��c����6g�	�C[�9$Nx�5 �d!4[�5�4y�7߬�5w$��� o��`�\�Ba�L�ixu@U|`C�GK�� �H�93�'#�G�'T1�e�IA����d$��c�d[N+APzH$Eq5���T	�`r�9��$�r�r�JSb���A��j |��$���L�!y2�X����U)D��
�-@G���`��=�H�6� ���'�\�ʇ�u�h�/ރ��!��l�3�FI.�K��i ��eΤ�d"}Ībi�'�d���Kp�9��!�vX�*��`X��j%̥!=�7$sԐ���k�    IDAT!�9��� �F�%�\��_��y���U��µ��s��#���*y�R�hFȥ���͔�L�K��H�!���I�G�0��d2"��;J��fH��F��o�����%��kN����^d	�A�eBv���/��v\�՜�L�i�bih9�LI��a�ԚN�b�����E狐c��	s�  ���{5w��}�[߂��o~�.Lz�R�(QU��z�B�����h �D�Qrlv��B_�"�r7����!��E�ov��"��'}�L�r�����Q1�JC�o^4L���Z0^dT�ZCSXPƱ4�JYJ�Y'!e���DT�yɄLɑ���1T=	��5V&7����ɗ�V�Cʓ�K<� �E�`����j���yq� 1ˁ@�G�\���BЇ1� 9�Г��T��R4R�/=`A)��&pa%�!��Ӑ�T	i�K�ϫ�ʤ�Xg��/ۘ���'$Ǭ��y�nv���=ͷ�����kѰ �h�Rb�^��a�� �LY+�h�F�e�h��pV��Y�X�����l��� !��bq	P�v/��e>_^���Y��\���c��)��OOIӊ ǣϔ�\2�$c�p�ȝ2}���/m!��Ǳ�������u~�w4Ѓ
_<��M�9���ݧ8��ӧ. <����~��Gl	�`��Ĕ�N�B�2#�����Hb���K���8̅��ʣ�&���	����ϟ~���������W���������o����;w��پwz|�r�Xo>}q�>�8]�>;���x���}tt��X{r+�Ǜ�nµ�y�팲�ݘ�R4�4�c�����y�F�h���jK�1+}Ȩ 	���0�Ib�U�`|ō���,��	�Ɛ/ }��ƹ�Ҷ�Ѱ�X��B���ӻWv�|d�q)�.^_��ޟx����Ch/Ɇ���'��N�i!�,/rա!�0���!o�?��׻^��}�o��gJ�vv-�W_y�_��u������'�̏����	��wUl�]���	�J]��gߒ�W}dq<���E��%���1��r��1c��NGb�����g8����9_���_�s����{	��0���\5D���%O���L1T2��'�b6;�1��DR�o��(q�y���=����w��2�t<��^]\^����_��~���/N/�����o���ɫ�M(_�3~=|db�d�����XvB���������i*�M<>�yqx���v��}�����������b���~�o�tL|iu?5>&s3��l����cŗ�7+ %z7�]!k���.a���tF�W� 1�ƽ��#Y�e?�Rz���_���B���qw�lrzMDl`�� 4�F���L&3���H�ax�a�$<M�\�џ�9��|�����f�W3��n����x�:#t� f�n�"qr1M��٩_Ci蕢$�	̀.M�x
G�8b��ӎ/��yMg��E#���,"� Vr�x	1[�d�z�3Qjx
��Ƭ����5����9Ze�	*
w^�2��$e�%�o^��3�X��҆�c�o^JA�VS�}^ǣ$�=�D�j������[Ő�����!M��
-_�$�Ø��ǏEi�җ�4��D(#W�iȋ.��1i0�@���7�n[�l Z��O>��V0�p눶C��9�����A�D/C�i��@%�T{�k����E�;QTFz��Ԕ1�e��ХJ��ڢ
����L�H`4J̄��q�<�
.��a��L������h�0��NM,���0�C.�����t5 6��j��)ː	��XbG��#�2�������Nxj|�p��m�К��c%�G�41,7�t9W7��x�_�ܥ]2|��X��$H�"�[ڼ���Kw+`��BJ� fg�`~��!��p���o�L H�@��9yJ�P�
wr�F�A,.��E��d JG��B��WjHV��`hW:���[���_���U�&��$P.�HI��@Bk|h��y�� OF�V�%��U|<��;�	�|lꆄ�<�-�f��?��Ͼr�n���: 'P��`���_�\�Yi4�̑�5Y�=N09� �j��!*0=kx����r�-.����V23(�yp	�Aj��e������&�ы���X%�	���	<Z���b�hY% �Ld�|�Y�oWX_eI?ؗ����V$&I2��PE�!9�慇@ߔ%&�r��2OY���7#T�C�L�ek���A	�J��"���5s�@�aS=�҃g�я~D�ک���2I�B��C�_	���/�d4�%��ʊ&!Z��H���[�40�Z��RbLJIs	I���!�+=l�͚b��Ȩ��g�1�5ԐϩAr��K�!X5Clz&J�*V8<�JV)̅�lS����Ԭx���a3�B�Cb�h
ĝ�!0�I,&�L�j"fZơ�Do�JV���s���s�FH�r�"w��+C.4��c"S6�i% aE�We�E�*���i⹀��N#��-�"���UpG2��B�iv3��VY�ir)���V�2#Ty2w0�������o��H�T����[ϫ���4@��̚��N���UQ�0�k�PU	Ru��U���J(��d(��EPi��$3ոp	�]��\���s�d���u��&=�p��iJ#�!fl�Z;<S�dÚsK�`�Ȫe"�1�k�͂����:�)�0ĥ'�5i4���	5`^��U�к`c�D��ƙ�F\Cu����+��а2��dz��)� ��%�LU5��F�ɋ<�e�r������'j�w��#D�9� ��j�����+�rȅ�� ���P*>�%Y\/��5�9O_�t/%^q���h��zLB��*�&|Q8�kH kA	�|��m6���.�r���D)O�=z�B�kW���GQT��;9B�&-@s�B�	Y�����+e���"�Qh���&�Z1E��a���F�J#����B��Sj`���N�\�2�����$L=�|��.��'z�����͐�[.B�@KohɊ�==�aIN!Z$���3�1VC���avd}`�K+.k_.�j9��Vzr�d�f-6. dzC�r&�A1�Tz.�@ rm����y��'��Pk�4���w�`�J`�S�*�9&��G��*��>S�H�95l�۱Sh0�~�9i�(& �*̥�$�09M<%	I����@��d�[��Ǖ����GR�(Y�m�hʲ��cL�<A�2A���;���wF�0	����C[�(����S~�����I�.�Z��g=���w��/ww��L��$�9(K�3/Xx�bK ��xؓ�&=zC�����(}S��zU��ds
���m3}<����Q,X�3 �����`0���"�H<��tt)�2n�Nn�\ޫ���۫���76�n�x���G�=z��3�U<������t~���|S�S�����t^��E�;���?��ԥ��25���H�[�[{!wQZ��x����C�jn�&7��/O�^��������_�����w��~�;��|�;�G���z������7�WG�[/_����H�<*A�O�k��M�r�8��;>� ��Rr��j���R=�o��l�� T���D�v$�s�V/m��)���M�Ġ��jY�(���>C��Sl��V�����^�]� $��^&|�3X T�|��'�|�sF�y�S>)[#[�bx4�xK��q2$��X��I��/�I4~=���2�/�7wƏ�ۛ�p���޿y�7_��~s�?��|���`����i��q�����/��4t�.�G}��W���6���/}����{_>>x~x����C̓��v'��P�r<�\;Wa�ҵ��dS),�
�4+�ͩ1 ���Hfx�����4�������=�]�/�z��T�/�ύ�NW��������H}v�7�9��_��-�g������e̛+�tp/��6�}ٻ_���1����m��x���~ۯ����Z���jǿ%;�X��|s�{�}xg�7N��zc��ou�{��\�z��4�b#�r�����W^H���ݻw�g��.�띫�N�f�ll����G3�Q����!?汜׷J`R%�\0<л�̊2-$OC��`��a�aJ��BՔ��f�a�$�[`� >_��V�󡼏	�3t����C�v7a��'I͔� 6E.;�"p�]:�EI���"�G�ǓH~C:k�2�C�����/�K��a�����p<�D��4�?9�<�򐊇�	�x�@v �
l�9�)���%$);�مi�Y8�h����K��Wؔ�� �Nl�Ry$�r�T��}���������D���b�Kj��E��$!�\�ɋS�Qf����H홇��
��<�Pj�E�bkنV��9V��s�p�	�O����1�	����E��J}΢�c�Hz���
k�$��A��eVﶠ�0��Y��ʒ�iK��Jǀ"�WFw�n�Qy,!����"�(�e�'�ԝUj[�([PA�w����ǎtE��:���������kl�Ǯ<i���!"?=!-A�XM��,D�d/��������F�u!T(����Q�c(K=�U녨��8l�%��/�����,KO� �.�d@"$��^��\��A��*�Β�+�@��l����[mbՇ3����R(���!e$ɔF3��A^���ǫ��9f�k5d��u2=�D�d���GF:-�A��(���4���.��­�0xQ�M��PSJ�#!جܥ͂Yr�2	n�l��B�4M�E)��_j5��䤹�@:̢��B�� �H����K��.�ҙA���a���`!+>�"c�����>c�8m @@���kDR���kmI>Λ��D�Ye�3`�8��9$�F��#� ʩ"�?��EP�c�oE�H�V��^`E&�* �u������_ou� �(K������#�`}�Hh�"�h9���)����fM�hܐ E�����$�0he�\���pQ��T�X#OO�z)��a��C��F$�0' 6zZZ~ N6'�!�`X�5RH��<Q�GO'?�^H`����^��Z,Y�
)<�x1 o]�2d��M3�!0N60�je�f!8��1�LZY˟NQ��㤖�� �<�Q��!0�!��$R,< y�4���M'g�v'�h5! �\g.i�e��.��@.<�����Ȱ�x􆢨b�a�2�� cJl��-���i�:'��٬쐨�0ʘ�2kS�^1�Q��6�a�Jg6�<-cj�ٻ�3�,!��0xhfw�6�i�v���e��-i���9�<$�.���H��>�`�G�f�%#yͦgA��.�^�Sl�
���q6�P+�L� ��SˮŬ����&�5��' <�\�����C�7��)�YyaF��n!��Ԇ��Bਲ਼�)VJ�q
���������t�fKz=���G/LO �FƬRS-���b�XQ<2�J<6�by��f�
�1?�Db�9�؇�e�61�=GHKK�,��(�L:/�E�' �sfO�g�!Sh���5Ux��Њ*�)5�&�N|��Ω��!��)}-m![|k猓6v�sQ� d3���j5+�!�نRT��M���BS-S��6��(�~����x�	`�S�H��'���<쩳D�JC�l��o#�SF�����Qq�7�;)�V"T�SL2��S�a N�&Jo��(vT�U5Oz�!�6a��X"�6�ؐ	��(*=��z~=f�e1d�;���ۂ�(�)�f���������?Х! <�2�`95=��e�i!�54�JO<X =��qu�M%��ea�D(dF��45ׂ�,|�l����B2�9c�rEȘ�����a"��\/���^F~Ȝ�	� \�.�[���B�pb���m\)Sk��0X�RӠ͐���Rݦ@��\" ��f��"L`~�l-{��^v��YH� ��d�2�����3c挐��l���7lE	k6f0F \oXqJ�'>O!`��?a� цɣ7�_���1k3T��˓�ee�����/���>�۱|���O+:�O��?�������}��k�;�n;�kj��Ŷߋ�iI�~7�����<:!j<�ֺ�*
�5:e��W7���*z�䐫��,��u|z�٤O,�_�{yr���7O��|���;�����w�~w��x�������\v{���;��Z{ut����F�A��ѱ�[h�Z��=�_H{}�#5%�
�-c����^�������ξpg聋6dk���>�JJ൲���8��qb�=�;?g��� y����K$�~����O����%��|2��h��}��! T AD�둲e�Y�hȉĐ�g���"M���n{˿�]mml�m�ڮ/^�6O��[���ս�����ӛ[�}����R���}���c0O���Dx~x�.�μ�z�)�("���8N�_R��Ku飜W{G>�������^<x�����S_�nӧN�G��|���ɗ�굧��H��Z5�Y�_�L�\o �f5~C�y�eˎ ς��5{��/!cv)�ƨ��
]�~2�70}Q�����o�V@����[?+��s��wn���]�%�?��a�۸��b�)M�����x��{�v������n/���om�|�1��<������|��/����[/��8>=9���̣M�q;��u�N�b�zY�����XN����)��P#����q�OU|4��K�M��@��"��yC���sBJ����������0�"8O=0#�>���0hs]�<M�H�6���CF��QikV
��c�1�K��S$�`�]� ��m��ԧ��22�� �KlEHF���+�a
�j��5�����f��ʏ?���4}m���K����95���Lg��a�E�c�-;���fՍL�[��9Qn����eH��GCc�Jv�<HLa�ћ��kvzƭho�q�,���L*����ɇ"�T[H�4G��y%J��줚�7����Sa����V*�|�޳�h�[]���JL����kR4�
C�E�I�'������,DZx/r` ��y4�D�%j]��r`��/��>*�t������|�>�ʧ��*�j�4�9�����Os!����K�����e��g�.�0Ġ�9�a��u���5��lH����T��q�)�B�>��S<L^E㧖'%U^��*8m�������_�*�@�k����xy���Y#Oee��#�|�`V"䔃�kl�
H��D��9J�|�.~6*H5�D(��4���`W[C���<�� ��088Պ`�T�N�����J�����P^E�W|�豛�2���>R�q�lJ
�H4ʿ��+ ��$*�Y$ԚҳMI�J��#�)���t�c5+r�7[�T	b
?��`��h*U �H�\/�TM��^GNH$ g� �^�R��R=�Ьtxв[���Z>�%���?TO�W./.Rh!�l<�%b@��=a5���#����B�Lv"a$5��!� N!zM
N��z!0����^�#~!0�cSb�Ԭ���V*��L��J��,DߪI��J���m�;a��ǆ�^o!�?*A.�^��<8c���o}n�/V��Ulh���EƆO� '�V��Z��� ���划-P����{��X�Ly� �0C�
 ��.�F�K��(!l��@ %x,�UX�&N)8�9��Om�	�	Э���;01 �N�H��ߐ�J�:�b�X�е���QC�Y��4�/��Y0Zx�oJ�!N���ζ �k�Pi�V!�B�#��b�a��.m$��	��`�t�i���vLyo#�(�1�rf�L![�)��K:��c3����r凤�9��0��1��#F/
	���� �lJF6��<<��E�*�_C�TU�T�b62�IBk��H��"C ���@HN<)�h��[<-���9N�&��1S���X��|��
�,/ ��XM`q�P+�<S�f�>Z�V���'��9�:Ҳ� �ohi�C N�`�����z-1� ��svT��,�>ٜ��Ԁ��T�_.XvH��J�?��Ǭ@H�X~3[��x�c�8�9Ӑ� z`~$���ش    IDATNY�I�0�4�Om4�I��`��Jĉ>=�����		&P�
~�D������R�װ�m(6��1��m��L�(�S ��䧧��aL��[6ԗ���㌄_� Vo�ze�J���o��0�3&�9�7�d��%]�x�$i]�QC:����1i�E�÷�2
i!�0B4����a��P�^@��#��V�Vԯ~�+~?xz1������[���y�c��<l�8c��Ƀi����$�²��h�4~<Z0SݲPq�a�l�[�\���3����$0'L�I��` �Ͳ����j�K
�u<��ċ-;m��IH��OCo?*Q���@����L�8SK���B���m*6����'��'KT0�h�lQ��o!��y�d_�s��ϞCF��n���G����Lj�����?5c֚�6LOl�c	�^r��b�Wj0�GI��6pzLIǎ�c�i�,�`�3��Y��-/��f�aF<<��7�f�f&uّ��x^��!�[S�*�����~��7�>af�ZbfF��t2j1�x���!�*S�	+
���ʫ��ب�5����`<��Z<����n�����H4F��r
Y&Ǭ�@��J�oM�vw6v��n��y��j��=.�9���_<;�͓�����W�,{s�[ o�����j<=��!�VzB������_Y���7�l���Wj�f��9�^�]�X�O*��T�M�4���d�������c�,k�g��V��_}�v�����7�~���O�l�l���k߮��w6�v��om^�������d|Ѓ0<�5.:)��D�e�9`{+���cVoi�J3t~H����d��� 3��NB�l��ek��J�5t���&��]x7؆�f��
	��x�0��`�n���x�ό^���^}���ء��\�J��+.,x!��`x�om*���3̚���경3�ɰG���8��ƚ��^�������~�'o�}|���E��TS���!X�����pԢ�7\�y�8p�kyï��D��H�&���~媨���Y�������_=������Ó��=9>qB�^*0���뒝���r�HT�����ʴM�-��_�q�=�<��ǉ��r,��1�'Z�4��K۸h�^ة���?*��/Ǭ_@ͷ�-�
�om^l�?�z������vϾ�����o���ѷ4Om"�뗶g}u��o�/Ʋ="�˞�Fa	��_[���.F�%�����?W�}������[�m����{On>;9<��8Y�ᅧ�o.�-U���Ce��XLZ�(�����(+�/�� �޽{>�ŕ�E9Խ�ir��&�;�`�����^j9��9�`������R���(�����,�\��[�^�b�
� FR�XNx N��O�T@)��{Do�u����	�Y���B0�F~�e~�[��J�Ȣɫ�+��@-01<I�at?�D�Y���|K�'?�	m�`fis�!tix�2�4�,�v6d!0!�+��c��528���n��Z$�d�L;~�N�������e1e_�ۦ�t8ݲm�)M�fO}�b��{5����)CH�z�f�k���5�l�!��M�[k��#�H.�?B��G�l��Z�%�H�$�>IΉE��Ӈ�~˥�i�!��hJ-D.��.y�cw�óy4<�T[�A¶"`ÇvV�ݻ繦��ԵE%��l8-Y/�Њ�EUk�dhV�YH�y�NR�f�#�l��)���ҨB+�)���Qi�b�.�y|���2�!�g�c�k-N�=��a�)~<`Hx�!RRlIM��
V���?�蔑����E�!��N��=9�F)֡�y��B)�5K�X�M�^ �SA[�X� bmI�Ē�a�JN��m�,��v�Z |�nE]�%�C�\��˂��/\���g��R+0;<�Bh�����@Sm�lSah�Tj�<�	������bw��V%<
Xv��F�)$��U1Cy���K�M�Fvୂy-�S�a�Y8�-L$�P��I�D�*�(C��z�Y8��j�	*FSR��ܞ��D�v��i;F	�y���-#�Q�����z6�)��u$�Y��j�F��O��x�H��/-�@ �J�c���	o�z�ԙ���r�W0:��Z�����(�z ~��g�SC�o�d(8���,J��يj�m�0䊃��)0'�!*�5 ��ܔ!��	��}�*��s��k�9�8�b�НY.����������z�D�Jk�$[�e�r���b��ƩG�~	 /%Jp��vHk�Fb8�0Jģ�@��H��T/�֫J���kAT���@S ��1��'�6k��vQ��T�O/])��Qa��-S�j�7L�,<*���,ԚU���ea�R:/�ՍfQz�Q����)/�T��$=��\)����?���]��
�$~lD*�B9�j����#��W(��"��x h��%r���"5�r:1 ��kC~N�HA��j��I ��i-���ӔS֎���`i�`����XC�����?Cx�I����(�m��q��6�����M��A.K�?? ��U[C�<��)R5C����fXj�`���0R`f�(��l�F�3��}� n�E	d�"��T=���:x�p�JR<���%^���Öy2b���אC*���1��)��ِ_,� \۠00d�ŀ�YTK�p�2� ��������<1�h���¦��	���<�!��?d��]�L񤍪��<aeD�r
�/�݊"����ov�o9��ښ� S5��pKg����GCh���jV,�ڥ���F`�	,D�J�H���%?�����zSZ�b���\�K��旎I*0�h�j]�q�"`��
�
�)Ξ�1�-�����۸5�@8<��V�!�Vj�#�6����s2PqN�,��3��%����y��҄Lìp�P[e��>*�`�U+�Rd�a)�)�<��x�r���zly�0�a����:fNl�`�hh�.�!fx�4§$����A�$�<�� ���rq����5C`<f�ek R�g��k`l~�`�<��xg2��m�S�(v���L6 C��:�!�v�8�h��q�:Q��Ɵ�
��Ѫɒ���4�$�x�4Sz�4����x� �d��5 �>��0�ė�ƼD��0W��*��(��9gg�������+�Q;(xIe�����G����<z���K?�Vg����* �i�G?1E�6�pJ���l-ن	�yM���)�c��pC��Ӏg��g ���D����$R�YN�l!Q��B�fG��nN~��� d*EΙ%|F�i��8��q�j�y`��8�w������~���[�n�딾�wx|���۽/�^�zyv~t�6ΛZ0�Oƻ��><�XoS�K��8���Gb���r$�-��4C�i�⌡�3��b�+� ��y�و_N���"�����|��p����7�����������Χ����w�<��j������������#//����H�闓JM��Ǝ/qR�b]��icvQe��H��)��h��K�,�&�r'�_�6O�P�Գ�V7�9�D�h������ �ٛ��&רּ��������_~���������������-}^�����`���ֲ�R>)y�"��Z�� ���!-��f��k:j.T��;_����������V�϶��ur����<��5�֕��z&����c����8�B�_�������ŉ�F~�9��m����?���'�O_=zr��h��g�/8O�U��N���d����9]��Uے�`y��U���손��א0��'!C"������A�3�?���˿5�t�z,��7�}|M�ҟ�<?=E��������r���6�߹�����v��X��ڳ�\E��u�m�'ͽP-2�vF�����s������ś�s����O����_=�f�����ٹ�)��_R��.�Vъ�-әy��q�%��)H�p�~��xw�y�V ����:�C�r�%�T�?���\1+u���g00��h���S��cV?�~��3��̊bX,��ꭈ�\��k8M!a/|�Cy�y��F-��.O�pw��,BC�ad�EN==���%��2��D�����s�|hVjHI�p��aT�:%ed#ԛ*�ޔƙa����JI25p$ɔ*y�֤bM�̈�,��MXC=�8�����|�&����-}	��`0� �M�����cv�X^�91i��,�؊�V7C~��s�u�8*>ѳ�{-��[���0x�f��8Kz��YH� |������٫�e��f�R�t2 �Y?�$�
'�(gIj���h��|��Fe]�[�G���xҩ�R�V�ٔD��Xf}x0��m�T	gIPa�O�f*�UX�a{���_���)����@32��\�z���#q�K6S`-� QI�W���&61l�\(�O�*�Y�#���?�$U,����`yZI6�v�\�z������c$���Ǧ�NBC{�G�z�ֈA`��Xr�b��
SD�%Eh�p�#Rl0�:(�f���c(P�r�ܔ���� N[�#/0�D�-1�14Ƭtʫ�A
<ai��>L�QQ�V^K� ���c`�dTm��cÏFK�m2%a�lM�h-A^-��28���F�����)
�^�x�@� c� �bk�Z�b6t]X��GRT�g��M��14! �Ud�"��<S$	��A��&�ʘ�I960Q�)�*�Ca<]��B��BJAs���h
Og&5�XT4+$[~`HyI�_괉E�l�y<�aT1�� ���r��0�,�� �!gk�E	7�G�	@���E����"�px�x~Ⅸ�Y6�U����PCz�֗�!�o��P.��zY [5��ΰY���[��*m.p!�4�n\�%rLA����)��ZCM�-�\icPխ�SRT��a���TFÎ"%��*+������j.\�w���6��?�҉��pr�%�{&6C��I���E���v��|$fEY>?~ʕ�_5�� U��%�X<z�vr�dy�*��oS�Vj=N�u0%��
��!�A������>�
-��A����D�TY�,�#�G��?�R���9��,
-X�ِ �56y��cf�)t=�S
���F�`�˜��P��{�!�X�j9�\�ah�\�8�؜U��be�ߢpj�½�*B�H��~�*oJY4�bЛ�\Y0 �W6B���f��굃��!�4}�r	'#f!��V-)=�.Oe ��G0l~C$��i���iJ,U%�����Ӑ�o�(�
K;�H�5vi0�f�G�;h�^`0R��R�G��H��J�Y��;b�e���ʫ'X��&;����!���9gD�qj[Hʈ�TCH	*u�R5���b��/�*)[�W/#C8~���%�D�8�`�g x���@�9!y:B��,�ZE0�N3�Jc�POL��ˈ߰t���?I��X=gr�l6�H�Fkk`��%��"�ȫ�@eI�,�����(0������X����/���҅����P{�U^l��c�s{ʃ��/#0@!r�IO �69�q�;�D�j��9�H�:�f*��tb��ɐ��\X䆉�W��d1�[�Z;60��C��AŐ�^�4�ޘ��1����(:�0^�DAvbi0�k��w*�y�4T�ҕ�'<ZS���� ?<���7g5������j���p{$�k����*�a�� f/4�B��i�[dᜲ$f"�9� �
̵0ڋ���[;�t�lll�`I2��\f9ٌz66���ئ�5��*Q6@�S��p� Ыa)L�RRK �yk
`\��� �x��Mix�"��O��)C�-$[/VH~CH�z̆�m*7�"��M�_jT5�^���(V�2?�4���zvlC^!� �	�l���Mku���6S�1��]� ��[,�,�n��3rß�`���v$��0Kd��&,��<���0�R�edDؒ�����F��9���7nlno��~c�CMW���ƫóG�^=}���;��O��k�O]*�(+y���JKH	��],]^�钝���9�x8q*�
	ݍ����]ZϚ�/�<��
�X�����#T���t�I�����V�?��������?�?�����o����n�铽�/6�OV{�;��׊g���^j���!���'�U�M��*9ʰ\bz۱���kI���� {�_6�2��30�ƞC�ؘ���0�/�x'�ņ�����D#�Ы������#���
Z��Lu�����F��X�Om����D��pz�&%�P-�+�����ʯ7l�B�a<)�GY����K__���W�o����޽���jo����*][�vR|��S��?_?�����S�L�oHU���:m�'i�{ ��_�fd"�_A��i	��������Ϟ�>޿��������t�O��R�~k����r�3T����miz�e��`kM1*0[���$�S�>�~��9m���G�A�>��+B�������Y�z��D,��S�����������1�?X]�u�t|}r�wjqw�c+w�g'~,q�n�B��mlm��Z��u�/xny�|�P���х�����ƭ�w��~����䫧������O��x�ݸ�6�7.��ePY:W4Z��u�����f���мt�a�$�q� ?-6�:����wu�e���g�	0����|��
t9�'r �>��ɰ���Q�!�`�Y;���f��&2�8���� ��]׾�����[:�,}^��$+(W}7���Z��6�-�Bk!� �g�s�=K�8�2��U��������`�c��P"��$��!���J��kS[��Z}`�B��wT��,�@���}��L����4%DoJ�֐1?�i��mw�B�����#i?�N4�Ϩq��@jQ~�`��1L�ɰ;�f9$0���P��D�Ob9�hȠV:G���|�G!�`-;��@:u��������uTU��ɣ�硽�}���>��4D�2�[��`C���A��
[�Yy��ٕ�Pj�2�%��c]�
1����=�xLaH�:X�bU��RO�)����\#�İ���!U�9��Y8=b�Շ�!�v
�(Y�	[Y0i�I��$���?�fe7�PO*r;��$k��;	�����WC!�E9QfUƩ�LT�܍���p`����D�	��T	�+�W�$��-�Y��eDK��V`�sJ��H���IWќL�)��Qb�Ƀ�څ�h�4�J*�Dz~�A��R�:E��F��r ���"�H$<�ϰj��Պ�t�))�.��9f ] v�xI{5�=a��6�%��by��'�0�M��I�B�Y6Z�٢�NyD�ꏏ�
Ue� L
W��렖�	�D���������!�<�e�A�N�V���GRŐ0x�+�^8[�ސ�� f�iȶv���#���,I0!���h� ��B�Mq��+��<ˑBjlu��KƊ*B:MU��8y̶ƹd���z{�V��
yͲc 	RO?���% H!y�`�` `�<��v�e����Y��-�\VM������X����Fp�$W�&aP��^�k�D0b-�-�m�!H=��?�Z�H��Sh��:Ң�9�f9Z8N�R+��fV� Q*�bBd�k����ұ�B�
P+��H ��Ie7���>���"0�D�r�V�RG)EY����1ԃU�d�d4�/�_Sg��,6 �m�1���z��V<��X�Bw���j�-��V���ڔ� 8<�EH*6~k��%�b�fE����-o˩Z�Ԙ"5��G�U4�`��:cH.�t�h$�_��_r�갱��C~��H��׷�"�%�D�W�.�;��i-޷K�Ҁ7�*(hX������6��ܿ��]���t ���G.��h*�s�y���Q�z!�xH���:�*`���6���b�q낇��c��ìb�Y�潇(��q����I�ng����'�h�!    IDAT�)~w3T��E�V��Q1D�*��� �TQ�o(�f��8���6���F0��<^Y�3ܒҀGa�lS)��~lr18y �沛��l%JU�`�� ���Km�ǔ��\T��� lI�0`��3� 0�)x�l�Ӕ���G����-p�`��2#1l�lH-@<l��ճ�M�,b��`}��<`��X<�XC�W�~V2<�6����!�'��Hj����u&e��֕����q���L���m��Ǡ�r��	7�`��L$���Z,�S ���/�??��$QD�4����Cz`l�>~� Li*>g���E�V�[��윲;lSD�c���g������,�0�L��C�YS��G	��	P^Cy�Z5���`��zCI�� �B�8.p��iX,*���y�5�؄a�7tsF 1S0Ol��0ج��̓�Q���������C6�Q�$�L"vy��ea �q^�E(X��G%��&L#lr2���6[�^�`��agL ����r2x��h�8�CJ��ca��1�k0b������0���p����*\�<�-��%P��`�ٌ���3u�͖1��x	cL@�x42�B���:d�D�(W!��5e�kl�d�n����J�^6s������-%�_�b�F����}=)��0@�<������R/6pz`�k@yVƆ�K3���s����4����,pmwg����m� gg{g�W�u�o}���O�����/�_��.���.O<F�|�ʚ�B��� ���������Vamc������.�\^ |r�*��7�^�/K�g;}mN�u�U6����}�k��'�k'k����7_|yrt����������7�3�}�vO��8�x��~vws�˽��'�*��c�j筄������-k��+&��.=��ܷ/]�<��Vg�͚�m�<��mr�K��V.�fq�K���W�Z�`�� 
����z���7�^J��\?/��G�_������C-�Tj�28)��zZ	C��`l~��1�O���z���y��v���^�<�Ӣ�|xws�x��po|�֕��3R�9�|����j˟�<=��=�T���&{t�d����x�Yvr��7O�N|U��d�����/�zq��
�N�E�;�k�:�ϨI��v��/R]���R���Ҧg�{}�4SlNv��ԧm6[3���83*20g�x�j���\0���Ŏ��������{�U�w��8/7��|.�b�=?9y�÷W'o=���:{{w��ݛ�[�^�
l�@�du��_Cl]�-��BY�百o�a��[�7��s��� ��o��X�����]����X�����'O.��z�����ӳ���ӳ�͍����vyV@
���qD3�%������?�����L�p+&�|Ap�]6�Q�D��:�d3�2$B���&�|����`��� �dKZ^�)�fV_�5��l���!��15XC���0��Yr�V�A�'>D�;��V�@�Z�j��BU^���<�a���0�$ ާ<~(��,���������Њ0S�7�.v��AF~-��l8�z<�6�e���l�0�bm��P���jf+�FR2�R��)k��^�x�S�ƍ_"Q�m`Qn�n͘M���繎\�RE�;�SW�jBr�4$n���>7�
�(�G-6!l|�$�(S9[�Y�5CxRy �����I������k\�D"Q%b� ����A��Z�`|ȈP�"0�z�@0L�\�I�����R$^���|V����8��M �(}%ғ!)�x��3��f)���l�q�(?*+��IIU��7�0��lOcP.�B��!Pc[���"r)�'fE�vf.'I�:I|)������(z ێʋpQ1>hsQ��T�|�X*��>_~��^��iDRE�*�.��B0 #O'"�2���F0*k�
~C{�'0),��8�8K�DyRB����2
�J� WU�b�
���CG�|K:� �UW�i�:*�Z21�=�E����gq��(!�E1��X�j�#�K�'�zy�Y�^�U0���d`��f�������
��R�	&��` ��+���q ��*��`9i�J�m6����ˀ�I���i���ˈ�u	���SIK�B�E��
�A�(ăP
0�x0.4N��kV��%�C�$�4�m��hy�s�m_HE��%Iz�5 �-T�l��Gn�if�J�%�J�P�dl�M%�*l�ͪIK��E�b�s⡁0�c�&S�qJК�9�3�[���� "�	\.�
�*I��R0��&�A�(Ǐ3yz��]��LA�PX��x0�h����D�N˼��$Ux�L�X$�h�菙�6C�6�X58����#��f�Iu6+@kOa(�wNK��[bXY��!��G�)��Kj���a�'��LU���Tm�_b���X��.GfCup�$-<����p�*=)�C��(�zʨ�M-�Nxe�Yb���h!����}��f�D�`��咢t<ֈ��L�e�-����l������Li�k�Ɗ�SK�\^7[5��(:���t2M	�ŭWR��A%Pv-I��-<� ����b�ћ������*K��+8I�7E 6=���tHx\kV�#֋�;1��\zG*�@:��~Q�S"lV��t��PRy�����
=yu��b����:i��*�<؀�/@K�^�����P��� �$�b�I��U�ͨ,�n�H�������xJ���������@�)�$�3TY��K`h�~:٘�S.�<2"��TՐQ�ڽ�E@�
L���2������0�b-Jx0I1Ӧ��:�}O*Nl���B`<�d��I�ֺ��sb+\F~� �7 e�<��-[C��FdYJ��Q2�b���Z�zz��[�,���<-PO�)� v�z����T.䉟��ZH�8y�/�WOƬ��5�H�֐3����"��j��S'�+��:�z��R7�8������"LK#���Đ�P+��R�ҝ��d��EM�!��]�� 0��H=H,-ͱ	%$f~�E�P�VlRA��OmQ0�r���!s�0xb@��!�R�+ցD� Ş-ZS<R/��6<Nβ�\N
�e����ƃS
K31�4s�K1�04� lz��m�D9��rJLQy85K���}�T+vJD�Ղan9�p��e)5��@fÛ��kh<�1b�,/��F�)$HC���8F�3QC�H'�*�64Ŏ��� �B`�dCT`U��<0@lN)���&g��S��`$� )iSl0j�+OHTq"�d$)fC!RGC�"�D�i��-�z����|W��08�f��"I�a&���Q!���e'�_�Mq����`�P XC��h<��s�d:ۗ!eIj��%������9��x=IJ��G+�B?꬙*P�J�9�斿!���8$�$!���>���֝7V�[�7o\���x�֛�����g����G_yM�/�;��@���/��ʗ�����e�Z�ޅ�#b��rhs3�� P�"[�bߤ�:Hc�vؙ��K���_�~�#v�����/�z�b�6�O\��������=�j�p����|��n�|���խ�����e>X��>�x~~q�{c�;��
+Ő�&���h=����L�fH���cE��p�uD��J[�f���eAW�ަ���t0�I�뤁��*Y`xL�{r~/:Bz-���=9����+I�^����W���޽{�g��{����M�f5�
�gK�k0���ؒU���I�)�k�G7n�Uɫ���7�{�'����^>{�q���zn&V^Tx�\��;Ίs�i�|)�C7�zb�k�G�㽔��T�+E^P=�|���ѳ�/�y��ӳ���f����q��ˋ�U��zȁy}�0�$��<���*WN��`y+`�]l��Q/<���Є葘]W��H���Hl!��.�Eې�k��P�����˗.������<�]}����;�ƣʍ�����֥_a}����!��Ɠf���B��/���C���/z���z�96y�d˯����������7������>|v�����O6�7JO����._�K��wf,���m�^������_%;�>��s���݌� 3�]G��w~������Փ66���6��MilNY�jC�	&רﲭh�4LF �`zN�pON�������hfcn�-��C�ϣu71�4�)ׯ����*�O�T�աz!�j���@C�I��-/�YSS6����>�����S|�D���ƣo!zx����e���H2��zC�(o��I0��)���i-�c̬�ܐ�W@�Bَ��hD96zN�9mA�D����Ǜ�~����P+��>��>[���d���M.��\0�Bl��~��'�8�d��kh�)5�k}��%�_v�Ô�L
�R�e���H�ph_|�?���uU�}"UҬ��I� IǌѬ�R��q��=q��K'�<���<��;	����k�0X�^��^�6�`����X���u�x(�o��o�&g䡐]#Cx�A�6��DM�5H�_%a��{�YeL��_��_�؎���BQ�l�\���$��;`�\�j�;��: l��pH!m�'���N������Xbl����߇�}2�ʡũ UL ���*!VaE<��T��f�"X�W
�����ac���2 $J'����O�D�̊�GFN �f��z��,B0��8}�i�����[i�5wV�����0��� +����.�lu�fh���Ԓ�s/cL0�!L��:��(i�BX�,�5Z�)~[�e̤*���}F���PI��8���4ow�+HQ�Ȱ4�
f-�ih!�B4�-\}d�74� -@ҿ�H�F��R�L`H���,Hؔ���P^�0�9�e1E��7kubՁl̲XHkn� ��N�)�֥n����/Q�bh<m1��Ў%�Q���`�WF�+�\3���!B�B�I���� CT����9���`��Θ()��J����Xl�+Q�`��R�̋�> ~M���P��+H��1^}���_��lC��~��*>��.�MPk'B�<���YWJ)��	i�+����9͊m(����p�3�!!�bBj�z�ף5%�M�:w��«��-�-
�&��N	�έ���>�N�US+J:=~��1�!���%w��M�8m��1���������M8� rC �-���Y�����l9��)�Y�F1d�G�p0;���j0��)w ��j ���*f�B��uX�X�&5C��yQ����'[�KCT�p��b�(���U���֐T^!���0�؜dHݳLHN0~x�I$�ں�8m �����z� �X �Y�N�4�f<� �Q� x�$�Y,�9�pxۭ�.~�%�\c�#gC�AQx,��@�(�-W������Ea ��q�B��X��diw�8ݬ,�`E�ڥ�4�xd�-1�X2�Ҫ�Dj�:�Z��`�裏�r� ���}ɔU�)��8�����G.H�	Ȱ���M�C2�o�HHoul
KV%�01PhV81�y��Ư,$ݻw�����_5��D.@ã��0;��`�lxR��o!CHu�#d���V�a(��}�ʨ`�JR�I��[�Ea�k��I	���s*@��y���$<CYh�J�PURJ��Y�{&�Z�Q��^FQ<0ȥsZ���5�0E$�l�-٢R.5r~��c�'�K�� �B;�x�`���%<-������l1�D-0=r	�P���;+!�\f�`h8٦�ͪ��
.)^��!#?'1�X`La��2k��B��Wβ6,�؜
Hb<Ԛ�(I�VCS�5U��H�(��>N� ��4�C�Y�5ţ�ά\��l0�l!�b�[f��S�f1x�\�������/\��V�-k���/�T��"74\jR]5��8SNO`ŖT�ua�F��<�P	H;#�ؤ��8��B�6��3���x���T=�W��	S,N-�e�f���z��M
$$Ar
���%D �ud<%��1I2 ��l��Jٕ�������))@)�̂��P`������e�Q�cE]M<�YN�1CJ��Lo����$U�2�_��U��)��<�.C+�Y@�z)�[��l�u�
��ƟF`T%�T"�r�OL`�$T���Ʃ���$U[���<S8�u�e\�����[����t�k�n�\�}��G�����g��%J0��V��<)Liˢ���h)����d����V.���a7+* !ؖ
\9C�r���#��U�[u�q̐}u&�~��'��������?����ӿ��;�����w����:X_���j�������K��t�h��O-z�y��ozO2������~����
\��t�4[;�Ŷ��7ձ��KR���U����~'d/��ce��z�z�����V|���ܿ��Ro�s�2I$Z���}Z3ީ�l�[@�4�Х�F�),�04��C��	�&��8C��7��Z��<�^��&��-u�G?��xv����s���M��Q��mŃ��-���ip2���S����߄<�K����Z'����e�H�'��ӧ//>����߼xvt��b}�'u��BU��{�X�r2 8�r,�sɌ
�h�:.y�e���V�h�3#;�z`�l�r���#��Tv����Gj7N/������|]��T�����op�<�ru��z����޾�OK7�W=o�nn�zS��vvl;��dO����q�4������#���t|C�]ă΍=s�rkw�;�o����r��|�h�{��ˍW������7�^�[�,�{�t��:9<��В<%@λ�|��Z򃖇j���_��s��ŊB�8�%J��w��ʈ�!��G?���|E10t-��`��6M8�Y�ؖ&Ŵ{�,c�P�3da�,�(���#�!�a��>��O�>����/����u>e`[�z��L=su�˂�0�z������{��# ���#h�!1����r�3�d��KY�*31f�0
���f,g~=?�2�� Q[�0[�Q�������Q7wUG_���SdVU�ʈ�a�rlԼEy�!{7'���H��e�����S:�a�f)N $?yhy��o��CM�,��qb#@:?��)ڲ�Y�s���F$� �:�e�g���L��p��,6'Izi�В���]M�jV�!D8xQ�#����~�)*/Q>�0��ft 5� �3�j�c�5���1�Z��>P`���/�#�%8�<U����2V��;	�Q�$�i�بC��z�VlV�<�U���s��9I*P"�ER%�w<(!Xc�C��zNo��������(�1+`!�j�Q9�y���D��y� xŤGF0kq�d��ً�bd`S�P�:@�Q�0����L�)���@����@�,�5Jъ?���l-jn+%���� `0+�O��O��;��+��X`}����D�tb�ڔe"'�b#��-���oV8%!���3_��Ha�uY{=������U��H��B�1�w�W�v�0�V�o�����c&�3U�e����BC��e�Ĥ��O0m"��sJ���VZ*z8U[.j�C�1tz�:Nx$r��aP���'�fuh+��m
B���`'�l)����`l$�H��y�/�h5[��k
�`�7�����=N X����vSh�0�A_����!�z<9{y��k��3<ZldT
 I��"@K�/a��7�(H����<z��4&�>"l�-����~IyK�K*\Ҷ>*�*,�3��4ː�*v�V%S�*/�\�B����O'�,��Ѡ9�O��(�\���pbf(?��$¦OC;{]�p�z!�:�i��ɋ_�7+�t	Xw S�I�틡��A�ĘB�6��)�R������a4�t�� @s��8��KM�X�Q�&�w�b1p�B���i�)T��b���Ή���ۑ��]/�evm�"�_/�~̪�ߊ+N�j]BR΃D��H����ٺ����[    IDATɎ+��UY[oTSI�Iդ��d[/3�؀����~0`#�%�f KbSͥ٤�4���++˟�����2p����%�޼Y�Y�3*K����ly:x�O&z�`#(�H���-�@�C�$� Pb3�N���L��a��"0Ʉ�K�%C)��4��Dli���Pu	D�>P�%[��J�|q����QCE�j����������MD^J�����+��(�t-���U�d�\�,k.f�I�# *��f���	j1�`�B�)UL�L��Su��1�h;6N��dbF"�~�/ʽ.�h�3��,.��LSJ8��GB�j��L�]2���+�R2h˜W��b���U���`i�Ő�� P�prf���E�7�x��IR��2dXPObb��B�\��0��)%C#g�Pf�,}Hrсi�3h\��0�ǛS��00^A~KI�EN����MQ$N&���!���B<�k���U1_��KfzC���id�4�}����%G5JI&FE��X��@�Q�.q�P'�;��@KI��`6ʡ* J`��,]���&U0m�F�p9m:/�
Oɱ�F/=M�̊AK�s�4xz(^��2���@0H`�J�0�8aˋ}�`�h�Q�%�� �a)n��%$6J�%�9~J�R�1t�F��I������_z���T�R҈c6�krz}��R7�B�E!K&ߖ�hA"����\Y��hp�I��������c��T�4m<�����`.��,ɂ��dˑ��.Q£�U/���.�I·��
 nE��V�B�K`��O��K.ׇJ�ܙp2�N�K�њ�`��c�I/JA�Fz$�F� a2�L���&?J�↟��@��v����K���$S��dV�A�a��S.�'��
D�3���\�L�����rf8�H����1�X��b�^�'K���c9����$cVt��xJ#�J���u�2 ��e�W,3+w`KY�9z˅�z��hV��+f�@�*�rk�Ȭ�ƿBb3 k��K2w�fBq��x|�q�e�o�)�`�_(�s{ou�����ٝ�/o����?������q�������!����
�I]*��4J�	×2��Q�0Z�Q/�R�5�b.�p	뺜Vߥ�A����u�#"�Oe�o	]n�~6Cy�9��/����o�s@������ͻ������wv�|������������W'�o6�G�7��ܼ�M��;{>M�IXQr�|��j���
X]UA�T�O���Q7�єq������ʍ�Xg 7d��.�T#/�^\s�"O[�A���O>���d���O���^�<���h�6O�y��JP���2����R�0�o������G����'_~����\�,�U��}��W_��u���o@��d���~\^��9��GtK�����i\����4�|���.|GЗ2O�O�.�zz���˿<;�����~�ͷG�����\=�P���O�*���8�_���:��CP�t�l�-ד����� �Դ�q��b3#�*V=)����q���lF>r�y�?X�/az�\>��9���=m����h���ݹz��'�����k�{�����7n޸}����<���sl�<���}.z��z�v.��WdW;�����W<wVW�g�[���>�ܿuq���kG�߾���W>�޽��?���E�x��ݯ3�'����v��Z��N�����pC�Z����{��^�rovb{�����73��0Nϗ~X)��.=�H��= Hlpɧl�9���`M�.����EW��IX8�)��a���r��2 v%rGEV����������(���ƫ;r4��#��~�JyW���-=wQJ�м��J>K)cZ8�|iC4�`O��g&KO2�_�2q_��/�|QX��� �9�X��z�W���o5
?�v�o�7�����Vi��q��x0���[0:�u���������T�l�4�WP�6o�;疼 X~x��Hf����h{�*�TŲ�	�����,x��JrT �(�" sWQ�(#��-rJ�|V�v�`L�Z!��,I`? K �4e�f���	�A�3k	�/��s}�W���%���</[�`�XRh���:�W���G&�4f�B�'�L���&ê\��_Q׎[�"�? ^�Q�kk�1Q�b �if�����{JT���u�/�T�-�sd��Q�f�vA>��e�=`���/L6�6 	"b �`�:zGTc�53��o{�EtK{l)�L>����,{1�v#������Y�*Y,A��u���z\5���Xt��êè�3a<x�<#!�!-P��A��ЖJ�����C������+�b��Z[�J�r�*���?6$����H9�7�  �i���N�t��S5���8�AQ,A�9����v��Iq!-��&#��cs}�΅����j =Z�З��F&������rE�ӏ�c�b�h)%KB����茠�Y�u �ӂ�ULJ <~�rg����Rb�����]Z�'X[���:<�����	8���k��2=��6�������;	r�!W8��ˁ/ ��Y�����L)a.mX8xVK��;��)����|���3�����N�(�����@��R���Z�G��1G`��H��������!�8������b ,�ݑ!��PDV��4f��q�b%4�jO	P���Y3�ͨ ��	��f�L��� ^D���3ּj|7��]eu�� i�J� �LB��,�`&��D#�)����kk&!�lstK)Tjd*rkP�$U
�_2��$�1@��CIC���,�&K^!��`�q��|zH.�dn�K30_z.�E�ėI�Z*A&��Q8��B0���ٵYuhe��n,4B,�_�B8�*0��f8�[RJ��<9i���.��ƒ/@t3'�<�+ ��������+��M��Ts�q����9J��i`�9٠������6�H�f�'p�Jo8��L�JX>1��/eEJ�� U�E�ކj#ݶ}�p�F�(�
�z�(`ȱ���Q܆p Ņ�l�F)�
��li`�,��f�$�f���* �#L����]SZ��I�B>�fI�R�ł�+�$����Ɇ��RP$^��֖�=c�$#+�D7j���Q��`�w-�7^:	Fc;p�v$�&��XQ\z^�N�nMBH�(aVIZ����	rS�-.CJ����EZ!%l�m.�p�8uɐ *�h��)T J��;o�����T�����D	/��/��[�A�xi,rK2�¹�-�6�%p�K�8J��#���	Rz
l��B&u���-�v��W��÷Nz��ou�5WZ�*Q0`V����0�6�ۋ���FNo �@{��y�Dj&��$	�H�4r���d��e[��=�=m��a�TZ�(�����&T�Ȋ��R!40i��I���%��� �	�̒,% ���]Ply8/�9΢ �y`^��C	6|�?��,��ZĽ�Z�^x�^b��u�	�|�`�"��]�L�~�?$/U05hتq�Om-����g�ѐE���Ҝ��WTq�i`�e�Y!��T�#�1�R�R����dV������r`��L0��9��(Iz<V�9@���a�j>}�٨'�	E�(= K3/�d�۲)d��|�e�����c��Ul�N1����fT��B`�a2���Å���4�Yc���;=�X����C��0fC	�ͱpL	L��+VT�� �0�8�*
<=$e�Ҏ�>@Vs'**3�2k��GR'���gg>�����ڟ�i�������;/������[7_}��������ǟ�_�\�]/�ۨ]3�%�sJ�^N��aʧJ��I5{^9�גW�d�X%����_�Z~�.�=aj��K��wG>u����X�痫���?<�����j���͛߿���p����[_���K��W�>x�8�����G\�뻸���8rZF��������;?6��Fz3 0I��溴p\�P���Z��L��p����e�p�}���Ս�/��lJ�k=�O~���~����C�ݾ��i��x@�8����\��f��M��B���t��f�v�z�Փ/6$�gogu�7}�|�ǿ���w���V1�M`�j�qs?��m-��\_�I����n��8 #G������ޏ��N��O/�����_^�o������'���+���TEƉ_~%� Y�$���X�c��r0,��4x~	?a�5$ � �e2 -$L��s���F�9��/�W�9S>׏�}��y��[�g��Uϻ�Ǜ���g�}�#{7֛[;�����L/O�V.���r�G��ЩT}'�U��l����&���ҟ��V�N�ѾM{Î�v�������F��Ϳ��_������]��ٱ�����E���KQ^�{��^��jHς���9~`=�ge������/\l�e�c��'�3�f�z7z@��quHz����|���xF��,g	p����BJ z3T]/���9$w���2��o`^|K�oO�c��B��gP�*�E�D�K!��:��қLo `�<��-7V#<eA��`P�av��4c��99 �ٜ���>�WWs?i-_Ԑ�@bg�JP�w2��s���nP��Џ���ߋ�Q�ꬒ�xzv� �Ҝ�G!4��鞞{�宫�}0�_D�f�{B!$�J�F� ������^I��H��_�ʴ3����4�����Ul���A�'�\Ȓ�5���u��YBD&H���k��艋�-0��#4{ǨW]eQB�eK#�4���� Q���@����^~`wt���?�yg�,a ��#o(��-�F���i*C�<���&(e�i4�I�E���#�p_M�(���Yb��Us)�
�����!iȆ� RrH(��n�	�JCFچ�9��Gܹ�6�?��(1Cb��i2$��+�p8�e�ia����ÒQrx������Τ �ipriI����5�˓�����,=x��3.^������KX������1J ��+ʧS����5�9 �L/(f�r�p&7i���*3��'C��.���սB&\$&CtW��`,�8�����;���b����$]5��= zy"�w����(nBH���#ɏ?��!	���W�=/mgeꢠ�	�Jɽ��K�x(Az.[�a��XeJ�96JQ(��
�nR�I�y��%��K���(e�4Z�ŏܐ*�� 	7v�f��W��}�]�*�uC>�=���/��L��玄6V��G=a/(d�#4ȕ�%�v�6$Y���$�􄓿~J��Nb++.b�K�ҾԮ▰��� æ�4`0�
)Iry���'�@J�h�G?|�e��T��)V�!�4�� ��Ez�^Δ ʇ�kIig��8-f��h)M�Vgf&���GfJ�H^R��Nw ^m����VѬ]"�Ҙ�.� 8u�#ن"��"��Y	��+0J�̙Q¨|BS�d�90z$"���nfHh ˬ���vK-u ��%H�L���A���V�HiXJ�h�Q�ѐ9$_���ޒ	�˓�f��0x�3�h�%|	�x�b�	 }�H(��0�`Lf&��	`�E�&���j 	��][��䣐�⁤�Fr.mB׈�����C���	Z�0��K��=���� ���.�d���.q9*gx.vJP�2�,�A����.Ki�'d���#0*KG�a�GuB�h)0+*	� ��\��5\�K�u	��6~�wz T��	��6V���2��C���u��!uL��t�s�����8��pq7+0��a m�
BF& ��%*�6N	��r�)m;B��.�c 6d2��Y�<� =$(�.q0�FO �;?��\̥���ÅR�Dh� ˖���.&.K�A�p9��R�I��˥�o&2L�2d �V	�m(N)��I���@tɸ�R����n+��y�c��!����X{�ĩ��p��P���_�Q�*e� �B	/�X2F !̬*e�F��@{�%��.�w�����m�7M��ĜdT-QY�'��GbvV����qx0��#aQ�z7QO*�����a��y*Do�<���T�҄c�y����ϟ>�W l�ɺ�����v_J��$�6�����֚��K^�uJF	J����PV��
 @&H̖�dJ�$���DV2G(E�k�A��ҩ��D+p\��G'<��^,�4�p��`����p3��
X 2*�dKzQ�i�6���I3�q�^��[ɀ��2/:~� z�(='�Xt�LY�?0��2s�K#>�,,	 ���e 7$,e)��҈�o�4��E1#��9}�����C�$/�x򂏇��-�$PJ�[2��Z�'���B���$�[�6[���dEk��0LF�eB�2Z.Ƃ�~"0ϭ�l�	��V���C6�g��i)+�i����Q>�4�E�� ^dle>���4�-� %3�2�U�YSϒ��5Zֲ�H_2�5OM.�U�����|)	h�'�9���9Og.f<�zC-i./�_չ��=����wo��[{��n}������>��/����K����qrj�Y6��!%&;�~��ƨ�����T�f�(�y0zH2e�4�y��a����Go�A/�8K?��ky��R���|k���w}�no�?��O��Ϗ���z�ww����;7���|��u��	�t*���t��b��8e���܊m���$eh	#����$�$��#`�|�(�7$9��u �`fm�,.=M���1��:�G<��pxz{]i^({J�:�U���w�<i��cƳ뙲�m�<i6ry��v�<C��!3H��R��IF#����5��N=^-؝��]�Wv���{��+/}�u�!{�9���6�O?�G�۾��ϼeG��M���+��s͝ՙ��*�rK�SXَg���g'���o��ώN�����/=-���̾=7M�R���M���l����i�h���>X��-#�XYc0�%C��
��5���a�bIn	C��å���ʱ�`�_v��Z�9�/}�sup��'�ۻ۷���<9����f�	eo���˵�O�}ysI��k����X���{)��lv�/��q�m.N/N�6wn�<޹}�~���y��滟]m.�|���ʆ�c�<U�D9r��ǵ�5Л�jT��n&3��<G�����g�O3d��LΥ�l�a0���P(�н��D�$.w�� ��;dט��vp^ /fˤ%��!y����	��6#�����07�2 6��<�_b4Re5]���X^=
�P+%z2px.�}�]F{u���� a�E�JА��PP�Z�4&Tb}�"2��D2���u�8���e�4��zoZhTD�4z�୬c��ңG��U�fjv ��B�H��9b�������A:x�b�����'�x���R�'�OD�w�(E�h�<+~������n.6��8UQOd(��5Q�|b�j��.\�f�
j�D�F<1GB�'=w�5Y&!�ݻgV����[�*ӌwoo,�
T=w.L�L�̳.J�� �om���+�RO�e�i亖���B ����3_�|<+0�[�peX�6E Q�yYJ�YKۧL�&hA�5��K���e{&��L�\&��� ð��&G��Y��ܓa$�W8�9�Q�Ux �U�#޲5#�wL ��dK���E�ќ����]bL5�%kY	��^��9�	+S�� `2�d���4��Hcw��'+<� �1(M`4�Ӄ�s�� �а��`6�;~��	�#=���Mf̱1�C����T0$6�� H	�(E�)gI�e���	�G}$�(��-C�R�.���Y����?s�fp�GkI��kX�Z��$r<�
G�W=����.t��MW�4�Y��ڻ�:K�+�?��L��=�b�]yZ�ڎ��$#���!��~/s�ʭ["'~������і|@���K�.�  �Ex�N�`j�X�h�d�2ˁ,~����H-��� �W�	~mN�'k��n�"b�w�DNI�^����c �'    IDAT�Ǧ/&.Zj)O^�`����RX���q"�1���\K�}1a��:lB#��U]L�k5�r� 0x^C���8J�`���\!�
Fh T^�5����5�,��^2xd�Pah��ʇ�"�ʡіL���Y�y1I���/f� d�Ff�t���a���L�^|���j�%f �<��)�
!�����4���/OG^�:0H�rH�j,�f	(ŅA��BK� (zi�-�X%�LV`M�$Glr���%0_x	�&(�9��)����	w`B��d���e�l�)e>s`2fɮV��іq,[��&70�#�T�{����ʝ�=���U�JC��	@A%�ؐ#��F�I�J��Z2��/C+�@  �ySA����bȖ�ޒU�E������4׬|$&��K&G�u3�0���)�]�Ȥp�d(��Lj�L)Qr4`(i���?��2�o���ƙǏ��	 R��n�`���K �e*V��%�' ���k��C��ƄADHi ��W:w�R�@h����I��wEq�\�ei����^����&�6��J ��C,2��D\BZ	`J&K	�H� �gK��̂*���E�MW�ӨW2�A^!�F>�	�`�a��_Ed^�u��@Ku[P�ȷ�,UKQ:E��*+a��������K!/�e"nT�匊��Y.^^Le�ڎ�1��� W��
ᅓ�WB0B8>��F�W[��ѪT�ȅ��j�i�J"�fHã��#FE���``���]0��G"�E�W��¾���(f����+�}�	K��@T����T &i���$ ����0CzQp� ]� ^�d���TT�:)(_����h�^�h/���lB�\\�4�R����f!�W]��# �e�dD,(+Vz��E6:9��fiC�lG�3q!��3q7h��
.u�U��mCG�� s,x�6ED^�M_�����s��\��1��' ����Ȇ�z����巰 ���	6$9��3���˱(�� �WY5C��T	
��H �Ȭ�!q��1�4,����)�4��≙�ْ�0$漄&��(�H�ᕲٲ@�ӑK^�`��2��b ;B � �I,O3�v��
/g���>Z3LH3��Ib�"f2�̥� ���0�L/��,�9�HBr�d-9�1�`*.09e��p�Yi
M(4��欨 Ta~�Kx�*â�xL�x,��be�����2�ܙ,)1��˞2q'3�9b^>���l�V/߽y�����d|��٧'���/O>�����wǯ�ܺ~��|�fY���=n�k�h-[��%�JYu���
C@f���[04`Fr�[�"!�O�6[~��(��Fr���u>:��OX��ы݃�g������ͭ��W_�����f<x����~ở>����ܣ���6A(�5�S�BmeiK�@��3+%P��� `LZi�wyR"ɗ\P�@�p`b��IK����C��$\��zG��=��^���l�f/����I��g�F(]&�Yr�KI#!2��X�^L��X��Y,g���j��W�������0��z�5�����U��M��g�6H.ΌS3�:~���w�؀ոn���O��c�.������t��x��h}xr��ݻ�\��a��Y��e%lF�ި�`3d�Da��1a�9���GY+^tY�F�`|Q�� 32X�fK.3Nʖ<�t	o���˩��/+o�����ӛ�q��wwV~����3_����套�=ٺ}������pn��͑�?s��:0>���� �m��J�V^"�G�76g�������{����o���7<�޹��ӏ>�����+��2������c�Q��9���<�.�z	�/O\t�U�v�+�gD}�J��/~��w�?����1�<�:$�
�m<�zf���s�GmrGHe6�e.yr�����r`e�F;[9K�0��:3k� �8ߔ`�r�2��Ќ�Fô�����3�8��.�8{6�/�jg%�Г볪=��#���@m=�������B��Ti\RJ���A~n9�	���`NO��=�9 ���R�g-�%�-��T�CRhǃ���t�s��NƑ3h?�B;?��K�>yw36V�X��g~x
��9�~��ͳ�3	@�-?�LoU���`��H�.�^BTGA����M,H�(�/��p�	�J[���	i����x)�l�g���\��A�Z*�zaQ��¹0)Y�K	C$�K���߮e�/��,ûA�� =N�͖�d�~v��A�m���G�2}VD�	�K��2�DD`�xa(����D"�7�Bh���"4���F�*Z� �`�F���!����@4�ZD���V~6'r^�\�$f	c�u�h�t�^,2S������*m����˙`�L��U�|i8'=L�\PQ
�:,'�()�if̄�<ѐ%c�$0%i&���Eu��������M��j	��z�"A��vI�EI��o��iX���X��y���ߒ�RV��"�璻�l�/��3u�P&�9_9�ִxDDPiL�����׹%��O�^�:�X$4� ^�)���t��@	�
�@H��ʒCm�$ tY�K�%ϑ�7V��(�ߌVsz�S>�Dq�����xT�ӣ�G��=�;�<�'�GV8��z��
26��	���[9�ߨ��d��@��,�X��	�6
�q��]TJid��e�T�L��X{貔!+A�P�E��3�WQ�؊B/�KI���#=&Oqh)�i�k+���삥;0�.P�σ$��pg�|�`k�,�Җwi(_8`s��&x%[�������
�L�Qi����L�X��Ēpg�W��pWN��-6�@j)��x�a� ~[O�<�I)*�r38�?+��&7���+���W5
j)Dl%#��ua9C�cB%�B0�*!x0����R���:Öu�c�T~�n�%i��v�4��\KI2�EuCD���$͒����L�-UAa
�3��Q��I�Ņ�(J�L4���+2M��|�`���L��a ;-�f�b��Nf��� �Q��"s�w���LCF�Ut��9d%(���n��!���;$�4�a�
��4dvJ2U�"�ZĽ�"! �U�X�)�� �lNi���A��	�= %���=!�6���Yb�j/\��dm;xI�&+\�� 	��!3e��"�(Y�{��/=g��Rz�"�u�(:/�l�В�}����c�K.+qm�F`t���������$#�� F���4d��n��AB��d����H	�4�v�-͆(��4��C=���fi�{��R��+M0���\z��vׂ|t���.[<�4���4p�V)ŕ*6��p1"Cb��Z��|��p�LBT�F�	��F�`�\�����R�^�tUE��`�]��Sr�/����4��ʖ,B��ku�/\�)e[��)�_II��z�s�M	oƬv��q��(YQ	�^V��_�����,�L*_ERHWݙ��U?�\?�߿��� 	J��i�0t��4�K[Q��1�h��LP�2]���=�X*�#���~��9���]�ꒃ��`��ÆA�Ґ $N	�%�3P�c�!pA[-\�c4fCD�����U�����L6��dЛqJop-%�MN�|q�H,iD�@ $ʑB��Ji6��WQ`�Z�`O�2�D^�ZʁL0��W0�⚫+~���'� �4���4� =��7�%��P� �B�F���j�W��̬ C6à-�L�R�Ii�$�ʈ�#e��!�FNIS��S��|�B��!���%N�������7[ғ��&��C@�\�`��<���ms2k�	F.��N��Z��*�4�p *�up-��0bY�L@�Ea�B�����9�Y�7�qυ��JHN,����������s�/l"	C��&Nʙ[&�`0��e�X,�hs����ן�bܺ3>#�߻����{��gg���?x�s���{U��
� Ak�?dY�d�LJ+��,gq��O ֊B�7) ���T ��K2�� ��3"��0���6����_k1~��ζ����`W����힬���~�ᗟ���>���7��_��Ν�vV'_~�i�k���]o?;��j뫳׌�.��Q�ݮ�K�q`�^2�Z+f���9�ZQa�����I��4fJA	��8G�K�0��� F��x�,s9��#����%�˷;+��/���'J��}�w��`��Q�F>X���,x��PV!w��f�jw������?{��߻������+۬�k<�w
�s�����n��Q���r�rQl��o.	�o_��8͑���w^xe?�8ۜ�o����OϾz����͓C��sJ����|�s��$*@zfe�z`�RFb�l�7���̑�?���������	�Y����њ�JL\m�/?�q�d*�!rW;a��q�|�����:6ԅ���c��ç_���ܺ�ҍ���]�֕��ӽ��Pl��'Z-���Y�{5�~ <a��c�oi��.o����{����~Vy�s�sp���y�����t��çw^�\m9U��F<��E9�O�<��ypQ;��y6ՄG�9�0�c4��]�	8��4.�"��Y�D|��7i<���xh0�O[\�1�2hR�d��`hX	�fg�&��&9f��ۘ=	�j��G m�t`ȓ�͌B�H݉�,@Yh� C�r��GNS��`�d �eT%�}^k�	6�df6ۂ�$G%�cȥ$��4h8�h�|�c��Fm+{�
l�SB`ށp�1x&x$�L���"�M���sX���ݻ׿��O11�G,?t 3�_��#���ǹȑfeBܝa���&K�S*���B��Y>\[�T�q) QDD.h�Zz�U�Y���Gh���^�����Ԑ! 4@˿��  ��b(0��z]��@��ѫ�;X��FlrC�_+��X���*IE�g��ؒZ,�b��ƥ>x3&+c2J��b��f
,"�����[���E7 �X��AH#��1Z�A���'(�&l�L������	9b��4���'$�>wK �܍ ������%�����%�%OS�Ҁ,�ֲ����Fg �1�s���� P�-��X� 4���Qq)�!��l��<,_$�z���	���J	�3 ��[\s	3q�R B`�h㩁��zE f�4�KI&LB��dIOc�P�3���I���M��Bn �R�NAg�TB�`E�K�u��B�ep!� �/��l����*1sw 36H��0�h�L��bV��U�!���^X��^��DI�f<�e3r��lՙJ�,V��������`Lܫ�}� ��`F��a 3��?�x9�O��N�.@�Q0� fqi̔����j�O.�t�RWq�H	ӻi��L�#s��!bY�VZVr Bq�_����[��C��� �R5�e�7�����6Z&32@�͐j7 ��\'��1W`$^��8�98f�D�4�v-~����Iz�\ ��4fʹ}�g0���ikN	㌧G��?2���/�R�/$��}��lWfxHV.�4�8!Qa�]f�����hy�˶!�r<�Ί��V8��S��U���^���$f.�(O��l�"(~0$�$:/V2�4�L�Q��-;4bɇ�<�©L�A)m_���N�����O��F�@<�J��S#7Y��;%wH&g���Q�Pu�2ǣ�"2�_���&K̑�#i�	B�E��נ�)��(������hX�2��ŝL� �4��HC #�H���3Ε��� `��"��2 �K/O �A����P�[�)����'$��U�'~ ������F�g���o��J@��>���a�$�T�:�>6xJ�J�*d��Z�d`zo��E��"�S�9���&����f̬�\�r�HC83���Y�\�1(ie�G����FoiH@-N/�R%H^��/"/��M�^CiRJ��3�MJb��;0���o�DD�� 

l��d�O�Qt�i�>K�;���p�Rr=���3GmǠoFE��Ǡ�`���'���|F�dHձWn��_�{�S�a��d.���<��*R���l�L��L�����;N�[�v��0v���9��@j� ���yc�.�A��s6��%�G �s��2*_>t��|ܽ�꭮T�y�lz+w��D���!���.�1�PD���"��"�q*�/2�X�B
�~���2��f���Q���MV����K ��m�����/�5��|��H�̗U,Amz]er*�	�f�	�Dc	�p��
�N��?!b�3rJV�Ɩ�J0�$U��(u��,=��
df�p3=�Kr�fq�9BV�Lh��!�%p	k�L���"���%���Jf2�	o&ӓ$��ؒ&���B��@�	�B�`�a�ʝ&pQ������33��.��42��Ì5��×>Z.a�|�X _&3E.�� �B�r�v.͑� �%f.B ��J	��Rtx�l+�4�04s�&�(����Ҙ��)���B�����_�2�(VA��)7�$�dJ[SD!�KI3r�L`�:0���r`5��b5,���LN���Z�U��on�غ������>��������x�QÈ���;>vj�T�/��Ӻ4��P�.[�4�LO#�)��*J	F� C`2�J�s�fV�ҧ$�h��Sz�u�>_
]��u{�^������w�n���~���1����W��{�Ʈok��s��	�ܹ�>=Z]��Q?gc�`���mD[O&p�!��T� �T��Lf!4�4�N��it�h9R 	�d� S��|xQz�R��d�1��K������+5�ތ��VO?���~�#QA��1^W�`�e�%�'M��Ejp�%�#���9Þ��(�
ݻ�.֯���˯�Ώ��׾�w��^z����}[�Cw����^^�j��Ε���a�^ه�ø��|���&ruc}r�Yo�l=9<���'O���ڭ���xE��*JX������Z�,M����U#���.��'G������N�)�=�ZJ��R�X)�!C�,�`�G�%Mz�A�-��	ɼkE�4�_A�+�~9���]٦�qͮ|s��'WW�W�{gO��yr��͗�`0v��������w9�w3�Y�]�O���Ǣ���gٽˋ���V��x��/
\�W�;W;�G�P}�u�����������No�����r�㚴�[��Ox>���H��g��Vꉦ�������Z7��������x'Y��ȔHȹ�뛇Hz�t����)	z��G�4�2[@FH�#X�����/[3@&3�e��x&�t�S�I6���%%<���;��Ei�EO�RV9�f.������i"�bŐ`��9��]��� 6���X�PFE�I�v$r0��k�B�V������~���$��S��V�'���b�!�pdi8�R�&��$ _�G����p����wD+PJ�fx�E͵���A���$2�`���)_!�5� (�%No��vi��0_9#���#��*J�K�����	�H���;C�<%���x���W�BK�	�昁ap���h0^� E|���U��#�	f`�	"j���رa��)���f�G�ǝ�m�� P�t\ix�yH�)������AhG��?��^2>���I��FDC�"�����W�\Z"4r�!�Ә��k*��Xc'��ɥ�=��ib��Z��Y�`!��,�����~�rt�[�d�!
��ajI��d�˜P&0E�^K�J�X`������@f�$����Y-�����ͬ9X�	�ʡ����cHiɝ&@K2� �8ؐd��ܸ �M�E�Dfx��̽݁g-DU�*`#NBzW�V��Ge�� jx&���2��S��cs}��m\�`��L.L3�ˊ�[��Y2iW�dlș̅n�4z �FIb���(x��[�$rKV3�nD�]�%&L8J!°r�\t��2{.��X��6��a��W�ң���ޠt듒Tg3)k/�e�
��$^�QV@zJC�s�	C�A203DV��H��S9�Vz����    IDAT�*��~��PS���S�4U���/�������TK�cHX�,�A`2���,��Z0�0�z�	)�"p�+�R�,���
&D��f��"����;`���֢�9b��k��HƱ�<͖��0��Q��褊G,�^��e�B�KPK`l>/��"s�ff�-)yqG����F&h� ��K���@M#�p��X^&�������4LF{G)��ɱkGzFih�$ad���#�o�)�y�%"���G2��,�>����O#0'A���F��.*2Ks�����n ����<α���d�RJ� fg%l�R��0��c���G>zn�C������P�橌��̓�G\�KC��y��D�|�'g L��ť᫴rS,_ 3�%�ِ060��ujĠ^��`��e��D���T#/$4x�H2� ����Bh���2<^j�f��U�� ��T zJQl��h�6�rqY����8
�4�*dh�z������8��3ဣ%H�bi��D�h�.��:EH�,���"x21c��-��˄�'�9���X�4J��O)46��i�u�MV%_�����$���˲��\�0�҆w��FeO�x
��4f�v��-U�����ؘ�pW>�Y��VT�}X�l����*7V�c�az�Bk*�0[b+
L�!�d��դ�h 5�{K��\����*z�/B�dh��Qbf�P��҈"m���iX�?X���b��:HvJ��!+�FI��2�R8jrS56��;��U-�5"Q+A���8Q��i��=��k����;���R&����ܛPoH�|Ɖ�I�`N��G"B��5P-�d��pQ8����Z& *2�Fb*E��&1JI� `�%O�˅�l��S�@�"R �`d^�	�`2\ �f�/$��Y���L��F�j�i%�0�	�X���ޠ�*3�Y-`\ȥ�'�Mȋ�<�E�)��!�hu8|�f$��*���ҕ��җ	_�@d�H��Z�e�X2+��k!�`��Š��)�h)2�|�Ҁ��J8�Y!Y�`���C����V�����EG%��ђ@	Yt��{�y����-6V�_sE��}�8�p`q3���D�4"$�� �UZ�%i����L_�2'���L�F��c�O�%?�����q��������}������;/�Y����闧���g�=�8=�ں���)� h|/qw��,�"B�VbUZ�`�R�)Y��`�l)<!=w2�9��E!:�0%k�I�9G��́��o�&Z���q��^Ҏ�j�M�#�����������'���g;������|�lu���O�.�v/������f�x����l�C4���+��$1Ks	��JY����ꥩ	��� s�̋� f2@'9| s�����U�4\�F�1p�[A�w+���s�{���~Gô�׋�W�~�����^�Ьsc��, &��ȼJ��bя��%������ju㍷~𽻫��3�||Ny�W�����c�_�����
���%�?���N���k#�=���Wz�����x�G�����/o��>�۷���uj����TH{FF88���#�r�P1�Q *-"�T!�\F��N��#��i�%�{<ޜh��� �S 乔���%��.H���6<���K�v���u���Dһ:����%^�����o�=��{��}����{{����W��_�'�;߻���yo{��=7���FQ�=wQ��\�z���'�N��J���}ߨ}rj��w_�꣗��<;��cib�ў�ځ��lGag4M���3ɳ���R�Hf9��ӟ<�y��ޠLo���70}#�`���P<\�Ҟ��=o��W�Bb#<�q�`��B�^x�C�dt� e>A�H :���Ĳ(	-˰���X��֬-��瘩�e���lИ�H�F��WW�$�e�B�3��Y��H�~�$@���O�d�d�2 �.��p`�h	��>��aG,u FD0$fJBo9�ȁF	�rH)��}N?�c��fQ�f]n���8:<�G�{��"G��$��l{j��7	x<�;�|!s�XK`�X��%��F��_�ɼd/�1;��n��c�6��(�U����X�
�0(��^��S�|̂r��Z��^Ȭ9 ��� ���@����#�CH1�
!%H^h��X�}Զ(��j��U��$	�G8����W���JV�W���1K^�8�Z�œY  �"V���F25�R�?Z�����]F�����E$SrL�`�.&0���X4J`�nٰ���9*�h|iXͲEBii$��F��A�he 9��F`Z��g�Dñ�K�2��Ƅ�Zr���Ĳ��+6JHz=r�,��a	��̥$-X�R���F!�I�X�u�܉�L�@��RhlFB&�A�3k-��d<Um��Jϒ �rF�n`@��O�4xY �j1������L0����k��q�ɼ�04\�S)#Ѻ�����8ZsBH��C#_��Wh0$�S�i�N-%C�~��V������
G`
�&rB����� 3%2w� ۩6=�A?]��"D���F/�=3w$���d��$Ш�;kzi''`0Ī䊊0�
$�|ĭ����-�c}	2��2)
=�H�����L��e���7 �A	�BA�o�A�4ӫ46�&����p��G�a2脀1��l6𘣕	])�
�a���	��	]���ļ�w��D8fsHz<�{Ͳ�g�\$3�w�����+$�����P��
��I�@�?N<�4�䐘)-=h񒿥��� 3<S^�d��~"W�%��L�
x��L|�������!+J3*�A	\�hJ�Uϵ"f0&�!H^FzxŖ|������<0��X ��6eс�d"�FK��iʹ�fr�'A�'H��%6�C�f� ��%+eiXb���z�;�/Obr��h!��b^_�	6�W z#���������$���gU, �3��ِk��Rj	��ڌߠ����Ç`�v	��|:�\$ m.�9��8�..xod(1oE}x@@[�W7G ��rF�PP�x;��Ŷ���$�	'�X=���X� èH�$)4�!�g�v�	��Q/D����	-S�@I�.�ޒ��+ςr��%3�ൂPo9
�>^!"b�1B�Q���u�B�p�\�� guxD�j��o!ɼ�6<�eM��ܸ��U N��:��J  ..*��\b�y��L�`�[����!oG 8�B�aF���;xdgX8�1KIxl��$O<1�"ʁ�7(�}NV���U�MQ�� �d8��F,o		2��(�q��S7	�K���tǀ��35Y�#�U �a��K���M���M�!5��PNM	B�b�HI��
�*1��P�%�7�`Z*[����E�8���lf�:� e"4�X	��S@ !�jQ�r�@�C���		p�\��{��)DVL��|�MK��_J0�V���w��S N<�9:`�L4]�������X����LXQ�`��:Sn��}��D�(�z	�������d��[L-h�`q��O��l�#�?M�YKr�P�i�� ��q��k��"&�S��H ⧧ &��%�	4F�-�x"Gbihfͱ�>��� ��ɬ��LF�`2�Q&R�Ҡ�]Δ��8�i�x�1p0���d�J���Ʉ��,C�.��г���$E� ����U�h8)�F����T�/V�>L$b%�d$����l	� �Tn4��J���N���\��X�y��;%���d7���x���7^b�����;�½��#���������?~������=� ��5:��G>#��:I�3q���bQ� 0�z�R��6LHm������b G�
����/��l�v�:�\38p���K���e��w������;�έ7^}�b�`��ŭ�����}6��9���e�0㔍�j�T���]2S�Ly�'��d��i=�nKJV��M�Ʀ"B�X����9L�4�ֱ�h��WF��^G(��޿�k������7����3����GH��w�5{��%!s��r,��0˸
��R1�Ǡe`f�
���h�L����[;O�^���fg�����}�p��ݕ�F?�G�Y����	��A<���S��y��ӯ������Ӄ�;��u�����~����;���3���ee�HɐBzs'�L�3K��n�Qq�ב���S��gx�V�z����n�9z�b-��gy,c�	=�|yY���g�`�	f�X-V3L�ȍ��e�-��]64�&����������l����ٷG_}yxk��ݗn�݈֛��վ[��N��&�0ܵ�j��c�Lz-��/l���vxuu���_l����+?z��ߞ~t���۟��}j��3n=�����Kz|�܇��3�fE)s���iV������#���	���\ 0�GJ� ��\g��Xj���3E�皱�B��/�~�䞺�A�g����Ui����y�q ��X���rHo�*
�Yf�\ ��'�4�.�40������Iz�0ѓm�bhx�k�B�1�2�͖�@I 64�� P��򝙔' eY�?��I���x�{n��E���"l_������zp��L��p@� A3���{��Ͽ;��dp#�ʕ+s�s��T��j>Gb��D�!7E���;C����1k![�5�bN�t����ٳg���o]�L"�9����6�$�מf�+QW��Yם<�ӒƜB�6(�8����(�+���1O����q��єV�&9�)��<c��+�H���,�25��rIA�L�M3j����ҳQ-+��t�tb��ąp���F-I��[��f��lķ����F�"غD�@��a�)�e]�F"�gVg-��k���>spe)A�rK�.�D����e���.
W�z��Έ��[��*���,
�~�\ ���G�0��Z#>��" �C�G�����ܸ��g�§h�Bt�HMS���B�FM∪S�)жp�0`�,��h��e��ԧP��ƚ�iD�X�h�p�Bh���x�
�f�Qn�BS"5�R66��u�Vi�ג�f)�&�1V�!�
�cK�ja*�,"K�%@X�h�%B�1Ӕ"���(��]:�qJ�K� ������5�'���b���ۈԤ��ď�7:��o�p4���߸����|!�DK��G�\#��[�w/1�� �A��R6�hd��-�P�8�dy����QJluht�z�$.g��>L�?���&1Y��sZ���ϩ�qLzK@S^{)��0��z�*:z<"�n�4)N���O��8�&>�)MӲp�)���]�=C��B�-�s���v�HˌV������D#�ҍ1CD� ��H����RW҅�#����oY�Լ�I����>f�EiԘ,Q)B-p�@/���1��9&�"å˂1	[�4�_��r-V�t��\q����wU����
�N��gdqZW
�{D4j�E�(rH8]'p�=�fi��R���D���ґ��J�4?�Ğ�#��(%_.D�D4�, �z� ��.x���Y��1�W��ID���aj�ŕ��t�|NU0��J��� W�p��tj�i���+j��H4: �뇔(rp(�L.�ԨD#3 s�F�AfD�e���U]�|�!�R�����Q�Ѳ��!�t���&�n�D�+$�!n���Ԓ��8�gdj�8�rd4�5��'V�T˽oI���1*'�{+��fc�ʖ�Z�z�wѫ(�+�!;:�ĘbR�щ�Z�
���lHK�\?�8@�:��jA���U��3�C6M
�m��(&d�����q���e�,J�(5�tR�8_������,��Y�%X��R,�=��n]�W��*:��ġߢH�5��E_�Ҷ���AiYF�z3�3�V�
Ս�\���>���Yon�u�{㙬�e�h�tk᤼�L�M�d�4Q�IԆ(D�>�r��%]��F玸YV�_��eK�(]�t)}2��E��<�@8)8}�:�\Ռ%`j��������>��S�k�ѴF4�n[Ҕ�	T����sՓ���VN�]�-�΅�B�>O��±En��/w	�b{1}@\!�A�Z���:v��T�|�탞=�L{�%u1S��A��s��
)a�j��0�%#s�0!m��#(Q�G����R����XcB@:z���gd�І�(�)�a��"��I*�v�T:�T]Ѥ�d��Xu�h�"�v�DRz(�hj�[��Ƥ���0&�A���Hv���5/��B�B��I�a���7��8�c�Bh��w��f]|eL#�C`
�8U�!����:��*�h"e	��+��B2�̔c$�б0�R��:�(�%�hF>2�B���<p��,'Z���XW�ƌr�z�г	�|��B�m��Q�H�^`���:�8fJ0P��2_
�����V�/1y4l_^�;vo������=͞_Kx��ŋ�~�٧_���ޥ�7�v���ku����(�2u]��7�D k���^�K����"w+����o���U�B��>���t�J���N �
��O!��Ӱ�Ic��2�^~up|��O_��/�/�^������|��v��=Ѓk�����=}�I{�j�����ߑ�o+Z�*��6��ԃ��8��PR���`U�Ӟ�%7$���#�N&�D{^�p����q:c����G^�>���ϟ���.��@���y1�*9M�P��Hb
d|/Jr�%�E!ʴ��ze^��h|)|������'{�7��˵S��f��v�9#����9�A��q�����j}�,��[��vg��m���.ܭ���7��^쿾��ׯ�����^=86���jlͯj�+������zX2�5��[n�Ӫј�c�*�'bjSb*��TH'�Cص��4�i�9')b��Qd}�<D!�4���u����JW�ϱ��t�������oo����������߼}������գc_��gM��\Jx���.��]��mY*��o�b�.�������K x��9pxsyqx�`�����_�������/�\~�z	Y�؞����Ե	�?��`�}W ޶緙v�F!8�9��������/~�#��J�tQ�Ҵ3��.���� b��N��!䴷�힨�\V��
̨=8"�5���t!w��j��t���7ߨ+sb�up�����1e�����U(�%�=�o���K��CS�h�%��iY@�ȥC8	
�F���m�*78��)4���x�DY:���mW�O�&�7H:����;N�%�)��[��y�g���ϡ�s|�Y�5��Z-�B�o]�K����ޢ�K������LCv�Q�&%j�cY����0�;pt�F��.c���)��VQ���_EG���!q�T�KH%l)\��(E�����XYv^�z���(�#�b�D�+%���JQH�z��tdcK*�h�T� ��s쌷@���*:oc5�ghT��o���唕Z�G=&Ym�8:F��a�C��6=S�[~H倜|��ݰ�O�pYM�Ah��1�V���!�k5�4��&��ߵ�Ê����+$�K$ej��I�sp*Q?���ώ����!;����z VAT�B��T1ő5ˉo��hiV�T{1�?B�� T��ZH�ч�
N��"b��ҍ,f=�!h���[��t�(#�b���7�U.��M9�!��~K�"�s4��~JoQh8���G'8��ɟUGF�7B�"��������XM&%+K�A���'��c�����-���9��>�c��LSQ#_���p����#;��1���?~m4���>��r*��:N�e���L�(�S��D�P
�����%B�E bB���1��VR�i�|U"Ǆp�ٔ��Fxmp�S�dl;G>��[|��HaB��6J1���}�4<��/����4�%A��M{��G|�+�4R[���(�+�zE��:L�茕+�&K?	ڮ:lāO)�^"��JcR�&�[g��~�8.����YR^٩��_�ψ�v�9Klc���Y�.���� �);4�%��Z{d�h��8H�D�v��h���iJV�2p�fueI!�"�U�I��    IDATЄ�hI���+A�MK�2�k]6Aj�@ʦ��� w��f�Q�U�(#S��B��W'9��Zd�n�S:�Ml]ɣIoL�������E��*Ǉh��p�������kT4�rF
���(���5ђ�,�}c�rk�\�tdE#c�p�MS}
y���c$�y��r���:�5�Z:X�C���#%���{*�t����F�N\̋z�E�� t���k�֙���u#��-�<��%��U=q��w�J���MHU( -��(�B�N���;m0�bS!���ph�-F�i��}~E�#QcJ�;�J��7)�C�z�R鲼��� ��$Ғu��{r�"P ����PB�Z�X�+'�sx�)(�O�2m�w��Y���Q
��!)�`!@�u����KY��L��;MS��f$��4[)�>Y�G`j9"8
�J��Z��k �p�2=���(�-$B�L�N'�k�Y��D��,$K�;���̱�΀m�D)�E:͚Ԁ���(�N��r��ʕ�(�1�d�Y��b�T�X��z�R��J)|��'�Ho�|��*��Џ�TK�s��:�l/��M:F��Eh�T���tǈ���F�)�C��ӧO����~���>ܶ""EE[�ɗ�Θ�巜��%V�t����=H��c�1#��}���t�,U��-������-B�"颓X:�R.*�U:_	Nju�C��V���~K�+�pX:r�f�E�E�AKE+���6"��:Ձub9����B]���R~u�Nc�C�(�d��j�0"��5V"�N���Ƿx�@�vI����B�T(����<G���T�����h��0����s��w��z���@��9�N���a��s�t|x��Ţ}A�����ۇ'�'���z�����������w~$���˶^뛢�ߡ\_�\w��߹l�����)�Ƙ|����X�Lg�,��P�9F�i"��1�Q�N�I��M��dZ2L�ƍ�֚�x%Yغ����:/_>~��.^���~�W?���Ӌ�������wG�����Ş���zߓ�Ǳ$ʬ�J+�2�uˁ��-$���^&�DuK���3�\������G�ӆxhs��Q.d-�����`�K�>{7���`�y�uڋ�|%�䈵����)�	�_U��L��^�L�)0��}B����k��ܻ�~x��/����R���������~�ٹ�Z��Q�{S���j��R�ʃ����>y��ן�����7�߹��������YF���/JSc��Q��3�A�ϼ��"S�a��BP�tL�)YO[�m���sr���'M�}+���G�Q�����E9MEM]I�:�d���ĉ/�k��W}j4W���
^���v����_8���|���W|����?zsv��ݽ=ٿ�WNm�Z��M�6�G�+���/4�~w�|[�q���N�����������~x������~���`�����ɱ��γ/R�3�A�3˹�����v톛�v����V�ӟ��ŋ�P��v�����	�%Q��=�B���C�u��0�)IDHE�HY-
]Y:4N����(czg�">}20jh���H���W,��uԷW�p#k����k����W�A��)]Ϫ���&�Sx��rkip)U�(!�2~�q�mJG�Dx�d�JI�t��U��P�/״�H�r��qtn���<��%2�M� qƷ�K�ԧGV��NQ���w�.�ģ�π�S�q�4��?��?���v�`�Qk�*w�x��[W��Q�Zbh��QE�ɶ�|ѶE���L[_Ѷ:��mx�PVE��W��)!��m�W�L�ZR��PFk��MAu��,G�Z��:�7�l3S��h�2��a|���>>�(�,��͈Pu�Ī`J1�y�D+E]���Q
�B-9�Y����k�ZqQf'�tTo��g�E'DY����+�,�\~Oh�B��G�(0`Ӥ S�M�h��9���q0�)>'�id�jt�߈o�I���0���ǁ"2A�Mu5#T�j��r��Ocu[z����[qt�P�B49�O���3p�H�|̑��dw�|
���T� �"����t��.c+�(Gz�DL+��q��6!F���MC�I*Y4h��/K��A�n��&Q]�f�U,
����-�Yb&��7��Ua�U�}��i�E	�6����N�����Q�񁬢��rpYBEME�L�ls*�-��p
yF�9� &��1Zo)�+�~��f�WB4�tx�qzNM"����I���ᦪM�
ߟ��O�rY�]f����lMJ�G��%N�u>�9�)�V�ix����[n���Ʊ!!~�������,~��q�B��� R"]�1�i�6m��(T3>/y��4���N�X����_���D�'��V��S�tc/������ĤI�%�	���(�І���K��@�(�fɢȮ8�ۨ�,��څL��1RF��O}Ҭ
~x�[u����T�CQ����S A+�?��!�G��U�4�L>r�|��2Lc�teR�$��gmĜ�8�᜘|����H����Z��O��A�G��i��R�,�J�(1}Mr���dW�z�)Ԫc�WQ��(���������F�l!F�6$��,�1��5�]3G-Y�H
��`Dn����6�9j�qd	Y�s��e�����b��Y
K��Z��������Bּ+��<��~�/N�T���R�����{�gϞUݴͯ4�B�A�*��"8��9�%VȺ�b����h�.�?e`>�z@�S:�B��~��WN!'h�=��ӑ���q�"W�5@����HA��ϯ+��8u����,5�ꪮ)��4j��@G3�Y�S�H��&↙�M
�RY:BȤz������Fg��J�{�P��rsc�zi�p��C�!�K��f����h�bK�EP?ڐ(ѰV�J��T�V�I\���th֞�|S�%A"A�Y�ya6�H�IԪ�Ą�[�����[4S��c�*p�t�-�qJ������.8�V����Z��䓲p8A����U�3qZ5��Z���s�����>����e̲,�)�����@���������"���9V��(Z�Q�*�\�Zd�����#s&J�a�)����i�����~-�@j	�
ĸ������h@9>���ӗ%�V�d1H�:A�[�\
��q�8�[#k-m��ʁK�HD��jMQ��N����0�P9��FRYU蛖�ߴ��ж�8Bh��(7N��bZ��L[��_ۜ��J��Y�PGT���ۤ�2=s"���� ����r�t)�o��F)���6)�>���ԳC�����OKn�W���=�?}pp�d�0{�j�_���:�<���o�Յ=�nq�t5�\S�)���|QV�SZ�S��rL#���f1��V$�<i�
UHԪMYx{+�\n83��>��΁�ػ���U̽˫7�?�_��|����׏?|�;0g�oo/<�{�˚�{�8�K�N:a��a-F��--������)B�ҹ�idiδG%�66)4'	�-��1���5B����	������֌,S�������<}����ÕI�h���u	�������E�|�=��$��FkN+J=kx�A�#H��\!w�����O�n��p�v)z{�˖kg��J�����~���o4�,�G�Z���jx�l�`�?�p?n��{|�_\�yw����?��k:�n�^��*<S�c�i��Lm߶X��K�@A"�o�q;� 5YE�@R,}�">Y��D���q��F��M	g�K&���[uU�2_�U���Jpp�t,�o]� ��O<y���/zn�<�:�y������/��==�w
�o�c�W��'�ٿ���.�o�h��8<}䶥ǅ�����,s��V�g���������_�>x��=י�/����w7��n���ʲ��Ij=M[r۫��m���d�v�eL�@��/ɱ�]�H��6
�M��A3�
RB��(�F�6��~�������sq����v�=���>���s	Ρ �(���i>)끏)�4M!N�q���C����j*�V�!H����_{����8y�8]@spTWMQN=�!������Ǉ��G�"eS 5Q�I�c�#(��@Dc5� u�����X�N~�)�~���s@��ې�kZK�9zn-�l�щ�����>-D]�NTd�Ah9�D��Nu��ǩ,}:1�L��7:�l���Bk]-?e�pd�&�'�)�ɜb$B������ִ}�ƄL) ���S��6ͪk�H��
�떲���f:+�ǀ,��K!edY:q  �&r�A�=�!�)0���PHJz~m�FLj	*��BG9f�8~�����V�n�����B�W���da�-$�lE��pӎ�]�YJ�!h�`��	��F��(�8Z̜d��Cr�3Q���B�3"�Z4ӕ��V�6*�h��LK�[�݅W)�K�����S�8��E+�)��(s�����R���k�?{�g��V��L�&ъ ��c6�TQ!N+��g^Ǵ~�&�F�QڈY!Ӳ��A(A��_��R�u\�IܔfY�.�ĪLu�)A��"�Y#��ȓKߣ`v	�r��v������S3��jJP��ݶ�Rtj�D� r1�U�h����rx�)�L8��*��vk�i�sB��;m��8N�f��)\]>�7VT4ǈ�
�1�P)�9(�B��C�&bZ'J����Xzk�����Z��M�B��LD�,�#��h>rL#�$Hm�)�XK�rMg]���s���B"�=wQh�hu�\!L���:�n�8J�%�{daz��I*Z��LJ�A��E��!m�i:r[Q�f ��(���z��L���:I��:Hcd�L�VÍ��SN�BQ��vGݶ��9A�9X���P��Dx�YSc��Y:G�:�Lj��ϒ�jR�`�(SH|ۢ#��6_�r98��s 8@ǿ��X����0&S��£A\w	Y�� �)_�)̻�>%rp*Jd[ �N`�qz�����9���&BMt:�	DC@cd1!gh��t��]�hO��|>$�t������"�v��F�tt�����h7���@ǘ� ���$rR-�靔�x���iF�[9�X4|�t0!]��KFkWKz�|��s�au|oh4��P6mx�h
�(�'�T���d��K͆��Ҋ��m�1�|6�(Z5��R~�Ç�jK�	K�G��s����[����[ rW������Z5?���J�f_�I�Ƽ9��9�Z��8�0%��w��`*d��O-L���W�R�J%��hSz�i��+T�����F'�n[H�|&��䢩�1u�NϘ�9B@)V�G��4�Z��s����hjs|��XX�=�'k�p����'-�VUQN�n.���Є��p��խ� �0�*F!��ϟc�y�\K���U��iuj�k�J)vF��T����6����&�BP�B�QC#ۧ�!ml��5���!JS�L]��gϞ�x���3���2E���-ڐ�ʵF�8�%�
q��G'�Q4�20_�D~�F=�P.�Q�?B��<%VBE��\�F�)�Bۅ�'5cY-s
M��CG9��)�H{k���Z'R�U�;(�`}�9�/�ȦgUD�Fǫ-rR�ID9�V����%��@j��B��,�a�N_�^��3&Nv��4�i�Ls���I*a��t:�S�h���	�X'ӧܖ�HxYR8v�=�H��*Z�h��	4V����C�z�hCȽ���#��;P���9������������o���s_U��.�Cz롷��~�V������6p�V3rT��^�$$gu�un�_�m7"�eCk�ȱ.c K��o�:3M��F�f�BԬ�	`	�w�<���2�?rsq}��g���|���?����>�;~w���������?���['�~(ו�����TK|��FS��uؓ$&ӭh���&��GЬN��0�#R�,�N�U"�}
�Hg��x!p��E�?���E���2��-p���6^��$��iLN��B�g�i��Z�H�LD��h���Y����^�|������+G���j}K�7n]������I����mn�]���[c���cpq����C��Wח�{����ٻO>���r�����~H�b��U��{S�[��qZ�ڗm��m�*�(���(�4Kf���v��{���{V�n+d��9�}����W#�aջ��Up��عP >}�Գ�t�F���d]gt���1G��׏P=���5��tWr�-RO�~2������������?:~�����恟�u;�z���,�������yx{|q��Ρ����u��Y�۫'��/�:���/��%֋���8��y���]�<y�r�˫��7=}���o
�M�b-vO����r�@f��e�z�:ѥt�J���з3 d��BȦ��KYzGӕ����@7�bV�� adsl�s��h�Ï����~fE�q��v�߉9z�o���ɀ#�ڑTY.�@ǝ�R5YmY�B���@#��_�pthSPE�1[�,;�D�?�U�p�����+']�Q�6Y:5�4&B�h:�P��fv
G�4s(S�մܚ��o~�̀K^��B���p��'?����i��Tu�ˏO>�ȀzC�Q��L�4�Y'����Vֿ�ۿy0�|��ij��㒎��L5F�VcQ�>Dn�h L'�̗πę���[Y��ԊR�aBpN�F]1=�(њɩ8�,U8�N�*�[�����d!���X �,>�O��Z�j�ת�%��R��)*�,B�V�2Uȴ�B���(�����b�hr٬���|Y�1�
9�U��E1	R6��i8f��FV	����U]4���J����K��1|
��Y��P�ALG<~uS(=~8��U�9eA��3&�b{M��'>���wW>�@v��Dj&r��X?���#��[lY|Q�����y:5��G��1�\���BÜD���>����dMG��(�6�������F6�rǥi!u9S=� Y�Q�r���N�h�z�!��0�M����pM��#;)�U~k�Dc�^�A5+U���j����B"c&5�Ma��cM©�����h	�	:Q�Tb��qD�G42ǔ�%d���M����Z��) ���O^u��UQ��2�Ң
A8�E�/nd��|�|�i{�N�Ƥ"N���V-g�V4�tL˭~;S-S��d������E���o�C�i|�)����Q���{�J�*I�Eh�{-���U�4PR�V��~��>S��i����=�:����z3�j|:=eE����$�T�O�i~�	�e���gh�D+�>hU'�ٷB\��o��X�:O�Ӕ%+�S
�ml���!	F��*jH"ݔӔB��C^�[n!%L���4��o���	7�H�6���hʤLV"�C\��G|ns�@�3e�N$�*��8����j�C����)�Q!#�Ȧ9%���T����(�8H�h�P�%�Xk&��l��LJY4tM�:@@֔~�6�&�e�NbD�c*���kLV��%��u�M_Y�����>�(�Ȉ�a�W�d���E3՘�s��0�$�E#��O��B tʒ���I���vRE���;C�*Z�Hy_l	�t�
�U���'�)��k���uᴨ���9��6D�v��.��C�S�R8�u.�>��#�J1YǗf�Ԋ[~!�A�C-A�T��*%�k�@��6���,+�i�M�%���S�t8�A�5B:U�Ȕ�g�H����� �ˡ�����K�(�B;cJ�2Gz�Hg�)J�T:8�"V ���D�w�Ʃ���5��TO���>�qnrM-�M��\jD�K��t�op�)=~�0���cJJ�J�և>R��>(����G4>����pQ1iب��N��~��M]�~�O>�$�
�d�
+*B*_K�����������	�с���#�)]��MKL(���D�4�9�6��w�?|��+dTKV)!S�6�2
1�6A
����B5��RTDpb,ŭs�L������$�iQ��2(fR|V�/�� |�F�:Lh9p`���p�i�qD�D�"@�Qט�/J->F��Shh�)㐒�/1�t����d�l�^�,A�8���A���<R�k,���    IDAT�4%>�:I��Цm�����0�f�L��������Ӽ}�������c����/f^]��������ͫ�~���ߘr��ˢ� �;S{���Ҕ�P+�ZX=��ָe������Y�9@6`"3����~�dp4~��Q��qD��U�My����<�[ p���v��6o��^^�����Wn�>������������
�V���_��.�ү��*T�S�[��FH�,�4�%H�@J�$婘�aFVnLO�	z��3Q#<��h�!�j�.=�;�����f_9��҃]G�������S�����|�kEIS#��r"@&�-
lkTѻ�X�}䷁�^�ߜ�˨����u{�y즦-r�ଳ�u��✸t��}���ݴ%��צۿ{����/�o��?�|����t�Js������ݍ�m��/(����a:w�A�����oOIB�ʞ2�kU�ɲ������xem� �C<�0�x�����8A)�
�g���������s�Ha6H�Wǌz�W�-�׼��lZu�	@x��?|��ã�wg�����˽Ӄ#��������ۯ?�ڿ�����o_=>�8�8x���͞]\��^=\�a/D�׾u�O�:~n6{��[���r����d�����S�._��?�;}���?��~�/^�]��/s��r$H�����B�T��Ta��n�L�B\�"�i{]u��R��P�\>nӜ08�����T��*g�q�A<޺�%U�����g�J���)�"��iu��p�k�#T�8�n9�N<g�Cϯ�N3�U��5��Y�>��S�Ȫ���i�JC8�yyUHI��v)�=�_-Su=ݴ�p'��*����F���Ё{g���A ��5����:D��bZ������r ���@���F�mK"B
�
v̈��Y�~l�r�S%�����nt� �`v,%�]��b�:�p�4���Q�L��R&(M�|"|B
��?��,ܺ�++�1×Hʴ(~N�� ��S4�Ȁ�솑�N`uc�*��[kD����ڞ����g��ֶ�4!;ֶh�&8�8���L9ӘPS��eU�nC�2Ƒŏ�O�u�-�U��k	^W�9���T3R��e�J��9UO�r�R�JA(r;&g���o�)eY�S	�B�kNsLhq��F��D#��� �HTΈc� ��@�h� 7����t��M+g�	j���	A��BU�,]?U��XE�1�2gʥ�LVh�qL�h"E��A.$�0�b�hF�L���)sv�����Q>����!��Gv^u*NQW%F6�NRR@3-��Z�D�h�
������)�a�l�Y��F-��P���Sh�_?���L)��K����8uqب�wi|H���i-�J���mTOb����ǟB���^_n�(Cf9p�#^-����$k[�����h1%�ZVݦ��MHnd�81q ��7��B��_?�V��ճ}���R�-�ZQ��r�S�F�<��J!�W9QY�k�X3�Ɂ����Rґ�%L!��b���P�S�3pX�)�7��I��p��`D���`JIm�]<Pn`L%8�H�1e9�p��Ň Q�ٙ�� 
��n񻓇��W���OJ�)'��%"*$R�d�m�c6��?� ��%�!���"�X:�!�@Y��!�%��I���3r�����I�b��g+j� �v�p���d���ŌP?��r ���§P��8Ԋ�3@�r����F�g�Q��(�BO�rMS(Qn��3�h-%[b:B8F�Ʀ�	Gh	�)k�l灢85	oOF�*��j'�J����m[W��9U,]��� 1SZ��#�!������N��7h�9=����#�\oTB!4��{�dU��,ܻ�BFY�Á�dx��S�N�#S�>�,0�(4jۺ�HA�)fk��dy�U��0~���r8�����6���nѦ]��u�$��B�Ԅ" �LWp� ����9Q��DukM�r��j�	�@r�eQ� ��b9�(�nE�A(s�N����)���� �9)QH�UlE���Ј'"+Ax
�L_:���� G
r� P�dm}zP���}ߚM�J���bsp|.dt>��?�3A�K����x�Bc��/�=(�4&����+��J{}�T]���p�
��4x�P��Ֆ/4��w�Ĭa8CH�Z�>d�C��u0jX�DSNʥh�h��J
����tN|�E�mĦq����De:e����H{h�㷺�F�E�L��õj��I�K��M}
Z?�p:p�|�Aʬ4���a|�S��@h	m#^c5l�M��h��Z��V�ƀ�k	���G��:����!�H�FV:Y�QQ�\��+����Ҵ6��%X�Sz�_	�:�~ ��'.
4&�.<NEk	�L�C�Q>xxy~ᆁ��'��<rc��7�^}��ş_�������J�=t;�7��^�X���^A�U1��:T�C���_�R���!2'�(�(|��{�Lq&��\g�.��gE���lo����������y�;Ҿ�uq��W��߽μ����w����9�͵�X�O�^���@;�koM7��_����uZW�j[W_�F���B�����Kw��19�՛bV�3��2k9�R�K� ������~��g��8�����m��r�w�w?��������B��Ҁ������ƦF
ӮFE�l�щ'���}}��U�o�]�{�]L�Ƕ���t���-�kg̱���髃�}�s�������o������Z�ene�'__�t�_�]���?��>�vks�����r��w���-�h��;��چ���w��IK�0�f-�Ķ��(�#d�$�X�R.n�xf��YWu
y�V���ʦ-��!
%�ɡ�;FpL]Q���0=�ܴ�L�i�]��t\I {Q�vc����7�)Ĺ߷X������<���r}�W���.��߭��ߺ�i�O�o�?솲oX��W^Fƽ�Uj�>Q#��q����c�/��Qm���������ы�������پ���}�k=��}����`�K�m���-֔�7�,���M�`�!k7JIǱ�h���:X1M�W�c�0)丳�Jw������~��B��4�7�4��iF�U[�
P粀_�tk�4
�"�?G<DQ�"ChB:�w�H���([�ε�6b;y��:
�"Y���S���T�B��o��IՑ�%��E_V�ߘ�A@v2��ҙL�&�niVd�	����D%<��,�(�s��QQ#Y48�}��(�sǴ�8�@k�=W(��ji�Jm�UT.�DE[�(�WTi��"jhr5_��#�2A[Q�|R4�t���)����7%�ɏc̩��� $N�12�)�чc�*ה�jLh�)�3���$<�t��-Sb�D8�R)u��A����l�[��m���z�T��M&�N��	�cV�h��ѡ�h:����J�!)��h��=������5�d�t��9!��0�P�C�SH�F6)&Z!~N+2j/j�D#�
����"].�ft��c�H�c��mEv9EKWW��]}H���0]Aj8f:��p$B��SV���"p������ i�r[T	���)k������8�MK7V���\^�@cr�P�&��F�AD�?GV�џĚ1�:���FV��l�������ǯCL����+#B�LW[�����O���Z��g�m�X��IPME!��5A�1!������)j�|+
M���"�՚\�V��1Ef-A"08)����o��N�J�W"���\t�8U���R�Wȗ�Bc��U�L��ar�!�83��o,^�O���f�)��Q��4)8��#�n�8�# �I�,�4�:͢�Rz:���B9����?uiB(8��q�V���I�J_$Z�	�҄�곐1<M�(�h"����#Y�F�RrS\"�tS!��9C�P��K1�3%v��ǡ!q��BR����&��a���S�t�r���I!�2M�BU�3����r�����Z�|��Ӗ6�Gvc��T��X�j'%ٚ1��>r��'\n���M�H�ަ�<v 4[Fb�o�3MѺ
�D��t�9��Ԍ�ǩV�EIy4�6GV�R����s��85 ��gŢ�����RX�p#��i�83�͗¨��,�3�9@H��IQ6�(��t)n�~�� �I��A�
���%�L5�߹�=>�ǔ���&=��J�~-��Ł�V��5��d��\�p����ѩ�\�� }����QL>��g@�:��4�HYb�3Ԍi��A(�����2�8��\ȢFS!|=3U($BK����~�E1�X�T�R�@:zPn��>�KX�q�@;o�j�n�h������ ��Ĭ7�J����!H�DdY	��M��+!7ASx|�u24�TAhH�&(��N�>��F�d��Ć3<{R{FE�>�Ғ�Ol|hF���>�)��􉩮Fl�Hĉ'��ei.��QT��Q)FS����AfLN�V�O%�pU�YBQS�Z"K-Y��9��_�݋ Q�$�B��E@��I2&c��q����C�*e�?��|V���!u�!nD��)�(��[�=!����ȜfMM{r�a�!�
|����J(]Q��7�UԹ�&!��~R�(+�D�Ԥ�)�b�%�l��jOT���2��h|c��M�a�H�S����b��+L�Ԁ,�6Jtj��1�}C�8�>�tJ�0!|֞L���8����p;������ţ���'�?~�_����囯����~t�݃�8�M9�=Uwh��*��"��7�|�����C+�ap�O������7�6)	����)с�J�>BEI�Wt�"ϻr���V���\��}��f��72=l����~s���GG?{�~��������������?]����K�\��Z�!�8�o����
'p�jL�} �SQޓ _9߶-�o�t��iv�<�E����m��8;�,�#�ŋn����tW�g/
���5�`��	�9�u��Bp�d��D�8�5�VALm�l˸�8;?X߿�U�u�	M9_��9�p����rcٶٴ�}rӸN��+���גܪ?���������ڭ��:q�?��2����y��7o��n`���6v��6�^��]��_�M�$� �f�YQ�N�S#��HJ��%���.˞Є`"xU����(UL��
���?�p�����r���ӧO)�����n�uP5f!RШq�-ߑ�A����1팱X�ʐM[����礶�ڵ���o���^�ʫ��B�����z�g����&��^�L���yq����C�{Ӿ4~�ii��99:�=��v믪��R�����'���l}�s������'G�|��q"�����\�5�g˱:k��d�o�o�E��L�̎�)��Rp�4 �&S�{8��G�&Ю��<!k���!U�u�
o4�h�c;�~�B��CЌ*�8|����q�Ы��ފ�p�4ij�FDr�҉`
9+��&q�DӀr�@fX��z��4k������ D6�h	
)*�AX�8����,A�|=�N����+́S�n��c�2��c�Y&��Ϟ=�#� 54m��=&E�����q���'P"ǨP��89���2�[B�S	������*� �d5�#e9Դ�ړ����\�1�=T)Z�5���m*��ӑ�/jjdx�hR����9��I�_��,��Lg[Z%�w8��F�B��i3i���u�n��M�s��-N�X�����
�M�h|���RR(5!�K�������IJ-X�|]A�i���nb�Dv�|�-�ODW%II�[���*4"�[j�-���G�N��\#��v��+B����VuΙ�ZUa�m`��1MS೤Ɖc�4&�8B���#����L���Č��� s�v���R��l$�s���wOY�	�b�����#2�p�L��8nʉ3YME㘪[bGS`|~]M�"L��|#�X��]��(�p@��UTȣ�(�Bp2�c�98f"���j�h��`ҟ�%[�ħ���r�b4e�z��>?fS�|R*2SY�,T��(#�&R�5�SzY�G�2E�܌�dq*��}�3�<��휩�T��T��+NYJϾ�A.r��h��R.eJ�4���l;���j�k�S8���7�r*ߔ�7-w�$�TW�y8=��C"�����G6�@f!��L!�@v���ZͲ��Q!�R*$*%�#��75�^m�Ȳ�:Q1�x|c%�mZ�8�Q{�"������r��(�X�X���5���V�I�BL9�܉�s��o)�զzw8ү�TD��r:S�*�'�3Y4QY9��>�Lq�k�!5P���.q�RtrEe1��ݍ&���I���p�e�J�[����)��10�4r�o%��C��FQύ�\�k���mՅ��dG�(�E�i�C���wI,�����ӊ����ܚ)�H��T��'�2��)�G7��O��󙨔zh	��]���1��d��+�r8��2�XQ����p�1[���@���M�i��,E���5�(��p�#"7\]N8ΐ+�3��B|&ԫ�68��G2�U@�]�Hgq8Ô;'0���t��7u�a�F ��m��V�n#��Z��u�X?��s"�/*K���ű�e	Un!Rp���7E�t��ڤZ�D�|�F�z0�
Ee	��*0;�#$�ܪ��7A�h�=@���B�P:���L�.%����r}ʄ\�d�KPT����OǇc�w Ф�	o��W��a5�Aá�Ϧ�@�B�u�pUJᫎ�aS�T�z�TH.��j�+Wbd>��*�����L�E��Y���u��+�ȳ���*�ѦU�CS!�4U+�,Z�e)mC������ѪC|�E
��<������-�(e���R-
�)PAє[8&���rh� \c��Sb�	M��p�D�*eڳK���OhC0�6����`�c6m��'�DӔG�S�f�΍�	!׀D��mb�q�|�{c���"��LR�����������{]��i������'�ݞ���^�������;W�~eS��}R>��(дVw{�R=z�D!f���A��&�J@�t� �L!
Fj��R�@#�6["�Xێl7��u�@����#)@DW[�~~��$�{��J��_^����߾��/���������������Gx}���_�[���^�v��LD#q���a~!Mb
�c�q��Lcr�[�k'�{-
Ynd#�)>�KI�O�؇�@�e�4#ľ���&�*n���E�3�}І{
�1��8w̓K�j[^��P���)N+�\�\J7N�H��l[�����@�3����w?��o�O�����_�D^��/�Zp�Dv��X�1��7]7�4����*q�L� �����w�g{�P���RTo��c�	YiNǯ�����ը�t� ��֟��'|��J�����R6u�|GӮz��?�L*��閧#8�)\Q�#禩r���-P߬%�AAP�8�"�J/r�����$֛ܲ��Q���]^�x��Z����=8����^]�������o?=���:u��n��ܜ���ݿ����4�=_�\��xw�Էm���u_����|{{����ã'?|���}��O_�x�b�W�D��[bN���jX-c��Ǳ�U;�ہ��qi���
k\o_j���!�:���2��I�a�8LE���YU�PH�)~����(H�;j��ph�����(5gE�9iZ�6�E�L	:�rՕhLV��F`7���'b�'�&�z�h	�B`���C��#e�A	�Q׈FӮ���1~N����������N�[}J��EЉ��@%GJg���z���8�*
Y�bꮧG_�]�(�y����+uȄ�=������,�Z����1���Ѻt�"Hw�B�=�X�q6�k�q(S�ND� _.p^G�cE��>���#��4�����b��	��hi���1��7�fR��) i���?�Vͬ��#D��[cp�JǦ�����O�i|d��	�lg��i����ѿ��6HIg|�ܩ[c
�Gt���	2Q����df'O8    IDAT��Ms�)!D��DjFf:����
8����9�s��DT��ș�) Y`�+�R*��BB&�T�Io䈒25�\�׏X��m�S�=���w8�s��J�="8h1Ц�)�1�$X!Q8����J�Ȫ�*��*Y��(jd��e5�9[|9�Ʃ��M���4�f��{��C����r�pF����XQS!u[u!�P#<fj@HG`�*rX+��\dN���YR���}�#��l�lT�Б�#R9�p��L�R��UK� �B�8� T� �χD��a���D�(
�bZW�R8B�b҇ӑؙP-!1���:�"kH�p U��oipQ>��5&}w7���cP����1���o*j��Yo8���<�]d��2������Ʀ��mYF��g�i�Z�i�M'�Dt�c�z�>=�I���s���y ǋ�x���۟*q ������M�:��)����D�Ï6=#P����~VԘ��r�wu
E���X')��JܝB&4�
\MlFV��OY|��a����T�X���Պ�0`�������ʹZBE)��B%���["ʤ�9������g��P:��Y+�i	�t�B!3rhbvB�T��X�U4����(��yp𘦝|#�����bY�0��m�����D�2C��	1\�-�cD(:�" 5�d��8�VB�[j�p���-�&�+�U�ogL�gw�W�Z%�L�eL\��?���Ƕ���xݫ��6v�-�F(	<��~K��y�H��C�4�b0>6�Ʒ�s�k��V��!1�7~�7Ɯs�]��ޅ���H�n���Y��8B��J�9d|��)7���D��S�j�X��;j���[ĘS�~��	�-L<)"e)ԯ�]��1#��	G�h�H�f*�\�%�H�jf��<��>ͨ����'�c���W	���A�`�L��ɑ(˔��ԌC������u=sDqv7�4q��U�_V��s�&Mi�pL�WN�Vk����ԉ��� j���?�9�Z��Vo"y���ҍ�e1�!�FA
�Ě�_	#&�~�Fζ��AT�,�Χ[j��6� 1u��ܘp�!��:�zn�Ec|c|����X�Z���RВ2�(Zn��#��T�§�S���9B�cKiJ�Țr���]�w��!��`%�WΨOk�����XѲ"�i+L�!e����! �p0�u^���Z/G@L�YH%��!�!N6RBD嶖�(|NAԴ��B-6�4Mk	!Ks�8��3��p�N"�0��P���_�>ʵ!EnjW�,Ưs!;0� e���;8\^g�g'�����������_|���K�	촏D���*Norj�vi��ݽV�^%ԭ7��"���4��e/���]�޿z���]��B#��	��=b��(��j���$�'�&B�F0e��x��X��<����ť/5u�\�������W�>x���>԰��ݿ�?����g�_�?~j[ס�p����5@YK
5v��kZԈ �f+����hIIOj@��#q��0R`�����]���%*�_	�������M�[�v�=y���ބ���3��\��gINUTE�nj%u�b*V�B�VZX=�^��m&D����Q�%'�k�?����E_D{��g�R�M���^�\��.%�T�.{�L')������g����{��/���'�O�}�}�p[vKXU��Z�m�3�;��f�쑭�ݦ��w}Y������g.}����w6V-���d��Y*!�g3��7� 噇�0?���zSKo>�)� 5�8EOR���Fuqt�r�t�]
|)U�&5�h��-B�X�����}��_�ܻ�7P_<y��/?����ó�Gg�k^�쭯�][�9t�k�v��u-�(�{Խ��d;��[k���.�^�_�<x�������8���<�t���M��=S]�\ÞHў�t����N3�Q)F>����hz�8<of.H��\N�]�|�y�ϒ����՞7�댲Dղ��kz�E��t#e;�=4&�hc������#���d�*�c0�RnQ�e)��tʢ��p��t���G��E����h�ja��96�4P�Qu2���������%��QЀt&�O���٩�s� $A����85� ��t�w Ԑq������Bj�a9zhE�h��7u�L���k�X��u��#3n����Y���>5cH�*����	r\r�vX���[�(2�4\{���S�FK�2㘦����n����L)U��M����Si!��4��Q�M���oD��>6��J�� -��D�dM����)9�C�]��R��($���Yz
!@����S�U8�c"�(!�,K�7M�_�!~�<~{K\�h������S&��PH��3R�Q��<�S���Ȫs����Ufk>?2���Ȓ�(��B�9�!�bJ��)���.��cN�V���)�Q�a�g��m��2�M����ء,�fD�8��@S��@өN�)1�����%�b��t��@Ф�G )VWhѲ���NYBEe	ME%����(T3ȢB5-1�i����7M�4��2[x}M�8F���+3�Q�G0)�Bt��+m�Y��r3H�%V=�Tz
��6Z8���䷍h#DM�Xj����6�8"i�1�
�XV|�9l�M��s�Y!>GTEG&�����͘��"�hk���WV˟�JG�+�_9c�8�3��2�����p)f:!+���#j�됝r�BR��5�z�'5�u�	d|R������T��KC��B�SVfY��Y`�S�N�q16�^H|NNsd4Sލ� �9�F�f�c煮�A�lcUd��G|v^�ju��'U1����o�t:%B8?<�K债�)�)K:�����"�3���1���'1�Ҫ�B3���I/�O'Z=c
UnwѲ�	�"|�J��Z*d��vM	�P
I�gw�(@�-��$Bp�b"��G��jLĨ"P��tN�ɶ�ґ�X���F�>�\M�����n�U"&�P)���|Qc����ۢB�D��d!L9�&� Pѩk*:�.�Q�H�t���p �FY�:i
�J�����>��p ���8����K4B����)�CcQ8+��8BSN�|�|��6�ÀLV'.�\n�h�"#L	�0�	�`�ɀ
�'%d*ٴ��(Ģŗ�o�Z��p
�;���-�4
�L�S8�q򷲋iZb>���?�)į���d�[��(�0�5�ŪR�mK�J+�էP%�2�cD�O"g~S�cH{h@�Ȧ��+�(_�S���͔����Z���Q��)�^J�\o�2��N:��I���X	�hq�/m*�	�N�����p�S�%���&���25g�7E�H*'�x3G-"��D�(K��XKh�g�7��DfJ0�h)F`k�O�T
r�5��ԏ1�|S"RL�D�d{#��F��W�ͬW:W����M�e��M���B��s,
���rYK�p2L)BF���h8�@���P��|��"[�D�����ުH)��\Q��t�rM�� :\��AJG:&D��i~���H�Jӻ�)m�G&������O	����g�O��?����Ǟ:m_@���q}���W�{����~�d��6:]�*����T��� ~�B ��N>�m��g+B�ȱ�D���`���[�Q�ћҦ�C=MEg��T�U�#�ҌrQ�m�Ф��1��)���+}��#ߛ��OϞ=������߾���q�K1�}�����c�ڋ����%q�k5��ٮU��r ��������Ň7�]��9}�M�sRsv4+�p�����Ecr�z/]�k@T�9}_)P	����Ӂ>͵��391���`�{h�W�;�4ꎹ&ڂ
�$WD�u/� �F&�<(z���'`�ᕿ�y����J<�\�=�_����X��GiG(�YO[�ͤC��ѫ�˯�~z~}trvo���§��|D���-����O԰G;�Si�պ�٪m��
�����=�KwQ��֮)��\4)=_�
�J�L�� (�w��8*���8A�_��NS�G��:/
:��Z�I��0�S��B��5�"b9��܁�O�������}vs�6|�K_<��SW����_<{�������Gg�$���?�/�� ���b=����П?]�z�y�{i/=!u� �ka߿T�N��wz���?�n�!O����g��W���Wm�I;fժ�ڥN��ApB�'��BsV=����x.�%��c;�����35}��7�*�m)��e�;��Y:�D[W�2�t%�L�
��VE���i2�����f�U!F4�!�G�=1��h*M
.�!CD%�_	Lו(§O���E�1R�(ʯs։��'.Q��L�Rd��4Iq$�rۢ�P���:���L7Y�8`�!o����U�B������y������M7q�;��]B�;E�������{�?}���n����T�oD�hXQ�+�_��w�z���zm�,8S��͔7M�*|x����J�tQ`&K?�!z�bDh���N�)�0S#2AMcJ��R�r�8]B&D�(1K�e
�����+�-c�r�96Y!
h-G"S���q����6�������'F ���R�j`�)eu�!��(H�E8�L�i�����L�X��)�O�h)�̈��r��qX�Ff��f+R?��b߽�Ky)�0��T�OӢ�.�-���+�c��1�H,�2�EŬ��ж���G3���Ip��!M���2UA�Eޢ�B��Mk`�S2��0��('BBS�4��� ]W85��饦6�8�72SL#�!���~R6��B�'b�8dN���k@z�DD#�*�#��5VK�t8G!)iN� �������̩�v/�����dK� ̶�)��/��[�hu�| 2gv� G@��D�.�@�Ȅ�%Y�l��l�e�)��5ںA����XJN[�_�Z�賥��}(K��#2����%R�B|ڨP�F>�-�n�*���ힱR��Fn�0��r�>�JSˉ�o��7S�����g�J�!r�i�5ܸK�%�T�)͏��~��MKe?�)�Toov�:o���4ߒ�'�#�8��ā	�\�1��������t�h��+7`�R��dÁ�N֒G��h#����d��P�%Z"@�2�� �q��Ţ��ԃ���g]��l�G0�g� �Q��"���X�3�D F�`E�3Ȉ ��Ʃ޴�Nj�b&8�	�B���O3�p����Dd��n-������p�,~?%����VdE9)w�zyG��PRjF?4"��H� 	��R8@�� �\��X��<6$N:��8�t���f8B�)'��i�I�@(��n�UT��i !8K�2酀��X��u��������j�Jg%:8�]M݊V+2f6:�BM7��,� D�N����G�B�(WN4?�	9F"��'.DGJ��5 W�DY���i�	�?� q �ژ�8tB��8>G�I� p�V��������35�� 4��)�oP8dS�����U ��Z�	
��+�,%_��)�VsXEEk�AȬ�	��i�"�E��*rsZ��l��B�IY-��tF-�g��5��ˁǁ��| B��SV�F��_W��5KS��ZS�~��U�B��G�W��р�<�J[&g:����#į\�'��W��Z���rE5���Vb�-GJ4#��Q� ����ɒ�1��c4ݕ�4Mq��rA#��>��6�6���W� �p0�,S6� |�|Ζ���nd�l�i�W�o98�"�L��t�c	���hF&ď\iUF�S�V���CZ��Z>��J_���Fג��Ԥ\G�CM]_ݸ�=8�wv����^?}����>��}������c����z�=��g�z|%TJ��IG���f���o�ֿf4i��==����sr-�hi��@����t���u� <ۭ��2q�6dye�h�!�!L�)j9���F�i�������&�U��g'���������~�{���kG�'g/�y(��������o}>^�6�_	<���IS��m?!���ABMu��w�D�,G �kl�qځ�[�u�w�еg�^Z���O�eJ
.ڽI\��2�~;ǳ ����iz+����*�q�����|�SET�ul�0�ч#Wh��zZ-8ߔ3�K �W�jW!vpxy���셏������˳��J��}\/[����a�NS?8./��V���;�5}G�p�g��=������/��/VK�C0�jI�@mm%�V��:4�j���8./��d��h�r�?���{j����j?=F���B�DL%*�RT-7�n�������**��i��(���?��OT��Ж�y	>�)�%�8M�:���j՘{X:�3��y�Z����M������>�w|vx�����������x����?N��V����tc��r�z�o�N�x>d��l����ޕ��)��s�{ǧ>;�:���ٳ�������n:�ti޽^�7mS�
�����Z�P)�q9Q����?��]��S�t*��bk���%�9z'�\�}BV�A��ش,|4d׃G�jI�C��X��3��D뇯�(����9��mS�h�-"E!�=Dns���`4��,1��)�P��@Lρ�\o�V*KS"FL~:z�3�����)�IĈ&!G
>#��+�;�m�I���TQ)B���s�B���Y{��<sЖ���^�J�WTc�������~�m'�Ң���z���$N�}j,Ko����p!��/q֢�z�o!�lo!.!k�ɤ���u�ҊΪ9ȍ*JI�,H|
JU7�e�o������)g��z�bm�è�s_R�~��r]A�ܑj]m�(��
���e1u����#�3x�kFuW�N(K�}�g�*D�` �#%�G3�j�+�(֕tN�)�Al��ЄTW{>�6:`|#��S�D!���k�	��S~r d�����d�Ms09�OS#q!��e�՚����&2VB�!�02�]���Ԁ�]BwR9hB֎����X���e!����h��6��i{�H���T�8�m�F�:��r�p)I%K�k��Z�r"'hZ��z(%D�&��D"��Z�B5V�i��Tj�JMPz:�)'�T��%�A�T��He�BM�9Y)�#jJ�V9�$V�Ȇ���T7�oo�#@���Jg�?Gn�RL� l��2۫J�+j-���JpHu]qX����.?A����qh�/��8�Bd�S��(#�U���yRf��\j	6�%X�!�*�� �O3�zXiۥޥ��)d�S���h�������A�&:p��V��ЀJ0�Q��!�I��6��M+׈��,j&�cd�	�фR�X�uk&���h]�e��5�H�����Ml�Rڱ��	��&�&g�~��f�s���f,1�|!Y�}I
>� �5(�k�u�0S&�QK��l����[�Z)�bH���G��f�g:���6�%�8���rLwS�ME����%X��q-��if�ڮ$�i2Z��Nz�D�BC�����"��8]-X�8|b5���CL��7e|�M��_��b��F�(��8h妖��(��p >��L��Yb�qL؜���)G(]�''�t �2�H��RH9���蹬��3|X�eZ?|N�q�rӉ�nCF*�x=@8�N���a�(�h[Wb�ʼ;tL�)�-�/�{�i�4?��V3|щ�| ���t>�Ӓ��>��\bKA"P]S >����H��#:w��#��'�U��:LYh�f��2�q�Z��P�9�I�"N"F4 �4e�]�Z@���k�amEx�~��gK6eSg�".�c_�;�����E��jg��N���g�#�*&�D.�)Z] ��IGVNQ��t;1q#�z]-8�X�E��.rd��ђm-��S:��.�] 8�\)tR�4j9�5@���U�2)���� ��ju%��y�B�@�;�]��V��h��pc�.���Bn�����(2�6���/ _TU粶j�;#+��\���URC����    IDAT��Lɖ�8�6��PL����ɄbN?���
k�_��(�(��n9����h��z0�I�SWD��,�8Q|!��"����q ǔZS#��de�|�8�H�8�R�����`���~pr��g����������kO?���?~��W>{�n{��b3|ߪ [�W��
"�bj�a+��&�1���{�Z���\�6���$���wh�޲���ΝO��(��Z��ڰX#�rms�|��v.��xAVOL�
Y��t���I��Zd�O|a�zLv�~�[L�Ͽ��O�>��׿�������{/n�z�r|tyv����+�j\*��ȺN���ĝ���nQ-���_WI�Ǌl�������Y���,�>{��Y8Vd���k�Ѥ���g+j�O.�����ӽ�~����D&���S��H��FТ��'N�p�ք��/*(�qY������^��j]_�go�Dy}�x�:�8Y��o<+;�^/���/�����xڋ��.��Rຮ�s�������O�XO��K���i/4O��U֡�3�Fm�(S���y�W>�3-{�c�\��>k�<� �"�)�=���QEWD*�%���Qu�.����
)!ѷ\ڱ?�P�L�7[�eO4��OG]��ϯ�1�����ݫ�@�t<ҳ�bDtes<�=����/�O8�?�y���}�8��o|���ŋo���'�W���P���Agg�],�%f�R�����u�x]���ԡ��x�ӪG'���[���ߟ��?��ۃ'_]����{�}�����^��V���"�b9����~�*�o�<#_)��P���1������o�Euk��@�R����Z6�u�y~,�q���S|��	��K�r��]�#��"7���J���2 %j�������2E�Q�������G0e�R\3[��MW"h�WG�uB*�)05�d� ʐ��"��-q;/������BJ"K���V3{՝H�-c� 5O��e�o:tq�v�t:�C\���M�?�h�k1��{�w�rU12��D�K��_U�t������l��UTt!��ji��ۮ��)H3�u� ��5c��[MR�v� ��hT������U�:<k]F�Ѧ�R8�פՙNuVnQS~Y�t�EV~��V�e�<q!H�ҩ�"��I��.��o�3��CR6��*���rEI��b6�˵U�"���W��ŉ_��B�-�Xn�K��)rk2���cN�p>�F�A��8MN���ĔK1���sN����맋�*��m�*-˴�ʙ�$[A]~`��4%Z`E�!E��)�B�VQ!:II)+fC"�NK��4��C�T^:2�Z����ZM
����Sȯ�V�,�Npd�!lz'����/G��j/A#�ԭ���Vͩs!;�:W7�,
D6�G�S`�_��b*�z�M���e~�C�t
�1�:д�I�dpR�g�qƏ3+
ߍF��	�Z`!4��^�4gi��Ԟ��n������՝΁��B&qwZ��J�P	S�!!��j;��r�|�|Q�F��BM+�7��4��MaԀc�L9�hD�:Vm�VoQ6)��3-dd��e��R&��T�3��]�8�A���qJ�!�\����i+��lu�R(̸e��B�[b�z�٘�n.�ngui�2�	j���Q#>�
R�9��o�g|PJ【�xS�=4����H�󇳋 �R�!�����6���0�3=L�q2��C��\Q-*|�H+d��~���BF%p8,��&��f�����i@D
��,'�m+��k	_�(ܨtEwu�Jߕ*����!�t�
�·V�@|f���[���/�}
�0L�td��~�B��*��*�_����P�ϊJI?��2���2�W�;�̪��%��� ��iMU u�&�OG���G"΄�1őũV]����#���9t��㘶WE��u٤�ʹ��Ӂ���
���Oy���3"O|H)��,P4���Zȃ󵇜�I(�U����*G(?YHE�tMS�
ј��~���Du��)'�� M�kL���Vat�>/�+�B����R���o|d4���d�i�Y��[���猙
ф����WB�C�Y)�44V.����E���m�-�����6�D�ePiS!�@�dE����u���9UZ5�.	Qx=t	%��N ��9)�o�8�~��2։���V�x�t����L4�L�{Pƪ+D�34�|%�i�GC�MS�빢�����N
���.��(85�ޯ�D
�'�4!R]�������hC�BƺBh�
Ĕ#��D�@U�F!�K9DW��3������I-A8��r�����5E(w�R"L�r�YY��i2N�T�)2e[�'���!|cŧ�l�YK��6~~Y����YRFV�Y��h�2#�`ʨ��uP �|���=�x�o��͇���������y�y��/�����s��~_�ce��D9���sj�tU�.o�y��ј,L��IĻ���y뾞�/�[�)�	�`r\�:��LY��m���a!��Y�wb��,����ŁK��Y)v��QHKFS:��V���=ߎ����-��ǟ�����o|�[ǧ��彋�{ǇW'��G>5x��|J��R؎���*tX���Uo3�hL|����%Ҭa�&JĎ!E�s��ű�#d��S@��8R�󔎆C���ʑ�֓,9$P�݄0��������p JB04���!4c}��gLOO�E�0���\���>w陘����
��NZO���d�|��/3퇵�=]q����s�����>xtr�ٹ�A>�?�$��q��ж���*���]���I�@A�2ݚJd6�'X.MK�|�;�Y~ϟTA���c�t�,{�oK髋�i}�wl��_JQ�CG��S7'D����� ����#��#��������x^��=8od�n���
�g{p�D!s
a���f�[���^V.�^������������'�8������`�^�˙{/|����I��t�|��ku��p�g�]��^x��1ۭq�`���=�8?p�~���׎�x~���ʯd7WW'G�S������Q�m2}�ʹ���%����&�|5= ��l[�틋��NP�M��L��Fm��媫�Y�WE.2�&��=�"ÝGcU�ɴ��D2霚�&jj��X��:4B���	7m[����Y��Z����U)%�ӄsʥF��mñ�5)����Rη,_�2k!e�� �zZR���T�:��F�p����5���ĳ����N�������(MG��M���B� %dd��igt��.�AҰc%�����n�@�m��5�US�
Q� �Iu��+�(�8������.QQ
]3�r�#�rZ5)�,N�%�1�h�*��g�B���))K����  9����U�Q�V9p>�!ȍ��s�Y9S��!�@��2����A�7��
�5�t���t�����O���N:�5B�LV[Q3|!>��2GT9ے�")�J��%B8��1�7�����!�N˙*�9j!e�\Ӝw+��9��,9����[�]��h"r)1�Og��E��j���a�K��U�B��&��W]�X�!�4B}N~4QS>��&Z�n��17�Z� T�]�BD��/�,�����`J�Ŕh^�*��S��?����h��3��!�*���d9�U�R�㘺1Ga֥&���J��\{�@S�r6�ShF"ь�WE��1�fZ]|x|!�N���8��S"!�:�L>�\�V���󚌆���\L��"єߴQV)���S��O�v�M���|��dY����I$}xf��d��-�/=�rCƗ��!�dW[wK�(&�H>�o�wj�a�"U�*�Y)C��d|�i	���@�%�09l�.���G��P��K�n� |c�B�4�*Bq��ą2�Bi�V9Y��Ɯ�'�i�˙��D�`:�_�F4������ ��)%�3wG��hF ���d�8	Z<��4>��y�&5��
i2ȀR��wGx��^ʽ�����V���4��T��i���"#p*
G��Y`���5�f���CЈ�h����]���E*�N6N3B����dw��Iq�I��?:LY�mi�u �ժX�~U��8�v�Q���K�]"(T�NǇS���� ���;4_z���G�t���uk��BL�8��g�6m�n;Gc��9V���%�G��
q�ƗU�t|Fִh#Z�E�ԄX��8�L�ru͘�čx;�Y�Jlڷ�BU)D8D�O��H�$[�I����:~Y��s�STb!�,_���j�C-!p��~䘅BR�?~�
���9�Bz��ؔ?=�1B�2��we�2�)+B)�]9�:LxS�Y���v�!�8��ߔ�"�r�u�~��rC�R��
a�5Y`���Ȝ�5Y��pQ+5�)pЌ9�0)w7��)�#��?�^
l5S�Z���[i���ʂlٷ�N)�j�5>P�/�٥�kX�2_�һ.Ƈ�M�B��p�tL�FS+勪K�Mu�0�D��0E�l�.2�Œ�PƯ���%Ƈ��|��)��(4
QV�4�9�E��� ʱFNcm�ӜD�0��(�W�I����ed�4YL|E�1����9P����р]~-�.J��T%GtwQ@d]qF����D���r�,�h��%����Q3:ocѦ�����ć�V������������[�z��g����ϟ��<{;��{q��!r}p��0�����m��N��3-y[��?=�p�u���zڢ7|��Z8�h�4l�_)��H�{[��U��}02�R�����h S�p�\�Z��G3�B�P3���☎�V�_��� ���������Ǐ>�ã���ƛ>�I��b��zu郛'�>��������P���q!V3 ˁ�$��-n�� �C�q��m�BL�Q�Q��6�,��Iᐲ���ydo�s�M�D��Ͻ�/��(��l�_p���qv�bm"�&��9��J�p�b����SC�!>>�Ҩ�W�l������|����`��O�]�^�g������냋��u�y$�Onڪ@�����'6��������C������7~�����/��Y��^vDЧf�+^����}q��=o�@��b�B�sG�[	S���F���v�1l2���4蓳n�����px���h���a����=_A��G�~�m�=�t�z>gi�����~�_xj�i���z5IJ'����W��a�<o���\f���k�n�|�*��.���<���ӋӃg�>b��a�N�dO��
���^�.�h�����;��K�4}��z}�f8Z��>��Or��?{�>�{z�g��ʷξ��������g�\�]z��p}�Z���#h7�vX��lfG��-�:c{�g�g�]q$f.f�֎��D �{��c�d�Ѵ���&�����o*�w]9׃�*$��Rp�|Q�9w�qB(�Ƅ(�ו�BV�h����
��.xQ:U7
�2�t��d��|<eH����[��~�i�=���U�BUe���#�آ��X=Jw�֏&���.-&}���=ǡ77���,�/+Y�4݀��O�������o�1ۨ��F��'9�@��$K�������~u�O0Mc�l��A�ѯ
MSQ�	��PMcB���L��K���O0��!��N���e����L�૒@Qx�u��4���a��VJ!R
9&8�}�6 �iޒ[��S��8����q��l�@u��QKH
�~�j�(d9F����:7M�X��H$5�)WKh�z�B�@Y�J-!A�M0�RpD�NǈY?|Ա�qQkO�A΀JW�,�+-�Ðc&b�q
����UF�ix`Y�a�p`u�U���MqT���B��s�����1�PExk4�l��q,*S�iTe�����C�E�)����i�H�[�B�$�2n�A6��U�@�L���+�2�K�,
B���h�r��g��C�C��0��l��p
�DbI���c:��V̗XK�gԶ(}�tt��#e�p��i�. �����d!�)Tb[�?�I�UH��FG�2BR*M�z4Mʈ9Y�o*�_{����8�p�FY1��@�h��Z�K�'e�Y�1?�hE��U�VI1������B�r���c���#%�2YV�E�-��T�?���Z'b��R'E�����8�##0�R�Ƈp&ʁH�ꇏç�)���C/�cQ����C��a�T����tj �,*ex���2h��49�{!��,L��_�	՞)�D�B��)We�q
5�b�G�|�͟����YW�[�G���BS1��)���RNm�{��)�(���Y:~���)�f���#ptb�O��.���KQ4���)�A�`�N��8�V*qꦜ,}>���$^z>�#�����7�L�Sc��۪��4ܔ��I�� 鴐�|�c���ϤT.A!�\�_t���	�1nb�)]6�l��+Ǒ;����T�h�r+dd%r
C:;���k��Wsa��JJ(�X4�:��@Xk���.|6���MC҉D��G���L�𤊚2��/�,�:7-���&%�U�]"=��@X)FQ�L�	�6�R��PH�hL�@�Һ{5�@L���$����76?���Q��Ϗ�D [�:VF��8�%k�J�E)��P�N�t�$^	»7�.�O'�.ڢ!IIכM	�E�������$rB��ն4�h�@drq��Q.Դ5F��*WE~�D��h�����Mq�b,���*�^��H
�J$��i���.��Q�����H�g��Dj���]��CM?pd��Ù)&qN8V^�D����,��n\�w�c	�a�|4Y���@f
og�o�0��e�V������=1mQȌ`�8#�����jrBh�V�IjuR	8q�n��_5�IGW2	�"�[����Y���)*��2���[S�����P�������勃/Z&�ƪ�7�ZKj1�Z���Pq@�bDn��k�|�(2���j,�B��7F�{|���ޥ�Lu'�G��������}�������>�̻K�'{��;{��OAi��z���R��7o�*GӊL�5������{���A�G��쭷�z'�A�cCz
#�� oM�K$h[<=�#�� �y�r�`+p��:�Kg��g�
y���QYH	�����H�&�@�Ȓ��������������g7������G�����o�}�̣��C��|~z���\ាxN��k�̚�R���CS!�K�����^.��"�G�l�d� ��"�5Zlۂ�&�8v"R<��8Y�J�����:�#0\
]:e�h%u��<0mUJ��@
���e�s<X�b�=���ۯ�r��˃�''�����_]\��K6Q��#�99��:=>�AZ4Ƿ��q�usx�q�����_}��㽃����������Zo��IYv�Q�5�g���y��Ù�����Ǆ���б)�+4��z�96�%��n�]y��L!״q��ð��:'Ꮂ9>O)�<���Ö�X#�{ �I$G]鶔�'@o����=)a�AO�R�鄈,��o{�ӟ���?�������c��zZ����:	ϖ]��������sP}�����/�9ust������g�ח�Ø�G��g������{/���G����D�7�ׇ�=��œ㣳ãW��ݓ7�����x����{g^��s�W8�qnȭ7�:���3�n���03eb]�g�ngz,m��)�׶���\�(dft�F�tLhJ�E �wy$b3�FQ��.!!WE:���j�wޙ��#*�D�R� ��B��%Ŋ8. x�E��BB]�.E�9@���!Tň	gpRB���"=�u��ܒ-�(�V������
ч3��Q����ç K�{�kiIi��qT��]A�YH�"+d����y�SȊD&é(�z�NM.}��ٖj[o�jI�Bqdq�?�9q8���]��z��Lxa�(ԊVۉh��&1S�l�U�!�TW�]+�m�P�r��Q���Vg�M[]x���RM��dӚ﬇SH���p��4����[���J�K,7�,��V%H!
�h�bJ�����[ʐ��د�    IDAT4�e���A!�@Q#��O��,�9bZ���4�ŜZ@~4u��$�X�ܶ�k���8j�j B+�#KȨ(��BN�M�!t���!��Sh�c�8���8�i#��-=�t��YKtG�
��)�!g�nٴ�A?5 ʩ(���s�B��L�'�r��ǈ&RzSj1�Qh�����ёbZW���sbⴺr�nH#M|V�e�L��*FfZ��:������#��t|4>�bv�D��U����Zr��Ad�ʇO'|`L ����J�'���T�^���ڍ�FHE#Hap���uw�s#l�[��h���3g	���#%TK:	l�|����d�i4�~"T�:\x= C�i�6��I"�[m�;�d�N9\4�G4�V
Ac#�*Z.DV�ʅT��B���`2H���ElQq�E�K�$�:\X���TtZ
�/�e���^]�z1�T7����a�Uր��ӌ&Q��(��i R�Jd�e%"�A�)p�?��ԍa�5f4g3Ѧ��C�S��p���B)`�
�R�j�����O9���)C���G6M_�7�Df2E9��ٝ&b���STu��D΅�2�]5~��V�J8����̅�4�K)#ˡ!)��l?	�ъ&^�e�X�3�����]������B�/:���63~-E�S'��~gN��d8-�!�fN�9��k:[��̮a�W�|d�-!�t$�12R]�#0�1�L'˙f0E7�ۃ3��f�	�K��	6� K�s�5&�ì�@��+d�%8���IYM1K����~����I�[�n�"��yN
B�\���ʍ��ڈ,�f�c|�����S�YV#&�(j���)�BY	N�J����NVCwF
M�[r�=���h�Y��#��fǺzG�2�(�_n���+��"�["���h��k��&����_6n��I�	!r�:,Z�T��h�gZY:,e� O9���3MOQ�A����@S��~ä��x���8��:�O ��)���H��i�����ފR�p�-G�����D!L����MS�*��f��5Ef%�����B����K$'�����E�r��TW
���n�rU�w�5 ghF)�l94�>��H'Y�1�j�!�]n?;�%XW��S>GV��Y�5�2�B��(=e4!"4���\ �$bʯ�tƑ�I��]�@"��T4��2�mD+�)Z�wi��֫I�eK�`Vs[W9�h�$*�_Դ}V�_��i9���+�hRm��*�uXDl�^���dwnߝ�y�wv��O������������[�ǧ�U��#M���l�#ڨ��)�"o&���o����-b�9{���d�.�G�l5�Q&o-F�8�t�@_!̌����AnM��z4`�<<��no�����V�C�!PP��m{�L+�2��J���Ӷ��32���?9:�~������/�>�~x�3��{/|~�ө����]��_���a!j��(A��µM���Ҫ�S�M��F8��Օ]
o��7�hrd�+$�{�qD����#"n��7��x[�3�P����<�9Br5L��T���L��
��<jQ�.��琒bd>���O)��#�ح�ϣ��s��<	�x��^9�5���]�?__lz�{��/�ܻX�;}J�gz�� ��?={��yz�}u�|ps�S��o�*T�Fo�k��&ub/쑵��:��72���Hk�}����<���������Z2�vZ���G�*�g��RZ�f i����i���)���<K���g����̩�֭�z�d�#�.�����՞��0�Z�n6���l+�Z
�2�\_����N�>]yv��s7���?=>��O�/�����|���Qa��ugW���;�]0��_�>�ӚW>�yst|vϹxd��l�w�������o�����7���ȗЮς:�����]�8v��**�.�c�o:!�o]n��nC\m����
!{bdR$�'Ԕ V�&����� ׀)>�r��&ܽ��߈�D�y�L�F֕Iǩ9ji
��s�]������+��]T��Nz�D�,!~U�'���H�Ԟ���BX���J�SN"sq��U F��2U���&�s���E�
�̴�t[3��b��԰�[�vU��{D�z�ҭ��K���QbR8��2m'�3)M�%�L���f��k��ٚwk�PW|�UUN�Q�DhrL�t7Ł����j����HY���T-���b��*Dy�A���bDX~��d�E��e@�u����O3�F�vCV/���m�鬋M�DM!Z�Z�XL4�(�b�w{k�N����|�Z�r��W�i)J�YmsD�dE�pںB(�f���#�Ҕ�m�֌,����8j�Ԁ=��&E�_JH�`4Ec�,�|�������#r���E�\x�����!wO'r���E�\���JWq�.f�OҦ�g����U_(<�ڐs"���*G�7F���a	8pc��_�3Z��G�~�9S�*$����2��H1�p"�!hh��,������,�Ӯ(^
ZLSF<�tB�Jg+���(_t��V�8�h5�?���K��������\Q�Ub;�>���͊V�J��$U-#���C�#�c�E�^��pҏ)�mZ�4�9�j��tr#�MʈV'����D�<&0NYq�-DS�d��Lє�v�+Ϭ�B�Ԉ�Ȋ�4-4LάŔa��%Y��X	
�B�j��Ԛ�إxwG�ZW������-y|jSڕ��K����iH��Z���"�[8_���
��m��9�Adm��	L??qY8S+�4r�r�6�S`)������!Sb���9p1�U�Cgơ�����BN4�(p4�T�c�5yJ��(�!�#dƙ�8��J�C���B�ۖ�G$'��M����&������yD������ܤ@�kQ�����]��j�݁z��4�_�_Gq��X~}��(�Z�L������A��[q�1���_zb�L1w{Rv���;��Qȗ�HO�9��8��9�R��H�iU�R�HSNDk: |:��L[��ݒ��]:�Bޔc�O<�hVK�h4~�F�ɝ�}�E"P�:�)���p�r��p� �3����N�/��)_?9��7�l�M_��s:'r;F9) ��#���DTou7�%�i��|�,\b�R�̴�����%T�Դ�R�\.f�8��vȔj	�j|rN]�>�V�/������*e�2�5 D0$~S�B�)w�!+D$�����
oF���U.�*pјU�tm��`���e�L��LQ+)���N8ꊦ/�S'��u���heSC(dqz��)��uh9B�`���/d?�i۔_
Ym@��Rڍ���b���Vd5�D%NmP	8&�d��!3!��>�@Dn
��R��e�Z\T:P�5�G�0dH��z�^I�c�\�3"H�Dd>�CD�ϊM0U,]A�ڠYW�5�B2�E�d�1-��
1~�Y�맕*�d����NPi���)pp�y���0��)�r9je�GDL8�[�յϸxT��������c�}��������|��G���{W�<�~��74����j�*:�V�Mfo5{z�+o�j���}Zo�z�a��j�vor��㹌\�B4�H���;��)HR�����HdB�.�zLR��P�<EnU��k���A擢�On�!|�(���׌����Ƒ�ζ�m���,�����__�|�>���G�����>�wxs�?>=ٻ���%�n"=w�Y����+�_E!Cc�6�i�_���tʚD �1%�<���c�U��e|%0)�N!�BFR�X?6���"��;�>��[Ԓ�&-����l��@� OR*/���c|!�Fks)8���f�������`��`}���-�q�k����c-��V�	�ZRt���=�'���><������߽�������ᕵ�wz�������V��G�҆&�BӢ��6^�J������<����<�VҴ{.�!Z2Z�ꁊZ.n�R��J�z��(�����?����1�s<%Ռ���m���>��Y����?�ɃO�w�}��/:�*nS��,�C����7n6R��Z��5*�U��?~�������{>���������W^�����O��Oο�������Cf���/���|��Ϛ������Ŵ{��'��mN�Ԟ������kڵ��6�f���������3�׽:�������پo,���ṏ���T���Ik��]Z|2|��)ߒ9cRD�X���oO� ����^��KVq�r�F������5j^c�zK��L�}jL�3�gW_T�6��6D9�r�(Q��,��d��*�d�0C(
��+:���WKe�>�����d1"���`D�[/��P?�$eT12Y�M�4�c0?M��m�MCp�[�D��H�D�,A?��r���`�q���-itÚʅ�$.%�� k���G}"($� ]���7�"�9�l}�$��V��~���Iy7�=��P.N#Z�����h>�,E.K:Rn7��-BhB�J�/��d��!Z�I-0DW��O��#�8�B>�)>B��Cٔ���.&� ɯ
f�ߎUT�*�1�,7YS B�����C
r�('>SYSW�JG`�,�*�M�=��B��/�Ι&�8���'���R�lt$��BE	
�#���-�/�?Ԣ�ö:���.�ZR4�g4�9�+S �"�ԅQn"��G6v��gC��˪%c��٭�tup���U��a�;Y�F��4��zڄoE���Zjxʙ�6§t�p���m�F@�.d�B�w͈�f=��HE��8�Xug	���>)�s�M1#h�_B�=)
iE�Ñ�LY%��r8�B3�H�o,]�%z'ˑ�c,���nW�\c+��T!U8,���^�:)�@S��|����AJ/T�.���p�� +DCf�3�w�r�[��d�U�y���]��1H ,n!�	ۯf^�{ :@ſ�8��nD�HtCH2��RWw�m~k���3�I"��|��\k�}��,�S�h�R^r����_4�&s�� QJf�@>��tj N�DN�q��l�m�t�H�&1�a�9FVoB���ZN=P�ϔ��0�uqY�XE:�Y38� �Xu
���p �f��V����B��m�F�g�⧐`Yu�g���R=��O�h��-��r��K�u��ñW�(TKr�P�/�K�&Ǐc�>>N�:��Iak`W�('f"1���T7dp4>B��@��FH�n��
��]4��L�>��<�Dsfu�w����j�7�c�� gB]
!F���FQ=�A8��RK���!�i[��C+$�!����o
�iI-Q�~G5E� kۆ����7C(@j�3d)�s"�֛�*�iV�t���X8&0f�6��}���k�H!B�p8n�3�̯����x�H�?�j��bS>+{�S���P��-?d�oms�8#�=��.����e�������?���G+w�(��NWj@�-
aI�`0�Nn��.��V]?D���	�n{�%njӄd��h
1�J)���CZ#�K�J	og��(]nKй(�R��BL���ȩBx�1'~j��NѦ�~�&UQ�,�l,�!�&���G��ڬ�}�1F�B��ԃ1qd��,QnQS&ň\�F�y5K��D�p,��
1N�p�uo��.�A�	ޔ��d�*D�ɶ�)��Bk�cVH!�=1V���� 7z�W����̔��C��M_c�|Y8kL��8�a2��i��@�Ju�L��L� Y~=�́3Rt���||�e2�7:"� �s�#�&����,�Z�`�`!��F��С̧c*
1&�#��.Ħ�D 4Ó5����"��,dՃ�j��!�%4���Цg+�@�\~C��d���3�&��X����cg��p�����N+��?z��/>r���=�����;�.(}
4{�ubZK~3a�)�+4o��H�s'2R���4�y3�	�;�V;�t�e	Q�E��֙�DfJ�x��Z�F��Zc'2�(�"�$�������A�
�;��5�mW�=m#�՝����5!�Pź >�fo�)j��8-r��3^\8#�'��������>����W�������;�<�wpqp�+2������O��eg��>ko�=$�ɷd>Ά��m2�::7m'1]K�(-��o��(_G���1>�]����u��|N��6ӆ�Y��Y�˰���]I�t�:Ц���j�u���	�S��5�H�ID��H�\o�]=;[}�������{��e�M��m�^�.�y9��.�o9��8�q��g������o|��z��߽����^\���p�cͧ�[a݅
����6�i�,�r��s�Q.ӭUX/��㪠Ab����$��ǿ�M��,�Ѧ�i��z�=l��Cd�:q׺;�#ڜnq�B�1J|d{��=��i�����y`��+��uE�hK�K���������>M��=�}��ƺ�҆���b]M�ן��S�ک�O�=������޷���������S/e���3���ol���������Oٮ��1�/�d��H��4���q��|}.���ˇ���7�ǫ�~��_?z����|������C������(��m��s �̆C�8m���uq�j�܊v�V�"{��[�������i��B�1���nY�`Z����f��h.���J�528"KQ�k%\Ec����q�P�K�K�n�:�W��Z�e� O�X��ڛMv7Uō���I��@_�JM�@(�tU�^� ��,�o�R�n����\R�ڛ=���V��7�(0
m�(���V�>�,MG��L&4Q�	��֕n=��A�����R����M�rS�s$�7�_B��r��!�N�(�V
m��M�8p)�XRJ�խ�hBH��h���إ�,�5��Q�LAVQSN���Ϗ̀Jq��2������G���C?&
Ig��������1�+G��0c��9�r���|Q�'ڢ"׳����6�daj/�L�P}b�2
��Gm�%X۫��j�I'�"���A&^�ь1�0M�Hqp�/���C0Ղ�y�P��4�H�[�%�
�˝FD���q|�K�c�|�|c��W���[�wǔ��\��zB ^#�S����hV4B������
�(ӛer��sL���;P.�rE����}R����ߞ#+Ⴎzw[?�&�D`;V{�QQ�h�F�4�1�Q"2И&��9�M��7fE�0j3�VjF�|�Y�n$��h#5֕""��F�PS����	ǔa����)k�BU��GNa��2��\��e��Y����"k�DU�p&b��M��F���	u�d�Lv�E��(\
����O?��+M�U륶�hۊ��Y4�,�v�p����:m�A�5�'D.����Q"<q��+�Z
��_�\�8)즣I1�����'[���� )4&R]S!Lﺠ�V=r?�K���4�:��	�nW��2�u2=`BZQ#�T�n����ar*ݘB���f��X���s����hxc! �ÙЮZ�/I��%Y�ݭxI�4�q����^����?��+��%B��il�1]MH�z3M!r݆O��ѦD�p>K$ΤWb��R@P�qD�B����ʷUX�<����H�	%�%{A`p��8�=b���U���p�4
qX�Q(>�����t����F>ܘ��8�q�tp�n�/a��L4d�/�h[�'?e���§��W(���6r��9�hR�%_W������8L�,��p�u������u䄤\��w�K�;���}U�ri��:p���0��0��&�t}9�\��u�c�C�1'�Y9 �\�~�&�S�bj��_!��uGP:�Ǒ+�o-M���D�ϟҦ!F|�M0e�hS���(WJ�A�ڍ�M��+!���4�f{�@
����#4����'=pX8G�.��)�t"���DLUd޻s!C�Y�h1C��_����^N9Ԥ ��\�_9��SAk7�w�gg�%>L�h�t!8�zM�OS������~O����C!�pNH~M��!p��Vo�%��    IDAT��:��	231N��)%G�(��IDh%��F�N�F�ȢI�'.�NI��~@��#����7es���D��놗+:?:���<B�(�8�8]ǹ�S�
&��VWFh�@?�/Z���h�z�Y��8|���N`=����@d�ֶ��i�dY�:�BB�<�ނ{�{��ԣ��{��hξ��~������@�#����cj����x�6�,�6��QeZ��c"���cf*�m�CKs@���6�7�ۍu�����V����X�7i[��ma8�w�f��x��ۆR0�w���>��>E�RH�p#_QR��:K���_�h:"T�B��O��t�[l;%�{R�.�<y����g��Q�񃣓��j�ӣ��{�'��������'N�����n`�bdB����tv��~�ZK��Zp1Z>���`꤬�8�j�RX%�]>�H\!U��R�\ΰ���<�7�xC��^;v��ب�Mp=�-#D����(ö��}m�t�A�ѐ��|Vh�������:�ˉ����G��[����2מ%:�tf���m���O����!��c�(<:�_<:s�_<�d�C���ٯ6�i�v�}���:;�D�5Z��	��D�-��g!���L�ŗ(����`�Z 2sy�
�e�ܢ��eW�U��:���\*��C��ȧ����uy4��fZ�Ҕ]V�)���/�������?��&�*'e{MX'IO�ί�����W�.^{����'O��>~��ѣ����]���������0�Ӡ�e��2���z���c������m�·G7�W>ع�.������ztrp~���W����O�������km�k�?帼�=�q�C�尮���R�7x;���F�IL��n�����*hM(;#ʗ�L�B�����2S�Iq�UH��FY�KU����t�Ƽ�J$�!j\AM��'D�X��Ș�4�Ȝ̽��[��m-���B�S	�D�׳E�Zܽ�8�Ɩ�M��p&��&l��L��sಌ:!�1Y� 4�qB��5m{%�uK�eVN�IGh���L��p҄t)�p)�Y,�������s��4�m]:��?Ĕ�t�	�%K�HQu)�uc�2No��'kZVS#��M������9hF|#��o]�R��� 5�������v�q��Sn	�#�Ңf�n|"�
 �.�m�:W�oW��+g�Ֆ�J}mZ�|�|�9SVQ���1�:��W+~���]�_�t"׏RW���h���`�/�h���j��C�LK��hC��8Qe`Y����	�p�ȁ�OM�O��#�t�\����I�ˊ9:1S(wW?�@S����6��Q)�I~"]��̈Iǈ� ~��z�"r��XY=V!8�RF"�S��o�Lӽ'%N"5�KG���D�~ ���#X��A�*�>��zHs�e�����&�>�(�Y�������	B"�徴-@F���Аk�����r�� �6���A�@]IG��Vn>���(�1���3Mf: ����%�p�8|��z0�ԕQ�y��au+�4.�͊r�L�]�rq
�|!~�B5�M��h�h1��k
��L�@
��C�p��I)T!�~�������uI�r�)Ǥ�f*�~"���7��a5&+g�#��D�ˢ��R��7�5�q�p���9�DE�Sp��1�BF�t�ɔ�g���c�Z�е0姹�S"\{�9�8B�z�b
I���*��V}�w�㷓])!ȨMzM&���H�����"�Ù*�5����N�(dן�PSk1��Rz���gӆ�,ܘ�K`��x�Ij8|)]2������"�el����2Y�(H�'�Y�1�i)�!�<x�1Kb�F�D��Z4�l��62�#R������B.H���P��>~�#���Vm�VO�7��t�|��h���\Ӫ���O�"e����8�)��8|���Ѭ�DÅ8�#1M�\`;���rvRKu�'�9}�X!�4�X.���WW��Nc�×�&H��8}rL���8���B��s�SS�#$��S�0�!G�P�F&��3+���J����ȶ��$�t��'>���t�sP��`��B�	N)�'�6�C�S�D�1q�Lt�r�ހ�
�7�����n�I�7���M�n���j�.��|�,)TK��IaS���o_�AZ2'��FH��᫕_'�3����tR#>����2�)亘�6���EY/�����#ͨ��9�ƈG�2mת��O�4)�>O�tj&~� �.�6�%�.��!HA�QS)!���nʨ�1�Ѫ[-��?�(�B�m�|������b���4
�-S
��a� ��k�ni�2��J����pZQ�������n>��E6�!���`�j�h�Qg��6gw!�F��)��$�OP�)�e�H�t ����n�~D�n��/�'�S�,��ɑUJ�Qu#�y�"<S���N����?w�ޯ>���?=~��|�����,|���z�M�O��ڲ��tR�	o��s=N4 �~�׃���8�!�7�#���,��Mu����x���l�Dk�U�+���[�r[���@J�y6Ut�t*�؏S"�Z�	��<ǧ ��kF�[����Ckt�Z�rei�&��+>_�����|j��O�/�E�����g�>���"��;Fy������s/l�'�>�v�f��=̦�-*��ن��X�1�#)T-LK����~˥is��ҥ�!#X;�j�:��������9�!6g}+qZ21F�D-�er�	)-BCL)t9��A%��ޗGp���w)����:�8�g׎�.�ݓ�]9�D���M'd�N;����y�1H|������/���ٹO >uc��t~�ć-;�Q������;�ҕ�#��Vd�TAh]�N
|u�]�B8�n��>e�����}��A�%c2���sL�����`tl��/��/E��y�-��(�獎iGq���G�wޡ��x~hZq�(s� �j��Q��~��_yT �>H��Om8:e��!����^^\�?x�o���?nzvs~usu�����o|��ѷ�/�v�,��\��.�t1�%T�v�h��^݅���?��	�_��8Wۇח{�F�	ݛ�{�_����O����}�����o�������l�`�|#K�h��ݓ��P��p�(α3�?��Vjբ��G����pj)�
*J�!�a��m��F���&1�{�����VDs��փ�}!��>Wn"�4�.�I匘D����� ���ժ��M
�\-��D���ў(Īe�n��x�ա�BnKQ˯�*N�.Y����ZAUʪs4�v���j�C}ᰜ���8�a�%�	ѯ"\	:�6�Ԋ���5��iCHq�]&����jIH!8���'�������$T������gM2S=ԛ�����!�Z�a��,���O�>Pu�M��h��&�~hC�MK�2N�vR`���"� ��(�l��@*����\KtX���0�"�%%�:!�\!���o?C��ucsT�!�C*�B�ͧPtDL)T�X���ҩ[H��)+��r�FQ���1�K�׏Qc��EM�2N]a���8��t �1�����TG�E�l����d�hOK��c6�J�U#(�d�^.�� �S-��Z�čcS(�z�S(��c��	EMN#���Zr�V�QTƲ8h�Q�"|�"%YH�HQ����*����'_.�h�+�&ME�19z�"���A02�I�D[��RL���rk�XQ�8��+m�z8�l
�{]�?cjF)�*�LS.5��Wc@x����5����(��a!�$��^��@a�mM��s0)O�ȭH�����p��fZ�������/�mi��r���M��Ut8[��8h�8������V�,8r|~������6(����ܔ�(�5\u|~�IDvE�+�6
��ҩ�\�5�h#N�LY�Y�Kj�H���r�S�t:���a���ctW�L?|e��:�d��v�Ø8D�鿴.���eFV'K
��2
5����aj���:����~4���l�B��"�l�r564N~[A�i�C�����ԸHw�6�r
�:|x6)) C8��v~�uŇ����ɡ�X��'20�9�h���btr���f�%�Q���Ws��Q�&J!��~i┻ˌ���\ќe�xLё���D$�3��H�S�Жw�ۏ$�)]TVϵ�j�*�_�n�۴ܞ��WF��⤟���_"Z;̙��7�3Q
Rk�E��8�GVV!���� 59�B@���.��p��?yt ��G����͡E��@�|�������B�n�K�ZUG��6 nT%������u�=8��7���x)���>�\�'�ϒJ�U���ƪ��DLs�$��Xx�FR�@~d�|�ަ�])��n�	�š�8��ƈΘ~Y�h�B�6L��R�O������Yo��I��R��A�kf�����[�z�U���� �t��щ�:��|8�T��Ѵ�u;�\H�hӤB���8F��i)�)���+�[c��oL0_Ȓq��3�8eQ _�@�B��ki�(#[{�  �@�BI��\RƢ)ȢV.�2R(Y{r�+By�Z���b�ۨ����6��D��'U���,~�F�D�$����1��%��12[�2q�0�&N�5���E5 1Z8#.��@D�Ĕ��PE���]A�1�^����Jo5o��pj��Q�_)�i�3-��ӱLcK0Z8\b�*����C��V?|��Ff*�2�_ѴiN8���V�����;~�����߾����g������	(�n�;� �j̻X�V�z�lOMKC���0Y-��x��g4���{�b*1Ļ٪�(o�M�ŨE��7]��6Ԇ��.�E9ޱU�����~��#���{���p7O�}��[�-�z-Si弙o����.f�M�9B�H��bz�����֡��Յ���>��'W��y��������O��^>��z���,�gۼu�1uu�Ҵ$ʗ����SQHY��%���B�T�5;i�]�(?�B�85:������Uo��ף�$s��T��$s�ڦDш�7Z����&J;�<���k� �٤Ce��;ڿ�/�d}a�?�������n��>��5���A�ѫ��O�Ƽ�x��k}��Յ��O?��3�9KPuv����X��ŵd���h�#sp�O���z���mB�H��|��������?A�n��(L�'��M�)��}_	+ݎ�e]K��Br]3��?��#��fL5,�s�;6=-'j��霈��&��Ithg	�ԃ��
��ri� x��!���,�������{����>���1ƫ�����������G��:z�wr}���ӯ��8����/�
?�n�|����#l���W�o����>q�i:>���xv~vr���b���ѡ#7���+�.���ŋ������Q}�t7ֿM�*�>[g��~ZBKF��.��a.�S�*��pD�ȉ��'BMԕ�i�E;	��s�Z��cn����RKo�@�*��|�'.�}���⺻�l��m�ʪ�Q�ɵ"�(����ā�li|E��1��B����^�hX3~��t�,��E�H�}��^��0[e8��BUt?[�\♐���.�M]�L�H_����#K4{�	�( �q��ɒb�z�B�8�dIOA?��F䍵~${�~��߿�B!��ZP�Y�BFH��NJi]J�@��q��ch	|���C�d���U����SJ�d�]���!!�k�ˁ3>&�	՚r�� ����Z�;�|�Kq�
!)�j���j@�8��B�ʲ��$Ʃ�:	7�A9ùso_[�!��b��5Y���B��c���ˏ�ɑ�҉�(�&�k�g0c�.�䒝���UԔuM�����|�m���U�����H�g��y��q&�����/E{��@��v�/���KM"TȘ�=C\V�B-V]�i6m��/�4��|�@ʅOVRFUp8ѨM(2�T�� C�д%�MSY
,~OA�.�D-\(&�-o��|#>�!�,�q�yF�P�8��U��!UB\.��D�P36�5�B�@�B�)'2|4 ��P��t�Cb�c��ɖ��0�5G�L�L�J�sRG6݈��/8�
�T>E��v�e�	H͔x�-3�h!U4GJ������,�B���A�J6MjRj�Bq&��"1Ӛ��N��2mi[�j���W����0>&���,ZJ� ������>���o'�@X���d���wuD�GK��dhQ~��p݆���A�\�FV�;!+Q��� L��E�L�!h�J�0HӔ#S��du�D��l|B���
��S�mY��b�Nj8�MSp̖�&��%�nJ*�1|ڛ�P�A8��zA��I���2Q�K�v{����J�J�	i[R���TȈ���8�J��1��b�hK'�X�3�30�F���gp������|�p��swM��BX4c�M�M���m��zv"H��dhF�I}̢��#��D�'�̯�!�+�>�.YS#&0�1GhJ�$�2�UkDY>�qs�
��} R��sR(CX�a�5ٮV�SL���
F���s3�k�l*��ঌ��ᴇB��|��OGVSե���k@u~�j�a�ˊ�)*��M��Gf��5V:�PSx�)�������K�i��r��Z�)hXJ�,�P4YY[���h�J���îNd#Pz�a-��>�7E�o4e��A�!���#Z:@N������S�n]�~������84�EƜ��=5��1�U
��B,*7M�,�l�(��a�B:_-���z��2֌�����@�t���p���2��*����"U,�2´��	�����GhL��롢jѷ�V]3)�*$kH�ˇFdg
ds�(�����(�(� �)j*=�L*�Hx����|wO�2d�t��嗮3eB)�M#�S�ۄ�A������
�X�L6B]��n2�^�D.>�w�j�XQ��p��uh��D)�U'�ε�m+k��,Ƨ���8���J�9�Y�FS�B���Υ�ȚkTR.Y��';"�ե�����*��=9�	Bp�;�qGl�N^�]^;�qF�p`�7E����@Phý�%��\���t��P�FoYK��]Y!Rp���G|f�[����Xo{���ށ����z�Ҥ�z3�[���~������;s�OY��f���ת�e�_�S�Q�H
�U��ܐ�s�څp�/�^���\�8p��������G����c������7'g7�}�����Q�X-�f�V�)�G�QS��G�)ڢ�0C])!��X�*�%�6� �.G"���>�j|׋uh�b�G�Qx��+�Vy��5a�P����4�Dg�m�B����u,�@�����W�Vlo|Rs��׵�0��_�A�u��<
�4�]�\\�<ߵ�|�uyps���f�N�>:u�~���Q�z�\xqyyN#�)n_mXc-�6��g?��E�:�r_2��6ӍhiD���,�r��cnS
r�Z���K[dꙁ��i:�t��w�w���?��{�׏:���p�|�v�!�r������������U@��IEҞ>��x�U8�qY5���{B-K��4;9>����Ϟ�������WO�=}qq|���+������g痮��O��=��o�җ�z��Ѽq�n���e�jzxp��:>���~vrx��`����� W�^�����������g�����ا?��=��~�����~׿źv@NZ(�i��@������+�a�(��́S@��p#�&��ĮWѱ�]+�0�p����6��꺠����J�2�.4�W[�(��t�(�Rڅ�vq9�t5]ֲj	�{��1��I�j��t{(���Dp�Lb��^%��Z�V���(���G�eR3�J��QԺ"C\&��P��󓢯
[�����!�a.���BD�uE�� � DFA-����������m K?*z�Q���㨕&�5�\[h�B��`��1*�o22#q�9>��1���RTV8��)\�?��W�rRp Ɣ�2Ym�d�������"��q*�r�g�ҩ�$Mc�:.�    IDAT|dQ#Јo�~��	��s�s�u�CDnۅf�Ќm)2��3�%FN�i�k�o��K�R������u���OKN��D��X.2N~ݖ�TnBLSC�_K@�ͦBь|���D�X"p�i~���pU�*���p`)�9����X��T��K��,>�)撸����F4�D�j��a>����^��F �P4��h=T�u��m�#=5Q͉r��<L8Ĕɪ�j�#�b� ����y�1!�Pk��{(8��F�[qt�7N�Pz�� ��s*ė��8�d� 8�[��_?h���͘#��FYk�No����L���ԡ(juwe%z��QBL9Ɖ�QDX��f��)��(�Fk:���ƪ  �����'�VU�1�x��$����*?�쮑�}���,~��a��m#P�n��#�uME4�ٷ)��Pn�L�FY�l���(�b���M�Z9!F D��#��B����L?~"`6�S
�p�R���%��ͅ�k�gCN����D�� �o�ht8ޘ>�N�p���I͔c�V���)��P�Wez��O��i��c!�0�9"+Ģ��8�^
���;�D�ǧ��I�)4Y�h��1�p#��-��*k�Yid��w�C�����R�M�>#L݊���,��Z�F���nD��Cc|̲l��T�r�M&%Y�\��RF���p^*���ɊS�1A����&��zw>�BM��2Z{��n�|7���|
�@N��E�*	6�4M����D��kʗX��S����0N��D�I!��d���ZIaM��ol��:A�OcHS�Z�l:I'&|z�0Ӑ|c9mT��1�DZ�t`
�R
��o�)]H��t����N��d���L\�h�p�rE�rcV��(�B�*7�,>�%07*:�552�+7m�"�n�T�5i��UP[��:x�mQ� �[���LA.r�he��ŏS�|����ӬNړz�� ��C���t�rw�tʊ&J3�(#kJ�h:"��u�޶������0�.�tYԀ��Z���K����EE!BFj���,�=�O���yh�Ji'�n�Rc) ]��B���j�ç�I��rmE�"���������B�Xkϧ�h��A��h
deS��1B�̴���P�	?>ǻ"�}���)%�nJY���������
�	��L��Vr��SW:�s�s��gյ�@~UH�0�Bp̕y�Wp�R"PNs�L���Sʽ#��t�(0����ͳq�0����\E+�0EE���X�M�W���� O�$K�N��!8v��J H����@&s�J>��5d��t�����|���������^q/=~�>�sx����JפSʁ���h�M�K�E�	$Ԓ�(��K7�4���Ď�%.����3AQ�{c�oi�����#��ܯ�k�B��I]Q2���R,�C��$�-e�0�.��I��o�.�o]�5�{�������/}��?~�����b�0�x������7O}�p;i�
:��z�-�M��ߨ\�&-�i��8�M�Ili��U���OU�J������+C�pd͛R��l�m�� s������2�v٨�oP��0�Pm�gU[dkj����� �0���C�����?w�s��t�W��H�]�Ze��v{l�c�>&���!�O2���^_\�e�������Z���������oG���u��A]iC
���}E��~�;!��[��PǱ"��Bp#S���>�i��FK}��/ί�k �Gڛo��Ӿ;�wӻrn)�'?���NAT���Q�wJ_V-�
\~�Rz��w��LE	~�{�sP���K�w�ؖ��L��;E�d�z�T�T�щ��~�q�x��O|�嗏����_{��7�g{G�~��kG����q��'�?���Ń�^���J�[u���H��Z��O1�n�\;%��~=ڻZ�\�����r%��FG�N_=yx��=���/v]{�p_�X�S�F��[��?m;�+��O����#�,��є��L�閆3�����D��L��vSM��n�D&���I��\h���Bd�����փ\W2:5o�AFsM��_E#}ʑ�!�2"�E��hɭ�+grt �a��H��I05�Z"+d�1jA���N�j4������ 6���DN�B>�,�O܍*$���)�iԏN$����p8핬V�FM���,C��8��v�!r�z�(0
�@!U����ZD�2>�����s"#��f�_'Dt�� ,��V题�ps�1٘��B�Ut��v8)�������T�S?FQ#�N�6vz����cTB
��*m����d[�>Kq�.e8?&YWM3��sd!�!���@v�P���pW��)������a�ShQ-D�Td�v,&���`lE���Q�*������ 7�(��L�͏&ĀF�qja�
4��4\�Uȸtwn{;Y��E���|RGd�Zm���)Enm��t4�$�gEc"X�1�ڰK���n-~8�,)���l�̩gNd��Be��p��/����z��z��fLG.��b� ��(�d���Cഢ�#M�W[�� �4	v�0㛲�7
an]�e~4���KT�8՚�ʪ>�}0�C��S;f���rz�5 Z�BiJ�KY����ѭ)[r�*$�����s���F"5S�R��%�e!H��D�8��$NJQ��*0f)U��V�&�?k�H���e���o�t�*����sf�1N���
AR��H�\}M#��[�ު�\��L���N��r�����jtR��V�*��h��B�P��������4���c�r�VQb�U4"DVh�'=f�EK���F`UL�aP:&"�F������S�y
,�~ĩ �@~�3�����1�r�-J<Y��4������Zڱ��]&��1�hi�ӄp�S���\12S�aR�J�6c����6F�KķXJOJ�h8BLxR��\��GVH�{ prK7J���DVN�T�h���O4<p��a�G\b�7��t©y�n�i���;R��=Y
2-M!��(��R)�B�B�~])7Y��#e�0��Q�1uM�18�������ge!9t*��i|���B7-�2��p~���5��9�[Ҫ�����})T�ݢ��ځ���tf���YLW$B:)v�0i��0�[]xcMR��pV�pcӹ SE
�@���F"+pw�#�q����X�h��h���,��M��b��m��r�ZE:B�BMA�����09SH��&��d	�*�-�&������(��\>:"�~�Jp�D jA��#���{��mE�� ���'B�Jaj��cr��©\R��ȳ�R�7I��R7���S>�g�^�D!4YW*B�'A�������Ei2:��ϧV� 1M᪘�@~�F�Z�U7	>G���{�8�
"�UWX8p�66P�bJU�	���D(�6�B��P.�M�r)��DR��L�Tjsҙg��0j@��mhZ?�o���K!�v�����zĔ��|c?L�� B<�,ReM�h�b�ķ���R���|d>q�)C�^�p���[����h:�6�T�V�k���W���t���7�!�mۻ{q���}W�pߩ��#�\���d�}�?x����O �><~qs�x��;c�����_��@J���U�5��N'@��>�)��y��~��������!� ̓�=|�$N��X5�:���r�A��D�*tL)��-yۼƼ'��qp��H�/���^�sӡ�hE�pG3]#�V��z��k�BH��mQ���:}�U�4�W�Ϟ���~/.>��OI�\�,��ѱS����S����)��
x��jd9�|%�0�����`*�a4�d���N�!+�)�kd[�֒�)�Z������'���]�����'Ď�bҘz��
��:��P����ƁK���8LI�o]�w�Õ�������G�J-Ć�������h�ݞ{�(�⾐�k�ͥ9|��ɩ�	��Ɵm\�i�tn_e��9�Vu}���[
S��e��������p$v�dɮ�������b�V4'7�!:j����E��ݬv_3�����Ǻ ���w���Q��]-4ש���S��V�g=[���+Y��z�@S�Ns$��D/.�|��=?�6���M�Y��w������_��=~z��+������/>�������������O�N������[�_~��'6����\��ir�z���_O]w�K�_�^��1�{��_��޶�^9����=8ٿ���+{�_�c���/^{�t��~����y�����~Ή�|݄@�v���vK��Y�wf\Y�t0�PC6ʲ��Xj��j��'�)_9f	2H�~B���"0:4)�U��I0\W8R8���g�vM�B7�r ����(�fm�F��7�n)����FWՂ����m���U9�?^3�N���lr[�&!Y�*�U碭7��TiߦYk4�sY�ů�RZ,��z5�a�v�=cC�1�}PW]#u)#X���w��#*�t��)��?)���1q��8��_
D�j�,��2��|���	BL���4ӡ)dJ_
��Mh��$'�ʥI��I�׌�T�B��ٸkr)FdG�Ԙ*F���8!�"|�E��)�Y�g��Z�p8��19��n=EPB���C4�##e8Rj`��S�t�!;��4��4%�.���"s�>���5����1m9�oА�Z�9���# 1eM9D�X����s)]�V��9LԴ��!�u�%�2W<ec]Mo�85f��FSF��6�/x��fS�b��Y 	��|N%
M-
B5_-!�4_(�ǔ!�ģy�Ou`���ax4r���L�r�
k��m�f*e���$b6�קQ�5J�#�1e��rD9Ԙ$���B���!�QH:�9��"�d1�j����N��^C��0)�$��6���䶥H���=HYv�Co]� '_8��-�*�Ԗ����R8z��ٜ�F�,~�VzHQ f��9UO���>SPqȣ���}3e$��(�!�gd��m)4�g8���[����J�P#�Bk�f���5jo:5K�+�"bӚEk��R���5�ڵ=�����}]����9��u���;\�M�E�FUt���O��
��螠yL�o��N -i��(8i�V���e1�[��[��9%5�<�Sa'd$f�qJ]$�K�HrV�|���s�.�4kY���S�6�\[�>��J����s!��9=u��q���8��A��<&�U���L]�f�B�+���b�Q���Xܠ^Z&f#Q1=��IGݢPT� ����A6�귒Xj��&��㍖UQ���?�:�"K�Ď�l���Ξ�l�U�O�MI�?l��&����b��x�J�/��z�ȓ.��"F^��aJU�ii � L��`�K�֒q�f_gޙ��r1{�����B7ޢ���l��@�ͭ�x��h_�}����@�1��A47~_��_�w���fk��9� 룩A� �d�J��.�	�n�O�"~�3#�������w1�'?6���L	�F��i�2�����K��Qibps�]���2;}hӠ�� _���w��� �$��)i���o����_]���c��S����u<�x���e�)U/��-,���:�i��=[:m�Q��yF��,�,|S3|u�A�/�"J�:��b�p�F���
ᑁR|���p6�^I�)�l��b��z�i����Oz��/�I2v�
ц��ł����&�XVaG�*�8��ؖ4����O]ZW˺�R�;����M�
��1�Q��Ѥ�:��:�燷7�qT�m2	���**.8�L��qv�F3�����Z���G ���z�����b*d�U���|d2��{��i��F��O6�I��Q$��_��a�ط���9�2	9ɯO�Wn��d�_�jdu�!�&$<����Z�=����&b��?�	�W��Ͽ51M
��1ቑ�u�s!:[;^ear?�'����9,^�C�>�mt���q)�����),<=|{U@]���)��6��z�uU����h����>��"e�hw������kwK�oQ
'��r>q��Z�ӗOf>���}LuBm �A�q�~�y�fscm
*�&�C��ܡ��������ό�ƽO|u�F�?�O���8���:&q)_[-���=�Z��+?�̵8�p��s�r0=,���,3Z?�*~����1E�U�~��bըTS~��`/��R~��R��L��������p5!
�����?��"e�*ߪG<���^gw˛fFA�EB:M�+#N A%Eӵ�r�/VH�#u��f;�!vА�&o��#���:�Z����[v�T�1�u�����U\��
�Go>���^)��#�s喝#�s�^��:զ��qI�����pS��8��.l���+�0�������o�BڃX؁�����G�m�,��{&����ˁ���6��fb~��U@K]'�f�OE�
��ϰl%\�q|�Q��%�`��F����W�������Kr����	���?�>�c�nK�>�L��tt3�a�C���}9^�j;OS��|y���y%��&�?�ǫ��k�F�r��ꐦ��VG����Õ'��7:TN6w���w_�E�Y�v��ut���Q�}���)�Knl�;8����࿙+!fW%	+U��z<�Ѥ�ə���W/𥭽�Ǝ3�-FV��mLD�M�£��(F���Ŋ�[d��2@X��$"���ck���laulTb�FOξ|��$B@I-���o{^�th�4O%��DA�)���+4�8��u
��-�<�� �K���K.%�4K��]�>i�Sk)0ָ1�p��Ğ4�� ��	�ʩ$�%��h�I�jm�Nh1��d1���jK@�v�߅iDTu��VY`k��(�·ؠۦ��F�i�ax���hĊ
��^��)�Q_���G�Q��(4���&�5����͟�����ۖ��p��p4�j�u+�:��ˈ��9ה�R�t� ������+�~@fǩ7�����A֘��U
��Ն|��\����ܨ���4u ZJolr�͞<E���EQ߉�YT�)�;��L5:SLjV���=(�X�;!Ë�&�2�����6,aIM��﯋MN�e�oY}1,�#��я���oKAyoT3Q2��C8Bkl�pEo���&�-�p��5~Ė����BW��ĘS�+W+�������m�4/k ��h<v�~�Q'�=}{,�Á���1�S'Gv?��f้�A]^��@:͓�]x��$�0����--�)y�,Ϛ�=&	�e�:L�lBp<N��~1w��~�˱����3����х/��(U��?{��ѓ��5R2��� b
�T����m����((Fưewڕ��ފΓ�>��ԭ
�8!$�)������klG�>̄R�Xq�Zo̻n����>O��|���=?�
��ݴ�u����w�-U��'���Vƍ�I�(#��,�f~؃Q��\i�^D���c��p{�*@�}-��g�a{�r�:�K�h�{˫)�A��8XPcjc��,��@�6��W�@
�	T�P��C�כ�1
�'�/'�`��>[ڐ�S���K~�|��˃��Q���e^���A%ԙ1����&-����ޓ�CK��e��>����oǤd�)���\?�X-rI�[}k�����!�$�3�-=@�B�+T�K(��2�)5�t&��`�����'��\W4E��7���{��Ɖh�9�x"NF@��v�@E֑bm��މf��X��( �rP���~@�����}�5}pk���D�!U���* _pW�b�aͽ��F-�ԗ�Q���Y��a�}y2kww�i�����hMj;9bN	wD�G-��ԓ�(8��ҽ <?����؉(����8f=���]�zi\���	���9iЛ�CXnbԧ]Yn�~���X�h������gJ�û7A~1!��8�;�gݴ��H ��p~�5{��R��H*D(��)�<�G��҅�<N���F�r2Ⱦ�M�S��vv�8Ŭ��UI-H�E�V�8hE7��ݧo��JQզ?7���L���z�VXכ�y:��p�hhu�������!� 3�����2ma"��D�M�t4g�O�P�8�}�LTf��
H�q���Y �45�,���o�xb������е�{��]iU�iv��%���{��Xq���8���?�`쟸�jn(���x�6�!WPY_|�L*���' �����W)�ԓW M�|u�_lKt͜(�?{w%�9����$aD���@��8��S�@�߉]�������-�tsF�+ّ�Sw*����J����ɜ��v�}�\�規$ѹR��_a�Q\l|
��ä���d&t��"̜o�zT��)�Ʌ�Y���R��fCDyyV�I��G��3��|
��{ݲFl�t����BSY?���n���UFTo���}��E�s������ũ˫������''�1>7�2O.~�No�����TL�5�M�sK�7�:�y�%{��?�wz]��U���<�{��!^�S����6zr[���t��Qfs|��;���Q�kջi2�o�	2�b�g�y\B7�H�i���/�b��.#ö�����jf�k��y�d��ӯ���k�/a���4��G�R��մ���������|�ٱ~��	�^�}䜾#������3Mi������)�a��mA��B�J��G�M�zn�^��'�!}Ɉ�d��6��W�v�zDE���A<3��j:�)�.5L y2�g',��H�Ҝ^�4Uy�g�Z����z�����>�`d����;���Ʀ1[�GA��V��@���������ˆ2������{}-v��7O�R�OF�Y��l([�|�"�j��Ly�n������#�q� ғ�������4R1�/ލ�����:���'!�����!a��g����_������s����m�?x4�Y�|߰ _�b�	y��M���H�ݿk7�\\߼9���ƿ�}��U(Z�)�10n���DQWe��"��8.��@�h%��v���-������y�cF���0DlQT�.����>H@	 �V���\����>�MO��GW"wX�ߪ�����q�iug��c����\I�\�<�@˷A\[�m	�b�4ދ� Q ��,�c������~�E-{lP�"�J˞׺�yK '��p
@��e{p39����T7�d�����w�ow�E�JLj�T�[�~���۵���,7S_<$�RŬ!_7��^\E�7�+x�4��GO�������;��@ �(4X�kS<1S}VL���KS�sLP65�����Sβ5+�߲��{̨֟��,qc��V�mLg�s���Դ��?_�:��:�+ݑ)�DWe�@��[���m�L͏�W*�lL���VϭP+qvrBt
鄺ȣ� �d#��(��Z�w�Kx�W!�ZI��X�{δ�婖_�ӵ��	>Bӵd�?#����X�鵀�����vĨy�
A,��-O�E)>ݔz8�h��- )��@�ИR 0�C9����T3"qqn�����+�:�
D]1�(�u"��. ��|<BL&�>�M��&��$��ص��H8����oO>W�;-=>�UԻWY�j(̰f^!�(�4lm3r��3)�њx�m��.O����A�IJ�olc_�&[��p��wqז�Ž���}K/��Վ��秇��{��ܱ�w{��p8[cfj��H!�es��Zd���	�!/M3D�W�̉������(���� ���
o��y(lw�Y�Ge�[��%Tz�JH"�����e��#~�t�P�L���a���X3ً�4mr�{Wة�%��@+�������?-�[����*y�؅�N��'ڕ�[m�� ��i�"?`���AVh��k�;
;���?H��2���[�(������X�B\�a�A�nJ��J���1i�쌅�Jd��7c���"F꧞�K��)ݢ���'�?t��|����������/:��,�V���'�Ng숡@+la�0P��[pf�$�[����y���
���S!���|���W_b�N�G�6 ����J�Nx�"�)�	7o����}Qy ���ʳ��-��܃O0���>Cu��;�DD���!�]fsZ���M�Bd�o�����B�܉7���4d'c⤹���N4�h̉�"��\ú��
r3����E�g��3�f'��mΧ��>�X��v)}�c>�]���B�������uMٶ\+��@�|o���u<w����Cii��S�g�m����Y�i/�}�~&߽�h)p������^�͈�y�����hD
�����r��{�[�ȹ0.1�?m�ld�[���B[�$7�ܾ�Pq��FM-��D�k�T#S6����;�r�|�[�z&�K%�{�~_����")F#i���C-�\޶�'��}���u@�7(ID���oy�u��U J����^F
L���K�ЫVV���e�R��f*������AtC��bs[�c�5�X���m���+��
��N G�%�h��{�iJx7������]���i)���j���u`y�=�Z~ ���t_όU������$��k�a �۾�x����id7�H[WI�6��)���y� f�>m͸_v�_ �凙���j����2y��׼�J �Y������dfQ��������q�
w�.�~��"�9� ΝըTgSJ?��85y��`���|L`��ߧ������3�;.�g<k�;�C}&�����'����^C����J~7�qT
����?�_|/VF��j��R," ���_>�^J�Y;*��X��:�5�Q<?�2�6�S����Rl{�^"����Ұ�6�X�p����CkAʸ���;p+P�TȨc���!c�������-p\�/��O�$���A�0��o�N�n�ma�P�j����@m�b��#����WWkC�Q%ro>��^m-\�M
�v3�;�_΍�ω]�X1wv���s���bУ������S.l�lJ<�)ۣ4�*O����c�@�^I1(��7s9���k�*�����r�}��y��y!!k���e��ih��96�z�����-��٫n6��˚Yۭ'n$uC>�!,�[�g@��|���[7{���.k*�ȗ}�i�<������+S�$)_(#��L�Dt�In���c�k�j'�;����Z��:�����N=��}t�T�j܌�z�S��O�A��U���Ka���A��bݮ�rp���E��������?��
枞��خ'�������U�SH7�o��W�j��9����|NЛm��6��`����Hb�G�r&���:�O��Hr8Ǌ��E-������"��Y���@R{2�a�k���W�8ߌG<I�=u�h~}��7U)���T�,t�(�c�)��G���s.֠ 㨩n��e�l��K�U��i����{�������|x)�f,y"7��8�c;��Ф�Ս�+�Z $�F���[��Tw3E>��EI�C�q϶-��5o[��:JQxx����'��:|�z�I�Pߍ��Є�R���c�WǞ�<�`9��ǔъ��Jv#�d����j�S�j�]��X��qv��4���Ow�3�C��Hal�:mQ�:D�'�����ؘp_p�;r��5���U_��3�l���4j�3�Z�e�V�1�H��R"�E�O+��W%@���t^b�'�������O!+��^�w���qB*�|�T��J�0E���;jz]����R������<�g0 C�/�F7P���EgPѹ�)���
��Fл�-��Q��݊ons�H�MF`"���ة!�9sytKj6'/~v,�[m�������k0�}��6�\a�����P�Λ���gK���B,�	z���G�4�0s�B�%r���eY����F��Go��ͽ�ʯU^�6l�&V�q�:��擧pI�t Ù?�1�%�ݒ5��֜�Js���y����O�w�x�>�,��*0���{����?�p!�d�sO����/���l�:�����T�<4=��/����N���ߕ�c��
� ����$�)5�m���m~m���oz���qm��f�{��<�3���;b�L�{���<7�%�J����x���gs�R�G}��L�-��O�(�磄��ِ�;K��#�Vmm5QZ2���[�!q��l��ù�����%`Q�
 �\v�	�5�Ϋ�Uz<w���}����`j�|�ҕ鉶���N�����yt�i�Ff� �Yr2�D(�Hp)Ir<ߐV��2^�W�.��I�ڇ�?�����j)�/3�P�K�<�|�v��/�}"�)�VH/�*:�v���#�[va���׳*x/� vADc�a2��{�����{��p$����X�d���[ϯj�:�x�`�Kץ�����@As,����)������PM(�����I���� 2 O`���f(%-�P�/)d�*>"���`�@��ْA	�M�0k��X���
��Jƴs��$�B�(q��r�Ox�AE~��'��NA���+?��X=��������S����[Z��E��~���Z�Yz#��Iד��؏͎�����6�P$h����<�ב@��
Q���Y��U0%��>;�sBsP�.u9���6�q�{�ʘ��\�9xǧi@�g�\�����a�͊�%��K -����wGd<��L6*f���IO�*�[^>����J��:0��)�B����how%x�Q�C�R0��m_�ѯ�>�UR\��[ʛ��Ҩ����(�=�x�����WR�;�_�Cx�T3U�4WT�t��Mҏ�Y]o�F��X_aXU.��b�f�-("�R̋�;A�<2#�s��s�[��,2�Ko��xR����y��L��k��ߥ,�C���[{�ǫ�[��u�b�.n��GU�x��T�q&�\�y�+n���'�V���p7py ʂ����� �Վ�B��)�b�P/����V׶�6���5�q������g��2-.��I6:Q��qq�Q�E/���i�Xr�9fدZKy��S-֫�V�z��� H����62p�{������7���q�{م�		3rs�r?�e���W�����6���3���E���#���d�	Ō���b'9���1l:B�U3��}��!�X��j����l%�u!�i�����u�θ�wL����rD�3V���y��M;v�Oa�d�����sٝ'k����o�t�g����Bk���e¯Ɩk2���/����\�����X)�ኯ¸�v��k�^\	�t�`dm��$�Q�μ����t���rW�?S�@�1l9Qii�����h�y�f�V�`��0;�%�҃h�j�"޼[���1Sr�
��`7��MkZ/)�	9K[V���PGH_��]/v�.�����n^��3��:�ޙ��J%�#6z�y��\��:���B�tKS}q�r.�S�oٶ���>�{'N[4S��
;/���?_���?:��Y{��������/x�m%�Hݾ�w���R��0�n��r}J�v�N0k	�S(;{�wu}sBS)�����Q<�\��*�No~v�Z��iu���>��._��T�E�}����7[h�(�
oU�V��}'
�H�G��^�����O��ȏ*$�pT�
恰��,�iy��L��ӂχ���͈�)��y���pV)gx*Vފ�2k�S���$?�/���s�E��ʻ�j��Ժk ~���%[Y^4W+}F}��o��^�������,�����ak�tۂ�1bɞ���t��ga�,�xH6�����P���׺Y�
2��ִQ���w�7�0�%�sD�� `_TO*��H�
BT��E=��Q��W��e �x�o����N^�1<�;��UA�4,����P�4�u�ةf`�5��M�����y���2�恳����rPf�)_����kj<��s�i����`uKS>�e������f'�cz`]5���R-�v��j��iƚ��Tdnc�����M#ۓ]�������s�_��\a]Dp ~����IƠ��7�^�2~,�L6������ag�*�*���Rٰ���I�i���10\^�Gg�!T@�ڧ[8>��q#�݇B��Y�G����U��$`CA�Ò@�aW
�Eb�;h
H���'ޔe&[�����#,;��z�{8�]��0{� ��nS�cL0tO��Պ�M�r<	�����\wB����J;�"�ghP+bB���f��t���:�gA���P���P	n���r�_�*�	ѧ�%/v�����4v�F����R����7���-�M�����E��Nh�@��O�p`�kO\dۗ�0�s��[�D]��Ǿ�3��u�um�n�H;�V��*���%;��
u�x�	W�mʉ��͇�������;�`���-J��܌�D�%���f��1������a��7��Cv^E�MP��`i���G�����y03z1~�"��u&8�/�����6��	Z�Y�\�����,���;�SS����E@��?�C�.��l;�s�>E#⬋��s�����ܦR�R�{����%�i%�"2S�Ym>���^�O`G�B���k�3��d.N|N��-+�K�w�l�j��
�
?_z����2sg�i��V��n�E�_(���ZF�t�a61���d���9B���wjэ�.K��b�Tz��cӪr�qW�������iV K#���}y�n������Ooy{�>S5�w�uyo���ې�)S�F`n�&d\!�>��c�x�R0�W�#	��+��av-o9e��^�[�8Պ̮U���~S(�^ߝ�Q��vQ̓RHΝ@Ϯ��%�������D/�hG�R����e|������
�i�_.���c'��P�Ҍ� ��x�&p5T��M�����j��į���]�09=Ntk�ҟ ��Zm���c���k�HC�����&���[,���W�����46��y� �)
���:��i��[�H |�+`�'�x{\�h]��T��1���oF�|�� g�ZA	�=��e���k(1��̦+���{�HZ�VX��!]|�V%��q���r铢��g1���nS���+� B�����Fѽ�Q��ǿ�=�[ܭZ/��/�KV/`6w��g��-��Q�����7�X3��jrn;��)��h�ҥ�����'MyՎy�7�SV���}SE���� � �z����Y�7�
B�L�п{>����F
��M�g9��B��M#
�L�g@TІ��y @N�ۈ,���]oFU����Y��8h��XQJ�O�$DOY�4,����۩��F.��(In����!E�s�q�yiaɥ��������ے��*�G�d�Bh��q�~v'ƛq����e,��������o=+%i 
��d��
��u��p�&h����+��F�W����
aW���z+�3����mn�:�%�ut��M��~x�x�øR�;bB��	���@2��Ǔ		M�)��:|��-&?$ͺ_Z|�6��x�zk����qg�:���ց;-�5��J�a;�s:��o0���H&N���U}��n�����ѯ����+���GӼ��Lދ�F	>����|��Sw�B���7���e��OQ#��3��A�g$Dx���%S�]�5s��oJ��d���H��ٹ�^� D��`�.Ha^�Hk��<Zq�j	��'aֻ�c#;';Cw�Wf`๾v�>���˗�׃.�[64�����_�Bo�~��i�^QV;��R�Z�P9�#sП�Qs��v��o��z/��:����z��#�xq�xgs��2�_������Z}��^�����_���/_q1T���[�-4jk�����$8z����������d^����ٝ$�?�-ļ^-���y��P��tR%�NA5��;�;#�Ki�>7�A8~�bI�ӵ�={}��-$l�o�v�t&����cj_S��Az\�޺1Ȩv���"�ɘ��-�Qd9p��d�����C���� �f�xQ!S������J%�ͼ\4��� �[3�r��4j�b�Ƀ�6�<�-5���X	��ԣ�����NTʹj`�k��?"SV*�}r���L�o��op$Y�c�Rw�۷P%>I��Y \���p�7`�m'=Ґll�N�$�|C�f���e�B)���䜍��W�n/Gs�$m�yc}�&o�4V�l�7H�*���T���_�'�ƥ��y�u@ɐ��b���(���6�OaQ�[ 8����Ē	�℘�Ey	����
�mӂ[���$0���j���ftTF�%ۚ��ͥH+%� �����c��8v�mt=��G�/oc(�0�b2*m/8$�(�&!u酌Y��(�0�8$��&�e�D�
_�xO���0��hS�����X�8X����)$76Pe|�ƳIZ5�$<�g ����P�z��Tn`�l�����T��͵�b�Mdj�#,��ߞ._����d�Ao�J�G���q-��3���֧��Ϣ�J~�j$�L	49��T��Nz`��w��0���%��m�%���ɓ�C�
cbHc[`��]]�D@��2��4 +�T�j����U�r�[5XbK��۵8�h��6E�:�G�j�[�FǻW���0�Q*��q���Z�f⊘`��"0�H5���7��"�r4@%�����'o!ߡ���[�X�o4$J�h;�q�~mk�5���/ᶠD��̕��P���jG�KN��x\er)f|Q����(#��yu��Eb��w3���x���7rE���WۖFE��T���$!����Dm=W�z��F��m�Ŧ�!C���:�{Z:��U���Q�IN�P�:�-�+=��l�qƼ�TC�|�m�8�
��aN[�!�I;.ā�y�����q�Wc�-p����à�]°�'�$�ް'�����m�|�5z��ֈ;>��t��Ϳ�fr$g �y�)�T2�m`��u"��*��|�f�+\W0��wj�7��:>C��6��Q���S�e��C�sZrg$�X\�����KkRM|�|��4�q]��t����Zzkj�4ݚ���a���o��߅������[�,3:��Q�"E�05Xf��x��z]a#Dd���]�BoO��Q��j�����\T/&n�^�D�+���T]��0nQ��\���$׀,="����%����"��Pl�&����)��N�[�#EVX�����o�Zg�;�P 4v���;>����
�u�q����2"�T;IaN�T'�5S1�wȓ�>T�l�(�5÷O��uYz�@^�̟m�:�z��䴷��y�x�D�o0C̒N��SҔw9�qh�Sk�/RC��O�zҗO��Zy6���z4/�՞bSU��-dđ��W��-Ŀ��8�b��Ѵ
��Qm4v�sF�{V�d��"�!�QV=������ǲ �����w��Nf�U2�^!�gN4���W�sݤ_K����uʧ���|�N=ⷤuB�+/��/i�Jn���~ޥV�bƪ�A��>wάRB�~���c7(�k|������%��l�Gt�pS��N��ゐ��.�h��7�h
�&{�_U	�W�«A[y��r�����q��t;�a~������~���l�h��{�uhV��չ�WB���E�KYU������Ѻ!ÇRMef͇�kW�/��^�^<^��{q2��ѐ����K����������W�H��^��Zu�0��;�*S�{�r��R��f�Z��
`�@�����z.͓���@G����2O��'`�j�lLHfm)��-�`����M.���]�Ӧ土��G����13Q;e��Ï�&����\���W=4��e���K��^zX�ْݲ�4�&�m+������2�����#�\'Z��~͏N�T	���B>�lUo�-d{�y�b}�����'ޤH�mY-��v}��P񶷸A�Fo��i#M��4��{���}��eV4z=}Z<l�&v�VJ��b�/���zȣ�����ہA<��DD+ɍ�䪛�Z��qn@箢,�B=zz�����1�����bɼ$f����l�je���친��ƫ|�7�·��W��ھ�lh�u�+�.�B��}�'�}��C��x{��wo��j�0�����b�G}.�Ң�q�ڶp|N����_�K���I��p�G
�?��q���k�aq�m��(5�����|J�Ǿ�ڜך'y.�k$�a�~�"z4��c�c��5`:-�K���R{��Ӊ�����b2r�53f�<�o:B���"�n���yJ��1���S9�!�Uz\��Aa_�J�E�U;�sm���Ӷ�U��}����{ �	�r�z�R_Za���YGg<�x����=��wC����w��
V��A����~�l�gV����;�:���6h�9v��L����X�m7)�.,�>�mY"Tr���K={�7�dx:M�B��y�*}C�+����C�-{��?�X!�˻�ǁ!$o�r��Wz��2�U�S���(U��w�`f��@X$� K����b��|������P�I4v���>�#�賹[����#dܠ���,S�Jx�ׅ%��>e�c|��?����IC�!]�����=�X1҅Sㆋ:�F�����rJ��+zT,tep�� 34������zqE�e��r
�^G�\��Z��Q2g�&�BE��X�`ۓ#�^\[&;
ŜLWYA����7��o��^r�v���E%L�a�t"Q����Pk҃_���T��, �3>wp��W�ϹP#��0�I�3�2������A�H-w���훞	U�=2��;�+�S7��LR��d*&-b���z�T�!��P)k���7+����4�:5֡,5�Z1�	�I�o
=y�z]�E�F%��=��y	HE�&�����ciJ/
��6Yw&^MW�7�3޾�d���� �e����e`,�ʰ�}�i��$G���g��J���Kև@,.K�zD���3�̘�[�u�C��62��"=��8��K�,-f$o�`�L4��i�҃|��a�D{SA4�u���2�� N]��vn� �c�3���T�f�"8(�pD��Q��\Mr
�߫H��!�ś>��z��?l8f��^*��������{�قK�l��T_r$��<��:�ѽ���?�䖤�7ƭ���H]��n�H4���1�a�y�x���;�j�C�c��ߌ�:W�"w9苿�о��ӛ+�H��,�p�._�*��O#�.�/�2e}nU �i��W!8\B*�|�3.��P��w��yG_�����h�o��~f����*���A8"�{!8}u�E&!�2Z���,���)�5�ݯ8��
����5 Jm\������X ���&���.�@Sbx�/o�Y�[7�0T�p$��6V&��S?�.�X��v�9�W�N<qjT!�v�ˣA$�	wB��$��q�mJ���˨j�:�(����x�7w��G�"L �Y���G���iDEt�S9���H:т6)��p�����8njq3��p/�S-�Z.(dPv�9$�9Y$�9��B�,�Ss>�I?�L�-�W��Ѷ.wm����5�4��T�M��p������N��	.ӑ�Gfi�^������10��s2��&N2�u�M�a�Ƣ����GjكƉ�ztT�4Z�E��KGQ}��̛A�C��>��`P��o��&�G&�J�ҟb$o��_B���ɡ�S�p��k}%���ӫ�!QvT�Mw��޶Ek�b�(k�{4�&��;"8	β������i�X��imcwҞ�y"�t}�z}�'c!4�o����Z����ک�����E$;g?p�ϳL8��q�l.5C�$�>�Z'�K����3����CJE�2.?$J�oY���w����HZt�j�M�f�6��/CpӜ�{S�a[��欸,.�!���v�)a4��W=Q+{/��PT�|1#|q�]�^��Yh��j�%��CG�vky}�/�`�����&`M�B��L�Ln�t��|Ӵj�Q��5=��$�����F�)�~����ib�)��bav���D_���Y�X�,�E��~G��hr|��T�ʶ�,�ͩ���?�|�|&Λ] �W�V��ջM�:_�c�wq�� �>����r��Ǘ���\N�����W��\s��8��w�].����_�s���GyB�=��`4�s�Us�������}��FC�~��vv�n�,����x>��8�n�mM��]��]Q��;RDW~Z�#5Z�^A��N���3�9���V��v��f��j������;|��ѣr�F'���p˱me%���t����E��(�a�a�KpB4��pA\"�H��n7�	)Kj��Kz���bH��M�̧֎Fd!6��_����΃˅������.ٞ��q?��|��_D������rC�ܮ�����?/E����r�>j�̑�Ʀvlg�̮�9�
���y���D��sG!淯'��"d�L���j�X�P2�fƚ�~�X����"�[�8>�}Q��q�|�#����Ѱ�����?���u����m1��g�,��v�9`����6�GCsv��E��+(1D��{M���4CI�D���zFm��64<ΐ�j�rj$�ą�w5�?T�7�ݨ T<-T9A	���ϕ~rR��ފ���3�8Z�KwN�T_\!����	�(N����"��vWw�h%�rjpɐGk��!�x����o���]
w��$�m���D�y�l����!I�-R�w��VkC���Vz�O�3�8S��S�X�z��|`9@�7� ��~G��9���H��#�|�EE�W<��:�s�1�]�w��	;���ߣo��U�J=�1�^�踰�DP���QE��K�r5lG�n�L_���f[R���ͧV��K�#7$G�c<x-�ڋ��IB�]��1�LR�X�f09�q��`�;�=$��)#���'3��ܨQ�_�[�{A�V�2��H���R.L���z�2�SA�5����3�_��a�%)�^�eߢ�2/B| gv=�}�P��w�+�
F0*u�uǽ�$�����&T�D3�@��;@��U¶�����3qv�|,z�f�%L6��u��ЮU���z�k��ؤӰ�q��{�?�׮m�wq���r�.�_�~-�`�	�5�/� W@����񅌙���ë�)jJ�o��]r͇ 4�[-�YE��� Ќ�@�5�3�BHI�E�'�Ɋ�K�D�Mf�p[~H
r���]e��4�o��)7���M����\ӑ��Z�KI�_H�#�H�3���	��Jpd۷R�E���3-������f��\��6!5QL�Ϯr
%H�Φz�D��3��xR�GT�(T�TJ��ń{�� ��ҦF4`)d%�ƙ�VN"�-͇�X��iO��I�XncL`
ƚIs��E��
MJ��JA�nрDi99m��r��cR2�t"*276�h����舔��%�SJ�aS��l��)!r]	)7[�>[Z��r��O���Ց���n*ϣ�6ߴ~�#�+�j��D���^�Y�zS���"��?�ZZ�MG�$�G�O�eb6��h�~ cB�!� !�f��!WEt�ѩ�0N
4%�-��2S�c�]����w���J��4!���"�[�I���I��V�n�M�8�i�Ä��f��W�s�J�%;���iE��bJ?X?�@�b�i�PȔ���r�	!�\���J�&K��ȴ��p�
�*�l�T�?�'JΪ�n/TW�B=��D�OvV�D��׭�t�U)�H��sv�w�������_��D(j!qD1����N>Z�q��ص��EY��$�K���\э��9F��̇�@�r'�����;�&���bR��Xj:�9���|�d`��o���>˚[+e�\���?͠��-S�Ԩ.�\Q� �Wi"�����(1�B|����l��._��%%�1U�mŴ!�s�q@�*��1SRq��L-x|>�����ݻB
\�&�v���t.�i�P+a!5��F�ũs~� J�REK�'��R ��J�:�Ɖ`���1����IST�I���dM	�(7m�c��p�݁w�})灃������3o�����>Դ�R��do�)s{�/o�>��u�ig�톳��ѭ[(q�8��0w�#4��u>��cN-���4���9��� �������?����5)z�Bʞt�ҭnCT��?�#�R��>����CgCJ���m����^��S$u�g+�����Nv��:O�@�49z��9�:р�v�ɨ��(0O�g�l��X����}��`}߬�}�ҧ�^�/��?���z���뫣�ӓG���ή��=���u;TY���߭����R�1\u������ ��Q���j=��h8��E�CX���1�2�.���hF�~A�Q>(h��.���۷��H�9Z�/��2���F5���4"�v�5( ʀ8��}Rͻ��7�9}z�h��;G����l��ܕ�Eċ��z,��Ub���7]ga-�o3u �^k��<0w�/?��ٗ��?]uc�(�w�R.�E�u,��nk���khG�1��5�r��Q!kw:�׉��=�L�3`C=6��e�)��j'e������Z�\w�,��n}����Qc���M�3Iʵ����uv�bK��	Bt��Y�iY]E���y�ץ��[��>��CA\��xA]RJ ub�Ԍsb�����>����ɩ�xs��'��_������ܿ�_��O
kc]&��9�|D�s���̛s��>��8���`�zr�o��OONo�n�O�N?:�:{���E����)^�]��,Y�ͷ����%�Y[!�7�Z�ɧ�U#[���FZ�)J�2�Z%&�;V���^��-�b��Q�.�۠rc���BB�S�*2�pF����q3�|��@>�x����*BMj&���UKX(5�9R4�7R�(����:�������Dl�YV�R�d� ��=�������jI3��&B�,9٦BLu4Fy6�SHĔar\9�>�B�[�u�Дc��a�ҏ��MY��=�:h��|:���T�Q���:�8m��7����+j�@�<Y��B��R�����0�r)�!W����%�ZƖ)�iO��pY��#����s��D(�`k,
y���V:�B�s�OL����`:��BZN�.�\8�D�e2)�t��F4��%�[/�t����rk�����9��,7�\n�-�Z��_zR�q�bm���8�qJ����y��?�L[�VcVTQQ4~�����r���Č��o���/+Y�6�%:�է�8��?M)|l3E��x4#sQj["�����8�P�R��V��KO�Vlk|k����#T�m�凫��B�HW�S��2�)�z!�C��1~S4)����,���i����n+g����IRmBVu�z "$�ɯ�p��)�hd+E@�3D���p<��H�4Y+�%d�N�|��gö�II�\"��q�pJ��"@�ʵ@
�9�R�#�؞�dt,0?}"�QB�4�B�8r�Idw�d��D���ϩ��_]U�hYE	N.e"��M3��k�t�
&G������9����넃�,�m������D01���8�V�M� �Hu�r7�r��tt��N�@VKi���(ʩ:~�Jll��*�l��	�U���U�
)B�H	qʒI3҆�V�FY��Z#��|d�ǁ��	i c>\��)ݿΔR�Ɗ�G�Z�F��g`m�R�eJg�C?5E�r�8�;��I�\L��)k�j�*�O��V'5$�c�m )6��tL����}�N��N3�*����(WbW3A���B�4����{�O_��uዚ��I�:'"Et�J4����pK�H�|�����hM���Nx~���B�)JٴÍL����H'�1Y�(f�v��B����������F:����C8C�o���%5Ѳ���9���eь��Y��L�����j`@�@��)��q���k�V�o�o,%N"���A�������w����>
B!U���e��K7.�|w]8����Ū	�KGb�pS���
I�L�8��_�@p�Z�D9���d�%vQ��D�ȗe,Z���|j�h� �Ve�LM����Ъ%k
�oC�D��H-|��B���Ԥ��_�    IDATِ�@�1'�>p�p���t����At:	��?�L:��@�B�+�P#�ܘ�̺�J�����$%��қ*�̯I�J��Í��1&�f&X"?�5m�!��Ɣ�Cmm�k�Q?B�J�cL����0Ӫ@89q��Q�?�����[Ȯ��6J��`�R	Q|c�-�E��A�ºd)�U���H�i	��4F���n��.��qDM�,��C�J#�K$2� �!dC�K�P�KH�zᢶӭvy���?��i��������}I�������s}:��ko����7më��կ�u�C'����x�OK�Soq;�pk�Ļ�f��p��5�D��Mu]q�%ћ�>4�(��U"�����N�\G�����UQ��^C	9���ԶfT�)�NTG��R��Y�B-9?�!�����x�^Ѯ�����?������t*JS�D�V�h�+��uH�yp|��ӷ}~���c�W�/�z�ۣ�W{�{��n�Uӳ���s�]D�rHQ6�9m����o�9F4+��0�0� 1�(EmQ7	B4�Ȣ�AX�m]JS!KuL�������l��ho�	vo�AA�j�(�xhi-����X�nZ��VR��@TSO9q���w��O�^?:�G��N��z�<[�9��[��$���fϯ�>�	Y��Bg]��SO�����/p>�s��>�y������3�GW�Z�j����)t!Z��� P�n ~o� �nb��IJ�j�����x��@��F7�<�\&�S�]�>��8
�� �ɟ��c|������_�6�ow�_��_�$��|@���W9����/��/�.��o�����l	M��D6���Գy���V��U`~�;���?�s+u�a��IE������ɺ�nnO�>}�?}����ۿ���^S�8�w���ǵ7/�sq����������ՕO����W�?Y�=nx_HKS3릺�r�9]�ʿ���>}vs�M�]�6|u{}s���M�ѪD��R�(AS�芻@%�%l�i��D`"������!X:D�-NuG��	�����H
���\AS����Cz�n]��C��e�C#��F�;�
�qD���R\�]PØ���E��\�1�J2�!���6Sj|6���A�����&bl!����6����`�-�&c�ŀ]��M�~S|�W��'�S)��`W�{l����#W��*�pƈ��C�F)���9L'-�t��!U�Ë�o��,J�8�飥)1��G��$�%�X"�/+)�� "�4�h/&|�pʪ�#%�J#�|L��鞁С_i4d�Mh5��7�4AK'j��9�妫�f8-��o+��R���3�,���.�Y�V��Q��)`��O�DH� ݊ZER��pN"���)mO�h@
�fM��+�����<M!���hL��|�Kn[>B�&;8'Ĉ���m��!9���Tzt��X?E��'e>Z���O��#O$�����T!S�5F�T�_T�̢��>>N:i���A������3NRp��R��!�CJ1�U�Bh���-�B�	�2e"�Uu�0�꫹�J)F%�h�M�-�6���#��N"Ǒ� ��@jY=@�q�+�Q��BDL��u4�Pnmw3TBV:���	�k3�I\�|Ə��� �(�!�m���E'�EA�	��L6>0�{ �@�.zM��HU^k~�u�Y�iV��A�X�B��@)��I��#=G.�Ok��S�oJ��Q������7�5(�n�r��-'���Ia�^��"�q�ġ�m������i�!h) ���('Ŭ�i��P�rM"���J*��.��� �	N�!@њ��y��(�	a5�,Bd`d�cK֒P=h)DѤ�=��ф"���)#(=A`R�Up��b���ix��| CL%�W.n�����Ĉ��ќ��S��P
eY��t*m�d@F��E#��c̏`���S
q��1�@pd��'�����#Ԁ�#É gM�sD����yha�ұ�r��"sX����ơ��v8Y�4�3(D�S�Hx۞��B��)OV����(,����CAn�m����!���a�RK����r rmT���jR*����ĕ�K�p��J�M�Gz
E+� B Z5��҇�Dt^9�!N��5��[��@Q��N�JѲ���j�����R�&g����i*�ҳ��R�($r�@dQ�\S��B%�I	���(j,�����Y͸C L9mH��%U���A�׆����I�%"�5�̌�*T(�Q{m�P��i#ASu'1G�,�dG�ݖ��C�~�R���b�&*�*DYS�)�D�cZM��]��2B������*P`�	J1�a��)��t���!��`jBr�P��r�%āX2�*i��I�p��wk�0����ld�8r�ȕ�輢FU��gWD��b8�FR��V��/j$��a���RH4Pz�ܮR|j�-��6�"Q�p�6�BmT"�0r�ve�l]�X&B�_uS������Kz[2BM�r��F�c�}���P�(A�ˉ���EF�������������@H`Y�F�Z� �m�eE��NJ�G���V9�gd���,���G!$5>>fY8#(d�ԛ1r`ϯ~,��\守 2+��M��5��W�ݽ�[�@�2>G���ѣ���������7�}�������.���֞wYU�M�xl�\t��ћ㏵��3'8z�q���p:&t�����۹޳u>����g���x��zP�*̔�nIIl]�t�vL��Q�HG�΀\Go�׌B@
A�@�9m���>B����3�V{�5���o������|�sn����wp�@[�F�ۙ��~2�8j�r��?��t����]>;y���ԟ~��7�"�����`��s����m����5���U7�}�ԹE�rD�,��#��.����I�Qp�!KHJ;li��,��7��@˷�*z�޾���P�
5U���j@��J4)1��K�ߘo���E��O@^�P���Gv���/��ݣ�ŷKt�ɢ��}���;��U�?����=��}ݩE�y`>?wv�٩>��~���o������/�Հ��m�^�����Z��3eT0��|�h9���w'���=�����L��s�h[	bz�ܾ�"j��rX蓚��'���IqC�������MQ����{ۧ-!Ȋ��]?��N�pO���t=��X���zf�4�ڣ��p���8�[j��q�~��E힨��`V}j�����e�yM����������/���~�����ɞ�^��Y/��+�O�=<��Wׇ{�+�������u�.�W<����/�~uw{�Z�����g�{Ϟ����s?E�U���:=E�~����l�k�G�����M��Ժ���b1g
�b!@[��j7�V:44 ����AD��9R�����-\��d�p���~3��E��ҧ���t5]Jd �*����.Ad
.�p��n{j���N�/��@��߶@<Fk�޶(Ǒ>��_"$H[T�c�l�,��
Qh��)>�t�q�'��$�4S�l�z��^@m���t��=�6M߾���|�O��80����W�������om>2\u�X; �+ǉ����e�l��IDbd�h!4����pÛb"��)׀PO��\!��dAH�F�0w��P�ӌ�h�VMS:���g��(|W9)�u"�f�e�|#_�~k�U'B�S@�4!Ul���hJ
�S!�c`����/��8U�3����L�Ⱥ=$��ߪ� 4�����y#�G�[��V��!��)"� ]%�ʭ�۩4:���'ŀ�YN��G��XLU��FD(���D�6�"���@"YQ �cL�Θ�Jh,B�Bl���j����i���1���چ 0
�8u��0�s��)U1�j&B:�N˩�,4!��KA�3K�����A"p�˝DD# 9���)>��)�=#Z`QS�V����mK�2E��U�e#DDuLV��!FQ4N N� 2�0�Y��"�U��A\��+Gm�P�i#&�S�d���1�O���o�謦��F���q�B�@>��|���R9���1ۍ����7�"�1�!�L(����G�n��OR��r��TK��L.0g�\Wو�d�ܺE�Lw;,�X��փiUp�M������p��r����0| �'hZ��pZ{1G�IGȈH��!������z3�g)CV���C�t�)G�_)>�� �A�o��_ E�#��O�B� 貦�/k�rd�Rc)��F%��ِ��#T|Y#��Jk��]>�AJ�G��1&�)X����rg*�:f�����5��&�1J4�1JQ%�����m�
Q�K a1��vH����
�F����_�1�1�P��ٙ]���]�r�G��Z��y�6���'qk1�crL+��@+m,���@�B8�����?N��4�pd4=����A��j	h�
Q��� ���!�C9�|��D���j�0�H5� �5m!�E����S0e|c�8���P��3
m���)+}F:��jaJ�n�L{�0�ݵ�P�j��R62V�f�5劣�MT����!ފ�j�!�T���E�I�9r�&��Q���0j�!׹hL�(����p�2 $�i��P= 0"�.BӖf�0D'r�L�1>Z����"�cS!dYE9�P�t� 1M�>#��F �vN�L:��d ή��N�MM"|J�b��j�`BJBL���w���������I�S.�cZ�*��J'��ĩ�\S���b
L_�FS�W��"�N�҅(D02j^��*"S�O�hc��98Fj�R%Xcp�1�+��A|-d�j��q�\YZ26��ܔ��/�J��q Rc���W�N����@�����J�Fd��>(:|���YuL�1�G7�e�y�ܶ�\��E�!����O"��q��r*DN�X.�O3YL�_E�C��6����O�r�.MSQN�8�8�v@V"���,8Z������K9F�8C�io�kJ��t<>�!ǧg�m|�ə��Wj��F������~��˗>i�ެ1�����x�����*>4��@K�%#��� �{�ֱH�k�C��:.zS�۹K��鐮s����8p�w�k�[CFʹ��rF�U
��� �z�#d�L�y�����z���ȁ�r�>������..M�w�=�¬u�S��\��'����ٽ�tdf����͑�׻;��;���o:�[�o��C���i�f7BQKƹ�.fQ-�]��@LS?N�Q� ��]uq]�J�S�v�θ��{�t��}p��S���u{gU@+@��ldL�Ԗ���_��oƾj�_L<����j�y�\?��zt}ָ��ζ޿ .��5�럗P��(��\�3�W7�
~�W����;<{t�DW�_\Zޅ�"w���[�η��wܦ0��&:�p8�P�酳I��MDv��B�$k����u���]G�����vb;'q���sG���ڼ�%`!��BⴏbcCH����~~c��+K9�h��SO=Uc�1�^����6ʶ�
����_�9�f�y��h3]�?�P�5p�x�������z�J��e���>��5LV�;�����.j�>�+�I��\%� ������bN��6��a�r�ZZ�;)�1-��.��������'��i�+o~UW�~��;Gw��~�;��e_�_��zR�����`�'�W{G{Θu�����t�~�����{ē��?�/^�<;?�{�ҷs�4'�������v�uo[�+)sftű^��.i����NT3����j�W�Ƈ�""��P�d�E���G3-1�K�;0�:-���wu<��;�rtT��ǅ�@�B�!h)�r��dV{���|� ��GV]A��5C�H_�ȲS`:�䤹*m+��dv��U(4j�'N�|d����rM���O.���5�w��dq���:K��7���o}���\7�{n���m�{��S�n:?��#v�mԃi[$����"�JK��[�Eq M�E���sXR�t��Ʌ[f:����%�V�9���*h�&�MR�!���ȶ�u�b�#25F��sD��ɪ�(�7�9B�d9�C��*�� �˥d��m��� #�ie�spD��s��P� M�΀�iE�ǉ`�-$�
D�8.����L���x�bB��u�7C�F���5��v,�)G�Y��1:8�4��\5CVK�D�:S>�k��Y%�C�,UZ�R�LV�C kSZ�7��R!4�薷���a��FY���ȫ(\-�N���L�q�1)� �l�=�F �I7m	�jK) �#q�!hm�'ݴ�8R���@��X�p����iJ�ϪbL3�p�FY�p�>��t�0d8�Ԙ�n��V��c�V̩�� �h�_4�����Sq+�굫5B(���ΗRK��u�ZW���S���􁲊Bc~�:A��W�$^�)���]�v9@�,�rM�4dQc��K���A���4�;c�6Jn8�4��� i'e�<�I�bO )��5w\��4!���>�oD.��C���_��Z�eԀ:�B�)g�EK7�L����8�!_�P=�5������đ� gS(�Թ2�F���� FLW����.SԔx�P�"TQ-�L�9na}�,~"5R��r��iJn�g�
���rBm��ݷ!�ȥPc�q
qp�h�	���5M��J��D�Qï(8�X�YڴbD0ֆ(_�2R������>�ΐ��!԰�D�C4��Ue�E�L�)$�VW�R�197e���+j�$R��o�I�Ƥ��r��*�jW�:��h~Tq��#Ou�J����ڨ��4F�ܶw�uh��`��:d��O�~��)�8B'D
�ǁ1B��IJ���vD��G%��h�'h��#*�`ќFY��9m�)���VW�o�e�n��Cz���yd%V��q>���1�mK%�cS��95���^�$B��ġ0�f酌�BE�w�L��z�����Δ����V���BdAL�m�\?˦�d��B~��+*���h�n���A.jܔ�]߆@04�]E�`dBE�4P.�m�zQ`)qVk8�v`Ȝ�I�T9��)K��p��DWVHi�Z�@�BX�ҋ9խ�|�KLh���@�r�S��1Ub�*2���->G(�)'Y#2�8��ۦ�V	>���X��ަ��}uڥT�Y��S�����5������1���� Ͳ�~�n���N�U�i:-!T(��-}#�,�������A(k��@��B����n�@�R����k��r-�5E�!�	�ބ�� Lz�ҁ�BJsX=�rД��P�FQ�(N"��7f#8!M�#p��~��T�g�P+ݭR�-�u�W��	��8#B"R~�L_��h@!j�/*�Z���p�MGHb)�B��`�SA�.�8��D�=`�KG�Tı���&��|��xy�{�W����=F����'�Gw߸s||�c��W�^���S�XW>B��U�sz��Դϩ���4�|����Yg�CG�GR�J�D��F��p{�㩍]��x�㉣~����cnP�{ߒ+W�h�R��M��x�s��������~��_��_{\jQ�|"���#��=����������
�{�`����-GEm0���O>Z�/�m�kM>��.�n��3O/�<c�:���������l�������Ycw�f�ϥ���n)�nbt,v��٦�~�a	r�]��,�D� �2��9�F�8�#꒹��tQ��G}�0�y���dJ���]�hUpZu�1��R����*�Y/)~����ˊ7oݻq獓���{~��l�
fᆴG�o�]_�K�/d��5��%N��~m��������v����;o������_8w*z$��_�V����R�tdu�z�ZK������/s�!N�ۆc�<t攕�@;����B�%Z�`7=&����ߧ�����
��Z�#^]�=����(;յ�u(����k��i<pۨ�0��=7sE4IY���"t��O�Dڳzv,<�� P=�?��?s�k��> EY�ˋ3O�n������o���;����z5�;�q}�/���~��ׅ����3O��ʽ�Zߑ>>�׾c��t�W��4�    IDAT�{A����/}�����з�_���~���c��u�I�}8*�����/;�a�|���dL�D�[���A@��K�	�d~3���μiw���7�����Xׂ��1��)��e.(� 2񌂢�5�@Q}2QSY8��!��W@/|��MW���B���Y�� ����ȥ�&)=��/��v m�^/y�K�6��)��9��ҍ@|HcAHV"��4���		7��c
h�S��_��Cм�^�mW��|L�B"G��%♨��pՍv�&�o��ht;�q�\c�Լ���r	*d�[#GT��I��.��a&Y���`YF)�<��TX�����2[�2�@�T#�~&�#Q%�/��O#ІH�L�,2�i�j�Y�p�4���)p�@�dY5GHE��}�O�`B�����Z�����p���)Ԙ8�~Jr�L���1re����!h�]S��M8]��p�4#˘#*ˏ��E	Q�Û9�5)�Qu��{��F���"'�N���JS�I��U �G�s�a�K��bwGLN���
�P~=�niժ�Z⫮�6'�n:&�������1JG���൑ ��r(K4�6�/Ħyx�2:1��/��%FƩ��q�i�1�2���@����qf]E�U(�r��f5Y�(� Nu9q841;�zh�h�B6��� _U_�ঁ85�~u�qTi�|/o[��&�H��D�P�C�M�������`��YJ�k)�B��T=���]��n�|�z{+W])�^�zY�|�&�3��J���������Y�s�]>q�B�M9Ç�i!�'Bu9l��/�>����Jg���%��^��ɬ�QHܔI7n5_�o6&e�1�@��h)�nq�%2i7� ��d�.c"����!�AV�B��huI��/�!@8FU����N��k�xc|c��N�EG�!�3��J�@=�����$5�!$���Z�������^�J�m ʹ��sp�����؇j����/��6NՅ��)��N��$dE�@�h�r[8NרZ@NL/})ȅ'Ru>���h���[Y���KCf8�3�B#Ҏ��q�� �kSZ�p�:D���>'���-�ߞH�F̖	� 1M�ęV�X4#�Nje�`�疺r�S�VUI*ڌr�Q)q�O!/�vo~�q 8B,�t�tWߔ!��
��}h��w�h�԰)�%��)���Q�����dd� �}Gt�,�R�8�*��>�".��Vq���Jy�ւ@G���Ԇ۱�0��)�U�T�Y�CY���i���Rr�ńH��7�Ce�#(��Q?�!���ě�V���G����R�`�D���*���5v�ҁsҧ���!��MEd���A�B���<T(��"����K�/�%(W�3P]#� L��Z����%�:K8�C�!��*���1����7xm���Nxd�ȢpcՓ��D��*�H�
�6B�Rf�P�)J���uq CC��?߈�+R�F�uR�D�[�P�[��6� ���	�C�p�,�M�i���$sr+g8�F`��c��GS�M�ɚ�S��F�3����d���G�7�]qS&��|�&D3�HA��
l,S:�t�9�D��B�L
�(�
��VִZ��֞�)PK9�t���$���r��r�	tX)QE��I4��P��rLQ
��*+�A��Z*7
%9����@׈OP�L�s��
�RL[�,
��V]?�ĩ��� �Zҕ���e����uln���_ ���3�����}�ko��ӧ/~��������[�ө��(M�����K{�0��������P��m#��S02�{c�<���o���-�..�'���߷:4��ɰq=;:".�{!]Q�y�ρ=�A���8F�E��� q��d�N{���G}��K:>.����桌Dx_*��Pi_���?�c���'?��6�c�r�I{NA9S�Tu�����n}W����o��[�O��k���w����`-�����gv�Z��CM?PSk�O��,�/8�iLE��Be1�;ષ�#�2�G��>@�s	4���v5%�	�D3z����|���ʞ�	��Poa�4g�רK8���6��Ŧi��I��:n�<�Dp#�ʦ�g޾srk�,_Ż��̽뵯��垟*�o�];�4d�f`��<�������֣��������n޾�ƽ�~��ɓ��~r��o
n�>:�~�6]�ʹ���&�_2��xaᎋ�B�TEL��
BTub������3N�3������O�E�|dR|�)�k�ٱ�PP:���t�����zB�iv�4��0F)Z���#�Yщ��.ĭ�Cw&Mb>z�H�����^�Ƒ�lYn�?��?ǱX�zS�0�jIԛ���zt�d�w�����t�r�����g�~��W�~��o~���¯�}|z�̿�N]>?��|ws=��ܻ\���?�N@k1^����Rv���՞�u_���.������_������зկ�<�[?�Avz])Ǻ8F�ti�|�D8g;����3�	��Q
&�a��1�����d
|!#~E�>�7E��8����o ;l�������׆B(�����/����j	ID։�: ���*q��H����(]T��h!J�%� 7��^�-$c�m)BS#��ŗR� �Q������.�Oߨ���.��P{�@�l��g2^�zr�a�G�v�#3�fˇ�O�i��D���V�9��w����^l�(s��F��3R�-Ͷs���f�R���J�9LE!�_	��QV	&d�Ӈ��5��re�E���oDc���v8ܔ�+W�r#��JE�|Y"�Nl�!�с�&�j�Z�Rf�pY��*4�9��[�,��1���Ӭn��QfpF�1ɚr8p"ٖ�R�N�����Q�xj�f�|�4���;�^�zN���?�P4�,g�ɭ�����K�e���3쿞�3��(Z���ߴ� �h�cT�1��1�v���L���v�1��98��S�D�񩅨^cmWu1#�O��b7�Q��5�Y�!���6͗e5!>ks&T'E ��� @$��:K.�3�����o����Z�r�pS�m?!�ZBK��]P�z^��5�PK'Y
��.�i�#4~��M-�Y)�D�h��:�B�:3UW����nE���)ڝBj,G�f:���3�zL�h��1�Ζ����j�bu�֧�AR���M��W+�����������G�lH��JH�#�U�Q�ai"L"��(�3"�I�)dl]9���D	HE�C�4�jՃS����ogt�NQ>д�(����ũh-��7�V�!5�h�8��)?M�L�I��B�t p~�O9'2�i���:ض�D#>MmD��W�rmo�
Y=Tδ�-}��hԤ���MQ?�+��(�j	��(d�[�T-㔮�N:�����+��}�Cؐ�>�BK�|��ʜ�1Gb>)��M+T�F8��&�R)]b=t���	"h�%7�f+�b��D2�
5����f�9�L�cp#�8�;�|pZ&�l��k@4�RD�t�fE� u�:JC&���f�ж���q�k���F!8Z�aV��D:��F��k�]���@u�M}> �6ov���"������,�����UR���*��zk4GB�Z]N
B��PPk���]�V���.~)��R"$��R���^��p�c�-9Ycm4�S�nCʥO�NR�<��Ə��aҫ�'k�Ƣ�r+��BQ [%�W`;��>+d�WQ"�8Չ�~�(g��."dZ��iզ�����m�>!�M�ަ�I�Ca�����X�-f��՞��*�$b�A�A���GH'&p|�P"��T�l���&���߭���D��NG���i�V�!�J���.Y%5_�rIa�6�
і��Z餌�&�(�Ld�4N�KlO��a��gV]#�^8p�z��G`r��8:a��9s� �19�(��=eQH�)]���e���,MT�R�2F��Ӭ��MӤ�B���#����r�y��7e:QBS��������5���ST�����*d��)�1M'&�����(��BJ�6[d���3�KD�K�6,mZ�����Җ)״+���/�����7��G.rB� �[�|�@Y�T�f]�Y��H�,Q�)�O�B�!h9p�tR��؇dq8B��L������afp|Y�]M��o�|d �+�L�Zu��#:�����Ǿ��ٳ����]�����흟z.pt�~��Q��㽇~ :��!��<�����m�u���YhUݎq����o�}8fE~��jIi�cQ�R��p�̞ѨN��Oq嶷m }��p����@��t�?��?�k�OL����S�O��������	��������_��_~��y�fi@w��p�Z�ѳN�����ڦy����/����~�ݷ�����t�Xw���u�.�?�s���Vl��QϬ�5E�����*h|R��҅�F0�2[m]]td
@�>��W�˅c��%um��o���_��O,=�[���4VF>6��{e��jhj4Ս3Q���2ڶ9^����>��n����g#����XO;�=�������C�y������]��^���]z}�y���ݣ}O͎����E��{���y����ӓã=M����whl��d[���{��S`'�1e����}�+��!�w�����u�l��p�A�=��Ns{|��<x��g��xt�f��/��%��JG!;�Q��6P3Dl#�4���&�Q%�������IY�K��{C�;n94U��~�}b�i�nu��Q���!���o�F�nH�V����:t�֗���a�ܞ�~�����+7��x������[���Ώ�-�]��ʮ�N�K�U��im�t�Wm�ح��}����Ջ���+����]�=<�}���/��7��{|�	������űK��w�ۺV�ym;�����rf��E���=&S�K�麘�1f�h���t�舖խ(�I�\�9^�\"F�zP��ON+��B�\	#�+�UH�Nґ�@�It2]P>܉��8<N��RcI��>�Ն�[�e��C�(W:��p��\
#�e9�-�Չ�G
 �_?�B) Mg�t����l�~D��/UǱ��
�l*�ꁬr��z�
Q㮎�ZZ�J�P�p���W����3Lm;-DZi��P�� I@���8��m�(�N>Z�r��4�*��2�K}S@�C���_ȴ(_"��Ӹ)�fJ/Zi�dE) �9^��9��s"q�?q��=l�J	�B�4�6�<����@��XQ!�D����E���S��Q�O�Z]����M�|QW�����V
�1�tMI��j�g�^����\��LjuB���*G��4i��3��Ϭ�2��!�'B'��[Z��T�&�f4e�C�N�(P�j�)B�dE0�2�3��5��+Q8�Cb�\��'b�(G�G�d'Wb�����(��kW����d����D���*�t�ScJ�E��H���#�7>��8-_�V
O�a-c�
�OH�j��K���~*M���r��>�'���Q`
�����,D�uB�!���G3�4�ʥ#*��T"M>�!���.�jw3�׳W��`8g�����S]c7�E��`&+�%@�qun��ąXU N���nQ'\�J�U՝�S����
~Ս�q�#e��1���H6r�\4��EQf!`:��[��,�����@��M�3�dN�8�mB>��85��\PS�¡é���S�B8��h8m�)߻24��g�`*�A���rW(�Q��|�ZU��Z��(gY��^g8���8�z��@^"�u5k -A���\bRS��ږ����DV=dw!�-uB�*L�J��k R�p�����z)	*�����V4��I)��m��Fn	r9Ѧ��WR@Y�� e!�B3��J=H�pD�p6Y�����N�d15,w��$�(Cd���S���d�e5B��"K1�2��^c�p�SW1��5���j�/Tn�Fm�I������2Τ�i-B�(���=,
7-Z�B+�_�F����q��L��p�oԡU��rL��-�K\!x�i��CX+�C�h4Y��i�ۚ��6�LI�8M��4+7Q�	U1)>>�BaV����yE��ǯ��4�9	�_z
�vu~u���j��I�]��i�jA�����J�i�TY��wqSR	�r" �M��6�v~��6A�i"F�i��E6V���#GгV�s`��Fk��t���S�U  CF�Kg)wő��-���8�0�$�P)�D�XJ��4*e�*�o{�hv�G.�D���.f����A8ҋr��m
|H�I��O��|�S�VM#��ʅ3)�L(DV�����[BL#N�8�R��F!�&��CH�4D��Ь=_4�d��3RL黴� �-����b�AЉ�(��1�2Un���F4B�+뜤�JIU7e��k4M��b��vQVW�B|Nw.>�@FD��y}�R6���fj�'>P
��4ө��v�Ul��J�5��@S 5"}Rh7����ɄT�,�TV��|��1q��E0��i��X��E��TET�6�j��:�&:��ֶh��\/
�·4�[��>'n:%Z��>G���9~��kxr�"¡��O!�M����G
2�ZR(#!������W'�/O���5�L�����������ϟ=�\hU�ť��cOin��-q�E2�SP�P�+�o����Cor�3�}���w�<����#.�ve1!>�e��-O^\�x>|����X�O�=��MW������:���x\�T��t��E��?�C��)��
�&�r���U��%���nRdX!m?z�ȳ�O?�ٶ�X�ꈓ�[]y<��ሿ����_z�ͷ�z�������W7o_���󍯿���ǟ}q���j�ǚ��j����ئ���A��(��v_t�m52�U�Ш.�Vm�(0��B.���p|�������D�c�6S9|�F��*��'�������띜�[�}�ǡ���@N��Ӆֱ�z5ר�,�cW������թ��>��<�w����_F�'
�"*z�u務�R"���$�� ud=�ڿz��'׿�s�������o�+�����ӗ/\�g/싩s�9��Ag�Y�C����зF�/��e[�`;�jZ�g����w���N�����J�����2d�M}(�����ua�-�hJ�9�n��]�׌���|�1�'�����A�q�����hk$� ]��hZ�37���x�����=߫��@㸠O~��N��M�_�|�*z�wzuy��o\���['�{�_߻����_��~���}��̿���+h��Y
���<������n*XӉ__�\_L<��/M\<�|���/�??<��q�)��x^Y�ū�ΜkKԧ&�eRo�*j��2m����
d��+l��0s��d|RtLE��zA�8-��%� D�3/Ǟy{���e�3)�19�)�"Ĥ��*��_'��T3ʥ���#�5QH�#m����(q�j8jz�U�5�L
M2K� �����%���t|K��L�M�.��������G �k��D_��)�)�U���V�p���#����#�U-y}pzIq[�|��H?��V=w`���(�-�9�0�Q����B��m{�@Ʊ^R���8K��J1u.q%l�M#��M|&��l�����h8Z�7��_���� q�
#脂\)*F�����w�F����~/�v�� ��BhM˂�[��Ԓ>%q84�8D�Zem5f� a�l�!jW��ǁ���\�����ő����w[�J%�F�B�sꄦ��ć���̹ed��k꭭s�q��@S�UiɊ�*AB6̢D�u��5�W���b�Gu>�k������rL�8�c���\Y���+jER�Bd!�c�ֿyB5�0ʉ�WZh��@)�����A6�kS-]�X��qZM���H)Kh�ҧ�,���p���ꒂ8$4>�%ʜ�p�uh*��B�X	`�tL4f�F�(ҴĪ��mS��gHuU��͛���K�g4Y���]=m�J(���k�[o�@P�QHM]\Q�M9!�e�+�1Z��U�T����+*�X�|T    IDATZ?�rI����_��3'������\`��9p�/J��\�6S�� ��߼�pZ %֕)��
������r�tX3FS)Ѫ��҄8p/����T���h*vA4V.��r�3}QV�tN��֤1�RL��t����&�v �(d'���/�:|#BQ�n
)��f��m�J���-E0I�sGF+�t��R3VΪs�6�}H�t6��(� ���ÄjozSn�N��@�I�ƹ@@U��L�u�VU�fLSN%rpL�i%�B��_9)�H�B*���/wx}�1e�vO�o�R�vI� #^?��N�U�(:�ӿƀ5/1q��1Μ�� q�6�9��C��z�&n*�g�[j%�0�9+jg�F82Z~�#5!���	gh�ҭ�I7��K��S!>��2�T.}#Ao�|o�3D���.}�^�������ui�&�5�b��`ZE#��^A�yU�	1]A��@0絔/�y�ɢ�9����a�q����;�>�Lgj�K�����ֆZE�����0�+m�đ��_?1�p��ͩ�J���!e��	���c�[��DL�B8'eMꧬ��#UH�h:�i�n!��,V�`%8�	�Ʒ]v�6��crD�8:��r���rq��)W>�8!�E� ��>��b*ėUb��6�-J�i�I2d>9�\S��U���S���c���E�v	|"��V:2�ֺ8�`�K�b�( ���k(
gq1Ǉ C8��#O�!�$[�R��m��0"p��!||���yU�����L�1>A��������G(.ޑ(7A>�60���Հ�F��i
�rK��Λ*Ǉx�m� pH�D�Hf���
*�����m�tE!��E��V'\V��Y8�p�̴T�(�MIa��S
��|
���j�W�O�t#�A�8'���U����JPE
� �(r>���~B0�������	�Ӕ�ʹ����6
��[GE���}@�<�`�\#h$Ҋ(�).�\���УL_;Ӄ�:/޸s�����G��ɋ���bځ?Cw�֑�{����ĽE���H�']���P���dՓjm�DQ��(�o�4�X>=�d�Ӫe�!9��(*���g��E���~�C]M=�!�����g7��b��#��|����VDܓ&�Z�5�����}8O�1��|��o9>��6��c)��Ak���Y�G^G�o������ڽ7<�����ӯ���O�����������W�<����6Di�����Lۖ��d;W�����I��]5XDTn~R����iR鏯���84힍��Q���q��
φ�#Kw	��}��Y?��airjB����b�넣v��--��������~�_Bz���٭�/��]�:��Gm{a��3�f����Ź�qnk��v�Vz���z&��t\����Ϣ�|���wo�x<��֍ӗ�~������k-�ˡ�P�G���'�η��af���h�}�|;��hk���)t�����CM�fV"�g��v����v����lK1�*v�Te)gr{�3z�aw�#����0"���Gp���}�\T:���g%>����c�z�"�y���]�+SQ7�n�z��!Kp;�h��W���@!���o��>���{�7��:��'�/o�L�� ?Ǿz���G�^V�j�������������B�{��z�;c{�y��mb
8v�{7��/OϏ��ؗ�??�:�?{���]=_�_=��o7��L녘��ޫ{ɔY��8��o3]n!WĔ㢧 �e,�Ǟ0"J�spl��]V S'�+N�7t��l���S��)n�3
�L�>�\z���1�����.m'ntZ\h��aP�k��溣qiZ��Q��Ґ��(��V ���O�9Y��>�4�R&���4%b��tp8U��� YY�o2�j?~l5���>�j�8镨t�h���<�z�A-e>�o��Ҍ��/$ܤ�nz����v����0���1e�S�L�j��pέZhJs4c�"��>KA�IA�Ch�)����q�k �/hZt��Rb}Ƅ�Ni�Lop/t%�׹�
��]P �����h�Zf����GH"0N��Dz5�$�Q')#�U����%���0�8J�"���C�tc
L��dV�f�~.��q�]D �3���Ή �u©yjm�Z�ր���]���)�I�W���O(?/>��C�V�n�UGƔX:'q#3ǥD�O_��e%2��� ,���L�IY8ˁ3��l�Ș������,��h~Ҵ�t~�Ĥ9!8"ޭ�O�r� G��Urۮ.\R���
�nIA�"���}ơ#���J��i�E���"D*�(r
�R 5��~J1���("�o�U`�l��*-�S���2+2e8)S�aF3�D�S��"��l«�d�ҥi�L�i�%h*�޶�FQ|&��iLNu[i��(D�߮F�;6������0˪�hYF��+J�t�ݶ@
��\K��L!ec�D�EmE�D��8:ɡχ�4e��L9?N�3���ߒK�4#!��ճh���IMK%3!V��Z�T���j&sV��QɢŔ)4�J �I!���A������^]k�)�č�����bU�l�TT�7l�<K��f��T�P�FH�V����ZpN
�##����jBh�QHN!/iF��U������*q�O�5Jτ([HR|�iQ
|Hj�9u��kI"}Ys�#KdB���m���UAk�u�2��u�V�HGV�Mx� �#>]U���h_Z��x+�n:h,A
��1A!�V��kB��K 4�m��ܴ}H�,\�F��U��$�����	1�1Sd��d����GAT:R����@��d������Dv���B#f�L9^�	*��^ŷ3ހ�4��?#|:�?������@L��"Sc}�f$����>�P�ً\�����R܏�Yk�����2G�� �
e1N`EM1�r�c�V^9�*v���@Ʒ-u2��ʭ.���$�*J���KM�'�2g[ǫS���H�V��}��JI���ᰶh���P��}8�`۽+'jɊڍ!sL��&G��F&���BK���5M-�8�\�NV��j��[+�+S�pS������,�Dح;��W�_�Rr�ҏ ��6���#�	�ɩ~�9�'��V�GnOʢ_��N!_�������dՏ�P݊F�(�)V�r�׆( ��̘ҁt��M����L�MU�O�6F'�H�&GMS�(Ң�H]Uzh���x�V�#J��I�*��V��~0��P�m0$����:�E��k�"�+)�^�L�NuN�1��e�3<_IQ�`2cj	*����5��*G�%BY�T+B(˘oQ�ݶ4�pY0�5-���f�(Dh�p�)�*���<�G!�(N�М*hB��G���A �b��ǧ�N�	N.���§L�>'��@����J�r���V�8Z�!L�h:���W;��}N���t��D��/�/o��8:�8_��{w�WǾ(��ubm?,�N�CoZ�{��&-yr�O%�+o9�n�Çu�y���{�)��1��m������{�m|��IGu������H\!|d�A�����~:�hQ��7Q��?�W���88r} ��]���i��V)��y?���'�>�󙰢p?�<�AS����h5���x�#�|�g]��hۣ�������{���=~��������/�.�,����ß�v��w����=�峫�[7=j��:��� {V㉚�n��QEѬ���X;�·:��"HG0��^p���YԶ�D�o�X�,�}�K�9�2��/�w�xFWK��	�2� M՛>�!�J7>�K��g��~嫳�c���N�������'\k�<;_��t�������Ë�%�^Q�|�3g��8�K�Z����x������3_<�}�����'������<�s8>=[��,�^��m�S��7l�D7��?��o��oII�;����A���z\��q5��J0��Kr8�t�o_|����[�vI�!V�}�Ԫ�p�b(DS�e ��
���A���-�ZkC��4�v� [Nb-�%�Y�G�h�Ba�M�H^P,g������^[�y�K'7���wI�|����[/Oo�_��l������/yv�摯��Ҧ��#���l]W�Zط�]��~p5]}���c�Gȑ/߮C��џ��_��{�o^����X�N}7w�V���������;�Q�B�w�9�)�(��%L!�4e�h��m�P�/"��ҡ/�C��j:hp�۵��A�H�N�h1M95�>���"��ZΒ�BΨQ`���荎\W3���u`G�9q��VA�Q0J��L^����Z�n�F�h@.#"�贷�p~�M	"$%d�%"4R�1� ���������[đbt#�"�v���1�h��5n�%XHc�M���*�^ʖ����+����3��=�Z�LS����V���5�����ƪ�Dk�0�ti�P��!eq�x��d4�I�98��8���g�֢�h�pj���T��1U�lx��Ȣ	�|=c�K���)K�CGVq�7b�]E	��C�8���Li��|`���I�:�-S����D�"���%H�Ⱒ�=�f˫��}/��E���hA0��D4j��Ҫ���9uY�4��L�T�1ӆ���V?+e��Eo�6�#+�H�y�\E1-� �'�������2��[)���7��L�t��U��B����1$�1٢ZMJ�� i	�U�)m?�8�jճ���VM�)D�f��u/�n�K�8�B�p��HD0���T� �ᧆF��Z�@�V�|��'4S�B����a��)���J�Ƒ(d�d;_W��`���i2��IX���������tPE�0�~p�����͈��R"�JOVnY�#�jJ��mC��t�
|�.!&��S{�7B8&�Yo�
i�UX
_�H�Ti4��3-�����0	B��@�B�����r��:�fZ��_cmRoFVi�����oE8�N���/TPV!N/�hFY'<D�$�u�USQ#K�e�W���P|��!|H��� @ԥ�Az�1
18�&�*
1e����dq��@�����!X��Z5Z! �ګ�lQ�)�����Qh���k�(��QN�^�!hk�73�**]��0�g�e��!�)>����tRਅ��8�*d̉���8�\�j����L9N�4��� 45�rX�5f-p.p:�ўf(0~Ս5�Pb�H�8�H�%���6��J�Xc�^�I	��&2#�Z�9 8S��h�B@���tj,$ǈ&�I�һ�N��pi9@�~�qZxd�sk����xK�����{B���*ѿR������I�̣�雨��LC��5�>q$��UK�0T�r��N0Mk�ffp�U�l��B�©O�Ξ��a
E���lJ����O�E��YS���"��~��i���Z
���������8̶��~"�-���8���v.�c�5\[K;���BU����g��N�R���,�R��J#�1�!W����a���QE
R�����r��hd8���r uɟ1D��/����St֋�L�c�q����v�`�@����RcB��Qt@��1�v�h:�ޫ%��L�h���@�Ϫ4ne׀�,1�Nx�NB�pL���	1��(����r]���:"g@&�uY�M��RNi
�H�Bh��X=Lb"M���4��F��aD Ώ�����CĔ/��f�C��|�çl���K�b� 1�㤃�HL`4 �+� �KO0���@|N���ArJ���UQê�C�d�
��d9�c�Q8���FۋCJi�Q�hE982��ʄ�m�r���B$��o-8�d����W�}�a����f��!�!8�խ����H�
�h^�
I�{���R�J��p�P"��\8N|S�8�Y@:�|$2gM�%�K�h�l��[��	w��ZF�"�89�}�x�Ɲ��>��uut~c�_M�ِ��x�{�A��Ç�����B6�f����g~����`�X����Ga-ܥ��~�_yc�'!�7Q���=����{��YH��i�?��[��)yd�I�-�buD�H�6|��=Y����s9|Q�����?�;MQ"p����R�&��X��OD�y���u�KtR���X�G�ӿ7rj�g3_�z���?��O�h���󋳋+O������������������:�.���j]�Smi��7��K���|�1H�F��2�%2����p:��0ͫ�l��u�zK��B��,doC�����+�dl!�'!̱��P�q�w��2���$��dZǤ�J�߼ӏ{ݛCS����ꋳ�/����G�gח���Ci��ե�<t�����0�:x=���3}�s]��pvw�������7߸{���3��<߻�u����ݧ��W3{�n9���çOQ�a-=С���9����3�i�,��<u���;���}�����R�e[Aǿ0]�x�e������sy�I
�R��G��	%)�m�ꖣ�v��Τ����G��1\o�_]7�M�[�,S��,Dm����`jMc����ٳ'�_<��[o|�ݯ�^�>?=;=���׏_�����o�T�>�=�x��ͯ>��R���`�6]'%<�ԃ/c�XϷ<���s�N�����i��b�׉C/y�g�W/����;~}������[~�g����9Y��׋)��;&+U�B z��PQ��|�Pb�o��'E�o�:�2�Q.������1�G�E��.�BN����'H�O'�d9�����6�.Y�g@!H�X�Ŕ�W���9�3��v�����^�41�<0\] _#B���l���N�Iѭ�)G󢲌D��刚w/xRk��[��� %�h@���q򩵟RT��7N��F#��6�Lg���e��+ʧ�m�����O��v<����D=TT-�o����g��V�
k]5���~���*�pkymP�����-S�	�W_!���rU��mER�8������8L�6�e%�A�=De��B���Ð�R�#�
i ��9�� �!c�V+f��E�cr��1"�D��'�X4�@�"�O���O��a�qۺ����DE�3���Z��!R�5n�^��N
�QWLj	9�@/e^����c��u��9���\-
�f��.�Z�L��߈�8�B8m�`�EF{���!Hi������R�N)����hF���&%�!"�/�l��[!��+��,�7*�����5�'M��ӥ4j��-�nuS.~%�9B�C#��N��(�,c=�1�U��8%F��PKZZ��PkA�\�2Ǌ�1��5 ь
ɢ�CA��Q�S��19��	�\)S�LCܪ��C�OA��ģ�:���%vVZN�b!��E�J�0!/}��Ӫ�e�8B*:�ƚT��L�p���C��S��˪�b�_���:���
��}�RIYJ��A����p4��X,��Wn��14
B!-��j�^5Y��q	���y�޵.
�DQ~ⳇU�M��|��A�Ú"3 �|N����U��L�K�7M��c65R jc@ȴ��\ H&7�8��C(� �	v���L�qD8�˭O���iE6���Ň#�""�bwP(f���p���$%���#���mPRW�m�Έ(����88-�SD"W35�4�_ۚ��TK4YRғ�=�ˁ���ΛJ7�˗k��i�tSF'�C�k&0�RD#�� p���Y]����k�E���U���]"r���V
�r�$&>�猯�����@���>�uk��u�W��35i::�bB�MK�`g��B�I�r0�� 4!�.��oG�3"������7��M��~:�)���1�Ṅ_�:J�,�;I�B��UZ�Q���D�B�����[�5P���c���˴�G-��[K��sDK�s�:ꢦ���'�)\{&�i
�]�� A4���W?�!�S�]/�,&��QC3��^4�)�m��e�S�O�����Y��n�G��5�j4�����d��[H9�P�oQ�*��/ר(�>䤆�(��lEI�B����Ln�,cuC�9�K��pHx�oܲ    IDAT
j���{'�����) @�k@ö�g�"�dpH��8�h"5�\�r;�����D�[�k��)�&%�K��%QE��hD�@�qZ�Z@d�,)������D�0փ\�r��7e�����Ϗ�����1V�gB��%I�>N>&g�0��D��Ѧa>��4��,�Fx:ue���X#�8��s�/���tj��ᣱ:W�7��CS����:B�~�#�N�@�h�C�� �P���V��t~8�d�FHd#�Lw���:���o��,A�U�h��4��1W��7�,Q:R�R���+-���V�UuS|��|%p�t�Ln�)�� 9R������(EE:�1�k�O�a���l����a����jp~K��	ϙq���˲�I���j���A�2S�8�*���i4�	���� +��DP���&e*���~��������,Ƿo�����`�o��察�>9:>��]ʹ	G�W/O��Q��-���E?�n�������P~��C\ew��C~:i�s��>��6z��+k*$�Y�Լ�	7em�%� @�G�U���HJx�b����@��Du���g?��+_'@��.�V���佋�4�z���7xU���݊��sV�*R�4jJ������>y�9���������޻{���9;�^�.^޹}�����}�t����'[G��.k���r|�jϵ����jl0E�g@��8��o��^	L�(��Qb�Wg���k�\A��.	i�%1bh����t���t�'�]9S�(*�c����h�GJ���3Ϝv���_y,�[�w�.����zZ/h�e�o�;������������l���ZG�j+փ#y~}p��o����{�������3�S�铧��m�>
hQ:�g���Epj���η?��x��n3�2u���W�ݖ6M:]��ԛWN���G>�%��*犢���J�´�̡����"d������"��+j4�US�]8�Jhբ�1t����+�U���`�h[�P�n!M���k��W)����_��������
w�x�맏�}�;_y��&��}����������.�_P]��k�-Ғ��d�G��G�p�:��N��Џ��X��~%�ᅛ��|��J��i�����ľ�k�~@X��)��^�p�q��eB������g�.��zu����D �x�M�~f��w�=�`��S�k}��@V��[Nm�">GEc�a�Y�UA�o����J�Iб��l-N�,��BN���(�	�L�q�Y'����tc)F:E�F[$��Z���)GbdS=�����[��dǻ-pRvm�S��P��*��+aBh�1͌o*J��K������Z;�8DD݌�[\��ow�����$&_.A&������>�ȇ���.8��ji�c�h���u1&"��C�C-ǆ�[8')N���ı"j�!XYD8��J~=!3S�k ��i;@��!B�j����i
7�v#S��:4���#Āȍ��|8U��۽V��4Sk�VQz�O(�Z�EC:A?t�ve`y���br�de�@�Yr�
�τ ��e*Q�ȏ������jU��������~X�Q���:�~�8â]�������6��kE��C4c)���r��B��� 9�1g�9�v���G���k�Ժ8�.��&��*|�"ȭC~�_	����6��r�
�N#����U���f�d
|�B��iJTEu�%�D��_N�rd#����/4�"U�B�Z�NT�t��/T�6�M
����&"�#�(�H�h��I����f�3?5嬂�ZD��ll��h��i����RB�֛�i�v��f r�'f�m����Κ,;�sM�s�̚QH�
�ģsxђL��m���O�Oh�҅�M��>M
@�P� X����3���f�x��(��?������k�aYM��J��b�D�H��~��Y���C� �>LI���%�ͅ��k��0�zS�[�Dɝ^�Y��1��"�Y�8�)Y��|ɢ�14�2�V��JVt�\ky�-�<�i�W��o���^� ���c�X^�)5J}���Pܲ�/�U��D�� f��L0�ڬ0+����fڬ�ʼ�R�͘$I��]�M+�	�F�7Ԛ,_��%C�˚Kٶ�`X�0�lH�I0_xCJ���;�1O0$/=Ӝ�!���&-%ZC <�K��F�]�Ќ$��09�Z���89fj.�����42G&��,7$�0�p!��1�
������-Z\�%��l�LZ�x�ܙJ��*<��ʤ� �%�� H�uՆ):�Ɨ���Y�s"�
�g�i9�j\j �` ����iDd% �G�E��u��@���I�&%Y�� P!�e���;��D�V�GB﨡�Ǉ���t}��%�<�zMq=��#��%o���Ӡ�[;�����ߧq����`rp�'^�E��ِ�K�ch"��K����P�a��3���)��u�s�8$Y���|	As�\��!�����[���EPw�RsM��>O�t�kE	 g�gb�o���q���Y15`^B���7�
+��Đ�'�Y-��	�Ұ�FΥd~�aH��R��	���ze�?�f��/���2iV8Ʉd��&F3�&0�H^L����iF���\��L���Enx=hl�EO�o���Dť �i����;���Noh
L��1�Q�jD7�SO��Q� sl�3���T8M3�T�sde�' �O�T'�L`by��!^=��0�˦�/`%��'L�ꅫz����z���L�9'4�`uT.�/�\ V�b�K��x�3�4Q�0e"=��)�A�,D)(�F�$�F�8(�`s��V��A�#�Ú/�?_29D^�����@iRL*F��>��o9�d(}&Vz}Q��Ʉ��a��������w^5�C�d�����M/�4�4�b��gh' ;���F�j��z �	Y�r�k�E1�盵(e��a!�&xu��"�Ӵ
͗��E�Zq	L�$��28�� `� ~z)ѐ�+���"O/X��2I��~�rt��e�-��#��;o�U~s����<��'�޸����?��C��h�+;A4q�Ay]vg՟�t��,[0��O?�����������~������q�q|�ˤ>|���O~�<�L�|����=I�c�±R��+.9�4�#4C�|r�5��ǟn�I@�� �[sm�Ѧ�>��3W�~���%lv͗�7����G�\rsk���b��[���%���W�����w����7��N�wv��/<6���S���ts��c�f�P�	A���iF��걚��h�jB�R�V�Z���\r[N�g��/�J�kdM,K���my.�h�=R.U���+_��$*%?,ӈQHCV=M�ZV,��MC�c��yt|���~��g~tt��t�l�u����#c�i��:�t�2���R������R����>�l�gE���Rlm���x��ރ���g/�l�8|�ڏ�������#��R[�LM��(�]�Q%���O��4��lJ������d����64p�����������X������G��0�p�ᨘ"b��
6��h)�{4MV�.���IM[m,���o-�.�I�̝����}`͔-B;؀e�,u���?�ҳHY����g���퇿|�����{77������Ά����r$,_���Hu|�֙m�M�Ǜ
'��|c��o9���(O��ڕ�*��������<��+�(~����4�������{���y�^�����i�	�a=�f�z�e�0p�o?�����o�s��Y��ҳ_�VPa�����J�|"Ts&A%@�0���e�Z�qK����LZ�\��&+�(���3涼`3Ab��4 �b��	v�|`�Bb���B�4ZA	��  M$�|�9=�/���m]V�<�TX;��?��_N�2�-�~}9�0�z^5��^&H6S�3@/<����e�&��kd�!+NS��c��I��* ��*��&ŗ��9������.
JQ�rN&T=l�h�@.�|��u<�����`8���`�/��!`�E��F	-��!�����iJ#f��"x���dAp�iVm��&6�"��Q ��&XJVC3ҋ� .��^S��/%qc�O#.%Is)72��dc�fdQ.���s�,�( �\�P���U����elP�0����`H��cT�f��,d;ٹN�6G���;�..�e��4	*b�iȋK�� wzC���$Tɐ���`��g�@Bc��c��p�s$k�q��N�a�C/U� ���	�E ,�4Y�+�	+%J �4&�ֽ�D��^?s���!Y#�1S��H����4��p���X���o���f�f�Ţ����8
])X�?�8�&n�ZYa�X��A�'_�L��6/��G��#ӈ�lu�g����j94^B�d�*�B��Y�	�-�\4���D__2�(͔ϋ���u/�|9n
��o�i��p� Y2���:f��Rl2�F,B5!����d	ha��E�1)�L�_>
Fм���K���R+n�x�˹��g�B!�(�4;�x���B4ԃ��oXn����!=�^�P1�3����m���Oɷ=ɗߔ0����L5C�&�E>E�kLr��"� s:ͱ�����Eh���Mxp��W1�Wì�-Uz/�44_��h�T��6a���9��s	Ty���\J,$��|'kT�搲Y�X��8�"JeoF�`(h�� S+
Â��@J��/�b��r�3�h�xfi�eQfIe�=ǘg�;:�O�iq�y��7_�xf>�υ��|p�?%�F�O���Uk7�`���b�H�+�ִ%�����-Z_J)[�j����Y��	Z��6ke�2i6��L�z�M��w�n�=|��'�i�FOQ��&Д��8��&����JO�7)A��"�-�p��1Y������|�h����d=�4�e���}C�i'��K�>%p�ELc��( $��5Ukڔ�@V�� s�|#᥹�u�ۻ{5��;�\Z_��j3:��	�n�h��d��O��c�N\�������f�<B�2'S����P��\J���,��	!퇘��KF�W���HF���>�	��^Z��H1S�oj��F���-�d^i"/7J. Z�z�Q^\h�V�Nϝ�4��E�?�� ;@Ŀ�T��% CI�L/��g�Kz���z-��&Y/Ul��Oȷp0��Q���s)+V-/�	p�&gm��2�|�τA�&U^qF��zc�C��ʞ�X�QƐ�����UV�h��\Ίo�=�V�i���R��hS�N9� ����*	A�0k��H��^�-J r��z<�%Ќȅ��Z�r6��Y�	[>$�Qqa���;�;Ņ��XT�6i�K�i@�����dxH�d}9�+Z&.��V��-� �y`J�[�)��t��_�G�a&�U��f�`	6�?/z���2��9�BE��bՒ�j"d� ��4%@���R"!�%(X�4�mʆ�U�
"`B�i�G������e�1L�D{z�������o�Z�ÃW����?9>|��ݻ���Y~�ⱇ�u����?��ͽ����x�a��Db��+
~q��8�Vӫ�ǁC�{��ٳs��7\;�K��Ы�l�!g�˺��fWV��.��O>��t���9� I	�K ٳ��H�*8��wsO8O1]P5w�mH����!_w�!�/"�)`~��	��Y����Y���;o}��ן�>�@���`o������/�}��_���[7v�ڬ�R�3�6l��MA��[5}�&�\w$��Q�$�>�mE�9GJ=�����2��0a�L�@� �@��rа"l�+������'_��-��q&"������<rPtQ!�M#=Ҏ��Xe͹9L+G�_�3�-漾�^�8;~�j����j�гe�676}[��nl��W��ys�B���MOA}as�%F?W�'v� ��瑙�y����V�s����{?��/=��E��g���f�皠���d۵��T!����{�d��߼45V�4�?��ϼ �����{�Ņ�2�����p��ѓTi8�=z$(�I#��Q�Ё����>�����Ao3J.���\�GE�����!`p[5��XMS���Ձ����W�.���sVS����s��7v7�R����������[w���y�������W۫��=�s������#�e�yN��u��1���o>�9�M',���~�v��d|,��������ٗ/>��ų���<�tJ�!|�s���Lgr陸�R@k��_�r0��L�����^�)�Ƥ�,s/KH�dVB��a��l�,�ӥG�v���D>y y�i4&C�jNX���Ym!�eM��5�-���d&`�
M��46G��%_D�s.4fڐ������ө�6������;_�@̅�>PY'^�͑Rr�:�!�@�L V^�S������7��\��i�+���pۻޱ�p�8@���E��CƓg8��U�V.k�����\j/!�!w�bF���Y\C���Ǐ��j��5`�4��"�FH�Ը��K\z��`ퟪd(��7�'6$4	2�q�4�z�I�@|U�kG�7����Ί���.aC�a�f�R����4Ȃ��LB�2DN���ʬ�&h��VgIa�+����A[z���JC`�Ib\4CM\ =u��l-WH�����ZM�����Pe�b��F�%��	9kM,J�06 H��ʐ\�H<�����H���3�YK��Lx�+Y,9�3��� |Qٽ=������4�JݼX��0�U0$��[��r��8-h8Cra� wS� al�Z35��K�ZJJ&��k ���f*�!'���(�$/��Lræ�I�{=�oT^nF����2��ij��L�c  �/���)�J*"�L�v]ۀư�Z^()eR��<Bb9Z�4|���U)�㟎i��h%@��.=��L��i
�5��)Ų:\�L�Y%oO������)���Z2|iJ>x�3+Vg�3���&�ظ���OiX3�l@�ט�%�C��R��� �bCBV��O`�3,卙L�������~��j��/C0)sg2�f�GzJ�� ���e0.3E�D(��St���;+<��̉���h��E%"w��@�-(M�4LFKFH�3+���e�9��W0~0lEgBX������ʥ���𥏇u��ZAq�9^�)%����,=@���N��Kh���2s��3(A����p4�fW�bH�o^��H�L�#��U NCB�VL��	�zʼR�`#���g�\�"�l�E_&L�Q0lsk1 ��b 0���4j SC��L�s���`g����,�@��E'���&[Q P�� �3A�8��̝�0KRo.U)G!h���EK� ��d^�Ȭ���7#gW�Bo�]j.!\�Gs�8mR喌ʰp�S�U�^ �!�ƱdD���C��[U���P�lxg�m�@N�zQ�?Zl�d&�%$9k��"j�(aJ	l�-߬9%9+=_C�W�\>�����ƪ稀�rs������u��S���@o��`�DGH�UB}+���M��N/7�|�,��⦐��wm#C=�V�8f%��f�/�W���7}����h��*l&}�L�!�/4� ���L���
�̊<Y���E�y�|PQ�o�ǣ�  �K��L�����X���PD`&�`�/����|Cbc�a��0�ZB��4h�l�2��j������K��z�i�(	�s/J$�ä/bQx�	�dqZq.�.T����3�1ЛNz�`ȨJ8�K�P�5�� stLu�l�Z\���i���'Z0�h�Q�*�b��7�w^�$��jD'�&J��^C5�,�	�S�]�P�EVM(˪�2~i �2%L$�,i�(0%��^��d"��e�\8r�]�R�T+��)��	�U	�h)�Д9=�ח	& ��L3�(��k�Z��0!YVL8�M�az2rs�:��p�	\,�B�GI�� Z��4GrKIiđ;6��h� 4䖲�1�̗������)DHL&��=k)�    IDATE��F�%�c��BF����F��+����S��ļ�{��';~p�t�����[�������ف����p��|���_�����f�~�K���0s���ϖ?�fK���nR��i��&.H��4e��5�����˿�K���H�vr1����*^��ο�˿��(�w/�b�50}���7����M]-p���˺4<U�kF2wEE&BP���H�-5&�_���ǹ�d���:��;�y�/��\��Ǖ_�ս:��zv��_Y�W����mȃ�C�l1uع1�Ӣ��pz��Lz��*�!A�R+޶a�Գ&�$�)bxzMD�(0ݐR3�:$՟̄�F z�K&w g���|��V�ӧO}	W$�f�}5���ҊyIl�C�U��JYr���9���t������Nm��^��.v6/�Ш��8�s��g�_��{t������ӄ�-{����F5��ͷ>��l<+��ϳ��3����k��Ύ����8>X�m����A���M{���{�G�����L�������KY�0v'ٶ35@�1)�}��������d��mk7v�d�P�P����ַ v!/Ϗ�<y�pRd_A���~�Xja<�t0��BX��6��n�8�����f���tx���	�%Pp$�Oq�C�(��k���h�%�����y��֝[�{77Ww�����;��__��}�ն�~�����k�xҼ�k.G]�'j��ȴ�����ڦ��U: �����Z؋3_=>9>�9z�v��sr���m���]n���:}�s�vu�I[D�P^5�h�IEK'2�~��i)��!����M���B��"Z���w*�hT���;^|5�uY�U�t��������_~��/>���x�fE ���Ϗ��޻w�y��ŷ�����f��u~� E2W[�g�▌ޟ65[��a�0�;/���h8�v���<�!�FoX 2/ &�zzC��i�������-���M���B�''��L����v�ù���PR1.�������6����ˆ�����(�w�us�rq$��^nU�9Ҽ�,�u�N�b�1�� ���DĲ*C��5^!�x	��9S�
�Ϻ�ʆҀ	-��9꫰���AC���UR�����_&8��z�3��7�O}>QYFh��;�7�W��^�}�ǘ��a����F���Jm���x�&ϑ�8��@�|I�e׏�Eg�հ\��7�3_@���`�^�H@c�L�'�M�4�H�8� )#�Y.� N)L)�=�����O�vC�\�`���Ʒ��:�˽�u
9>9Z�'�7��:�l��w,�h�z�	��G��?�l�|=�{v�u���g^iGe�̦2��J�y����wqX�o�����}��L5!XmW�|��P35��^Ñ��C�`Hh�U}$��f��%6�@q�ii�R�%Xx��ri
�aƫ٦U�υ5��!FG��)���ǟ��A8���U��P��\2ˮ��[��8����Ųs��H`L�̙0�	��8A�%��ח4b�Ws�J\e����A��HO	Úf�K���/JiD�$�S��C��a�CVv,��X� ���=H�_?����xmw�}�'?��:~��b��E��εɶ����ؽq�=|����l<����K^��[�
NY�Kbc/�� X�Gb�� V�%F�2`�y._̼���<6�/V2B��\ʹ�Wʢ�C��a6�y�'��o��7dM)`Z���'���m.G�_�شU��i��
Ly�K_�Ŋ\�i��А �i�M�U�)a^Q�7$k 8�P&�b�/�a��ɋ��P��$�-e�+=Hldb�:��5q�U[��`��u	wz+go���>:���pUA�Ҩ�W�
H)��F_���)�oRS�V����P�B0ѐ�y5���3���
���1[V��UL���J����S=r���&�)�'s\`#m�(�)��
�Y?����@z����[�Ӌ�p29>G�6^�ږCY��P%��M_t�^�������L���Kx2��2ZIF��pz�dH��y�%�V!�=AmC.%F���Q��A���Wq�*�׾8�
�Υ���3^j.���h.G�_�=�+<$~2%��14�&%CzmV |�[�����S≿E�cN��'A���䛵(����d��-kg�����N�#Lo-]��rt`seh�zy*[l37��FHm{�li`���M�m��z�.� i:Q�"x9�~ʫ�ܼ��nԽ$7��h-��gip�L�Q�ҌȋfV��
�ojC��'�$k��E�����U��1_�&��f���0y��wn�۹1~\Gs�����+og4;�]�Q��u�(�����ʷ��8n^��-��h�/,"���-'�ӓ#�~=>�q��7<������7��Vj��`|�|V��
g.�ҐO%�SV���5�/M��Li���DB�В������ʁ#L�4��1�K����P����C��F���W�-i��(�/�-��d�>:�j���?'�vwQ�l	,/���5^s� �z�` �Q��	�6��~�׶���k���,�E���!�)�qL��͎	�Ɍ!S.L0*��P#�K�Ұ��)�>�F���^���^,���E�#+=+��R��SzxØ�r�ϔ��0�B' �ϒ�8���NOC.}�a��f�!W4�v��IU	L�)�F�V����p�Y\Ts���F�_OL�*�װR�jP���\�D�6���\-DҔ�u�X�
��Ԙ����dJ�Zƌ_J�ɼK����ͺS�4��ɉ�;�2}�Lf���(�Pc��L��`����/M $LH�xJ���3�$�dm5�U��[���Ȕ2��% p�:�(�~�Qy��M;�=�Y��O��no=���������uCu}�����������Ur���Gh7o���U�.����#�b��g�r�3!e�d�x��KnH�[�o���ӧ`��O���G�z��S��s�c@%(�x�{��ŏZɁU.��[����te.�Ȭ����Ph%CCh^�7k�\ d"�EQ�֨
Kñ@������߾�zkg���o��@eο�����_������ܻw��{��MY~������޼��oB�[�˷~q�o2� dE�KX�4�dzR#0�Έ�������5���A�&�	U ���X�[��������t���g]l����Qe����;�t��y��/�G�����9`on �'���WF���O7^��� k��~��{[���C�x|C������t�����[����x��޷3��@�7������ɑ�v�nܺ��;o��o|��rs��5׷|�tw{�&x������y9{�P55"�L�6u[�cQ5<��My�@ �&^��:6lnӷ�<WwH�y���K�L��\U-�p�1�d���������8�o�
�	�����.�#R?]����cۣ�����Nnµ&"k��}�X,�(�ߌ�	�uy�������J��"�����]��w��~y����c�����{�x��{��/_>��g�~�vck���xJ96��a`uƭJ?�l�c�7n���m\�7�6��=��V}+��ۗ��><?�5o�#�ãc����:'�q�)C+��)��RRj�*�<�Ӌ�m�'�d��Uٳ�WvO�5�;�l?�����K�	�\��,6=ي�.N���b��,��gV���x�� �����?��gy��dw�����|z����q�Z&mW����L�`Fc��ζ�v�Oƹ��xS��_�6���\xU�Y���4hq4ǔ�aH4V�c�s�1��^O̷)p!{Q��?�#��,CY���z��*∰�5ǣ��j$�&�.+	*/"G���a0�^�1��������}Mͭy���S�J�RR�Xh���I�����{�����P8#KϺn���0(��cE#4M�?�V�Ֆ�!��f�'$' @���EO�M<�"ʤ��R*�]#��Ӏ�C�.")?I�Q�+Fٰ�s�Bx�اZ�bg{<6��b�>�r���)�����w�Ow/���%ۑ�X��W��.+�Z�у�ܤ!(�@�U���7qxֆz`z`2=Yy.-�U
�
E�$�h`���S���F/['aM�F���.JM ����9#$D@�b���_���ū��mo�샃�	qh�i���˴��R�������x�GW�����C�{�'>Azt��5�%8�]s�-���W^�}���5>���C{7v�ݿ�p����>t��㐁�L#�吟S�15Jd3e�L�������H�'sg�'����[���\�d��$�eBr���=�`��1g�D���G"=˷aƳ���G?�?�Zxh�\��-Ш���;N��O�	�y�,='��-�v��e�E �b�S��BC������DeQ��Pr�W�L0��Pc�N�y�Q1)2/�1������;�k���^����#�%���������)���jlg��7wTod�q��ʸv]��d���ѱ��=�,g�k���D���:��ds�D#�&��XJe����"9B�Ѫ�kL��Tk��b��*dR( = *�M�\m���y�`��o-�۲��j�K��F3�Y�T>�6�g�,�%=�Q��+��}�V���r��U�R*�[Ǣs��`�LM��QQ
�Q��^��C���F�S�A�ðԙ�%kHz���s̥����  �Q�ū�8����b^�t���r�y
�ěJ.��>��L������1q��k�j�ѐr�ȹ;���6N�T���D�j>f{�� �c#�,J&��ij��ace3ԄȅP�ɦC(�d��1���6gD� p�b(�K/���0���E� �x�|by|��pձ��n-G���so;V���<�8;?�T�[���=���S�k�66N��r���&��@��1v`�U�0�-����x�q�+�4S�#��A&�j0h�%��K#!�Ԙ&w��5H-�%��1�L� �<�u>���G�JFГ�En��ѥ��z��ywoQ���g���R�.�dȦS>��j���|�0w=��k3�iT7^�5�HD�7�Rb
@#"*}rQ"�4Ԑ��eȗ	���4��"�ՠ��qƋ�+7�`��.��2�|�Ŋ�&��(��il^Cg�ݭ]�m�����UGyJ���B�e��V'k�x��Ve�M���Y�i$Y�+���rZ��	V^��Q�U0z-$+�(�6���9�a�y���o��6���A29g�o�bk}�M�ظ������y���?��q}1����V>�}v䉧s�8���������k�����]_����[w��rs�������i*�Vt�U3J��׫��T�͔�mF�Q�M�������� � CQ~=��8�~��>e�)�B�O���	4y����;
"�!�$)�xQ�u���X"�d܃�t������(������y	��D-`2�+��a�Q���ΗL(��s	P���T+�a��h�\"��7S���C)"��'6e!hdb+�c�D�(c&��D,��>�&��!L�	�/��F��5�' ��0zkJS8-�T��Q�	å!B�(E�swt8Z�g���4Z.���0Ӥ�N�Li37`�{�VL�Xl8�ȡ�����>|��́��~�/q��I�&�̷��C�^�0�3	GO�P����W��Cɥ%���p'�'��ф�×I5�p�F���^��ij�PP<�K��R⢶q���e^\(��q� �sr����0��[�r�����ar�*�$L	�!���)��*n.�7d}YMG���X�:	�3��d�Ah�<9�������l	����[��n��w��;�ܺ��������|�{�#h`G*1_Gy��4��^D��vk�]t�����z�w�w����N��EwKA�r$�.Z�#ï�r��1��tȾKC�����DR)<�q�0�-gP\9<^����9z�h�d��mޥ,��3eB�q�ݤ��|U`��[���Q>� U�khM��!�~(�%��;�n߸y�;�}��j��������Tkg������1XO`���#l�]�ح�'��F����BcB�(Z�
��k� ���m�D���<0|%6�4�`d�M����s)��ӟ�T�*�(��,�f|���c �Uh�y�� �iRh�������S�c�P�����˷��k�[�[۾��M��e�ln���g��$!;:8Y��0�	��^��KK��w��TFg�mx�������߼��·޺�`��
����w�^�x���O=j������kv��L�mGch_��tl�͝#�=g�{�=�=�E�>��3?쫔��XR7�d�dG�/b�,�g�?���~.O�>�/E����a��ߏ?���g�P^[Fb��,F�	���m~9X>x����4����maR40W���Z�G�9H_<-����k�>W��'�^�z���7{�o��ߺ�����;.�}X`ug�毾�z}÷��0��/;���@q�M�ɲ{���Y�?Xk[8��O�{���]O/�^}u��vo���xK��o����C�e�~3C};P�0��S��&6��d�1�����^C��������?[)o<��rԀ�%c [bB��[��xp�ŗ��7_�:�8=��Ç��O~tg��;�����?nƎ�zE�����g���ه����{>���g�R����7w!w�oܽs�՗�l%�������~� �s�����j��ɖ�V1#�f�d)���$TCl"�
�%�^���W���h�بj*�c�Q-���� C�q*��	S6�$�pJ��̐2=��ʊг%��vR+�B)����$���kh�LN\=�ym$y;�%i��%s��y2H'%M� ��cz�5��D�L���(�]�[�����jh	�y�B����~_[�mR�K����u���t�B"i}��&���7�^�z����9g����3;�n�;wx���ݽ��y����6��p��s��Ł3|I�Df�$�nj�4ՙФL���4w`B�Y@N�	�PO���5�@��(z���7�a\���=�v�q��0;�����X�EysmY&����ӧO_~��Ɏb��Zm��^~�o�oo�8��嶔�J�$7L|(m��3����;;���:�o�X��ca���O'����sC����]^���{]�[��uh���)yI޾�+J�f���$�hj*/ȹ�+Q����|5�+!*=%��dm$�%dE^0��D߁&�E	�E��H��"�Em����Z��Ԃ�I@߁�~g��bf�j�ޜ�}W+.i��/�`���D�����z��3�J1�͊<dz��%���Lj�)��$f� ���Ҧ/�嬗�!;/T���d��
���fT���"�en~��sE�˗�6��������2�7�����n��OC�V��w@x�fF�NQ�xT�1q�ʿ���2)�F����נZ�#Yf�*�H�!<*=}H0LH r��&Mʢ�d
�:�"�~�-�ON+T��U,MV��d���[������q!4*�f1u��)ء۫��f�FEN��	��Ґ��Җ� /_�`J��V��Y\/}�a�c�f�<�v��򩀆*�0iX�Ұ ��J8>�U+��|Cꭤ�Z̏W����%_��bˏ�>�C���9�8oا<�>N�냃��2ӗ��V%�&������ғ�^�1%�o�Ά��D�S"@�D�JY�����XzHyv�a%�#aj}�J��Z�n�l:���l*B�r�2���1�fTA�m2�
�/��.ߔ�^����N�f���r?tks��������b<�V��3�6�U^_�'�m!�L�NO�J%�'�R�&����� 3Q�3j������{�L�֫0�I{,g�Tm��'�(��b�%��>s"������3jK��*��N�iƎ^Boy��TC�䣕� Y��,�)]��t�    IDAT����F�~qfK�5}=<w�a8N^�&!�r+k��J_8S@��ej�����ë?��V /3�������0�J��L���E�Uˑ�,C0}$���,1�>��z0�+A�E����]������9&�z���P=d��J�	��#��L��Z�s�14͐�����I��[67^��r�펊7e�	�A�q��ۧ�F&rUu�4Sq���u��Ym��$�7��Ѥ1���I~~�ęd�z����s�>k�s6����3k��ޭ㣣o�s6�KC�l~���yگU��q�p5	-3j)��Pʙ,ɚĴ��@�E��*B=L��`���	��/ģ�)�ZzIr,�)0�;�};*|�6-G�E!�&�ċ`H}Jc����7>�2��B����})�H�I�l1�B9s���H�����H��XzÉ7̅�����ȳ24�	#4��7@!�K /2A�Ld0s �i4�a�4䘵㋒{<� ��h���֑��;6�}�%̅�M��/Ss�!�Ջ 0L`�4���b���㕒��d⏄�#ʂ���M'YD3�3͠vB�h`����>N/K����@����n�̜�!d�T�Ӱ��̥M/���PV����HChF`-A#D8�PЅ���~�f���KK.&�H��hc�C�}b����1\"��%�Svb�!� � ,N&N�1�3`��L���ƫ<euݑ�z��Eї�jH��E�Y�8ɔ�e�^mˊ��Rz�i�̢E8�ǃ!�RD��-�aGS!T@U5������h\�g���{���l.�R�8����n����g7����ޝ{��?��ӧ��)���Q>|��'�L*�Wg�0����?��?z�a�པ�ګ�Ws��<�q{V,��=�`�~��Q�k���K�{򢛝c��?��?1Ak<8����n�\|����rA�U[8M8V2��T>d7�E@%������'fy�D/.�/����>@"g<�9;?rp�k������_={������p�����=y㭇���7w�^~{`��<o���#�㘭q���eT�V���c�Z0ʦ_b�\�`6k���z�ҘBb�i�@ָ���k9Ɨh� S���u��OO�l먘��\�����8)��v�02��G�)��Q�,I:�J���O�n8%l�J�t�#�����ť�,�z��r�%�ա��V��?�9���2s�u�ۧ�g��9��硤�������?�ϓ��������.�t����x�b#���[�v�c���F�7)�z�のl���r��A�
�^������+�
(6��BӘ�]���H���ۿ��cW��O���'+#w���g�b9h%	L�P/���@B8\�a��w`z���1�=Q`G���,l#^���NƷ<��G_R��vv�^��'���?x���;[ϟ=������i�o�h�� �7��賜2|���ڨ�=<��;�R��C�Ɂ�.aD��[*ۛ�>�q����sҭc�НR��x��z�e�;�K���ڢ�ci"&���W;CH��KCK#Ɇ�PH�!w�[� z�3=��*߸u�����T/(6!Ȋl�TR�嬂�i�Л�x0�y�#kss�s�[�k�^��z~�b������+�~>���������?���gO>����ރ7�t��g�����or���~�dnÛ�FBP��9Ym ���@swR��4&[(�
�ě&���B_��
�t�Z/"@��E���0�����?��R��!�m I%�Uh$ώ��t��$uFK��țM	ԛ2+�$[��D�'�|�3t���2�p��ӧOrf����xc|�@����m��&NvJ!wD;Tz-�Pz���w���������4/zʩ�Eäe�����°�@V�h�f�\�ܾ/]2S�����;Vw�FI�{u����^>��z2���h�b��}�]@S��֎��S�ǳ���?]>�0�l�_��èk~�v|$��6N�17��8w�l��&�Yȓ#Y΄&�J��{VC��[,ʑ���G��@6��U�#$+�^c����@ՓҐLc�i�Vyõ��;!��^S ��p�'��6BhL�ͬ�n����%�-͟���j՛�~������w�w�7l�����xoi�X���w�ܺX'��zT���{��ǟ�l�����g7��8Z����m�����޻�,�m���[~
tg���/�=ϸu��qo���=\�v_>�Ja_�\���2���1���_&w9A���fL~i������8�(�L��47s����Q|V��6�"a�8GfK���|Z�y�ʬ��E'��L�N�\�ì�i���&v��A��af� F%PVl��\�Z����B�JY>���4�i"�b��Fo�Ľ|� �͂X�b�元R#kKF�`(e�����(���N���vv]�x+��ةe{ܱ�K7�d�3͚�k.��Iƞ�T[ϓ}����աM��p[�=���]�x?f-tө��.�zy/[x���4aTC#���3j����c��I��F\��"3�E�q2DB���p�Rr���D���(o=Gr<�eB�K��6�e-\x��������;"�㴑�xΣw��0d����@.�DQC�������r��$�`��ò5ê41`4LV�L i��i���0U	 +�@m�eFc^Փ^C[�`zM�L�f����S���}�xd3~Ě�jS,��0��Uw.�	W1\������3����HD�r��w�O�b.�hi�&��E��_:./O��J�K���?!+�F�$05��K��1i%C�,. ��� �jdSC/�酜�`������/��K������.�/|�^
��K�0��s:=�ϙG;���%ϱ�_��Pޥ�ѯF2���'4��VNA6��*�%���	Z�O�9�p��#UBs���e����4h�h�!DN(���I0�8#�'V2��u����S>�i?o��6q�肭�7��-���*8����8�8�!4���R@��S%�&[�z-���d��4�4���ez�V���@zC���,�KV����W�����)�.���4����F�֗썀[��x1/��E�GR��Р��W"KC������n[�Pu�e9�[�H|F��IkE��'kr��$1��������St��r�R�H�W�v�9I,M�	��s��|)����06���j��}��oo�4w���LP鏠^�|��a��nu��>0+�Y��t��[+�}��Nui���^��{�3�n���������L�rZ������H�ܻy����ou���j��~�ů|��-<�:���2_�GzKa�d����$��K���U�a"W�x�1Q2UC�J�if�A�K����8�� ��R���Q�!����K\�oیU���}y/��0qa>�f�e��(NT�;��٘�ə���e�_�,��t-\9�ŕ�F�*��H�4�	��!p}����Mx�� �T��@��^8ru#0�O(Xx���s�$4�M֢H��� �Y�p�sTH`$zÖ�(0��9�L���{&9��)`$@Ӑ��ܤ��k1ƙU/C�P:��p��ӝ#�)!�	���qg
�%+Brl�MQD4��YY0tnؤ�xh��Qi����5L���P,��#+�`��s'C¨C�>(�ìb��LF�/���!��pb#Ħg����6L󂁧�cȥ�I����U�/ G�N$�"pI��(E1A=GC�\(qZD&`zJ��!%�RH�� SkJ��hld����I#%M�`ENS��Y .�c5��^����I&})��i�a�[���&
$�|c�L��n9�z�*��\�Lx\�O�����#�?>w|��w�˼~u��cg��~���/�skj9e[D��E�^�*ls�c��/��G�0�ōS0�=d�j�g�g ���`�*m x=�������K���A��%�9Rܥ����=y��ݣ��O��k�U\�����d�K����C����׫���HD��H��,[!$�\nU���f��;�䁑����=���s27�.��ҵ�o�޿�����駏���Ym����燎�co�}��k�զ�^�>�hzrg'��S�����5E�JH�'�������b�Nf�Y�^>����J�����J�Ң�Q"�u*<�x)^�0XTWQd�r����Q�ǆ�2 �!��<4B'Pz�y��71k�+O"W��'�^�x}tw߽V�ygk'�X�i<]��ٸ�z>�2���������2j�}�o���t���|J�����틣����8��ځo������;7o��밒o���q3W�7&��>���:�)(����|v�c��:p�0�[�wel�?z��  ���"bP�'O��b�4�挧#ǁ!=���,<*	�A��l!-fxLV�[�R�����.��eR7�u��h��.~��ġbj�����(/^~��v��<c���<Us�{��������s\_�r����ޗz�j/�_�\�TiI|��K�X�qS��}�s�3��6���K�����l�ׅc��չ���w����`T{Lt8�6د��9��F�&0d}G�N�JJp�z	��J��c2�=���A�Tur�(�E��dM&�i��S�V��1���о2�p]����?���o������/�9|�B��G�ܫ���s�b}�#�/�_����������;ʫ�_��&:Bn޹���_�Yڳ�w�����>�K���Tˣ��S�d	(��`RZO���IX g[���c�����x�u�F��^.�\�C�4���i�7����mK��'������T���
�ɡIqU��ɩ�+�4�VY�`-(�r(��~6V��p��ˡ��������vK�~�;s��v��;�y���M'�ʂ�:�k"���";;���U7�E3��k�N��������2�}�L��YiZ=}���ɪ�b���uB�vDq���s�����<�}�;��mn����f��nicw���u�T�����Dwg�h�AA��s�6ֆy��^�u�|�߳�Y������m/
NV�%54��^���q{W&��j���d7.@Y�J�*Qj�0V��L	�04U����!% k.�Q��QY��H�P]B9��!�L��"�;�9��^�ѻ_�u�?{�O�~=�����_}��G����?z����ٽؿ�����OW{�3��,<><�^-�}|'bclB..���?	ptp���Ջ�/~� 4@˿���g_�y���w��b�j���y������Ӌc��9���:;��q��b�����w�[�6��p��⋯��l����ۢ���r��Z���z<!����;� ���R����4$k�42rѹ[�E�.8[z�(��NgC?\��ėR��X��I��'�Bw{�>�.��x�#�e$r s����S��f5��@
ǑR#S�9�BŅ  Y3,���Ѓ���1�^�Z�|a��|J}z�2��/t�qJ�P��	�FY�WiX;�8����������[C?���c�ݎQ9�������u~�S�{�6���8����;
�*gx
�c�iui�=ƕ��rP�K�� �!�F�S&��0��" kL`04�խpz � 1�3���hxʳ&̐ Il0��ci-ӉA&�\L\��q�㇪A��>���H��sFJ��h����#�.���m�s�Uh�bt�TX$�4JHq���>��xIFO�g3���00*ӧ9,���{՘��4*+2Mi��1���p����v;d�!'���G���[n<v�`<��1��E;�ؿ~��{����v�����+.�������i}�+�`��	���)5a�!P�V
H��X5�D�E�!��U,z��50r`�.��V�L���UJ<����9|+/�)�$�^H�j��K����G�ܗ���N����r���46����~�3�q���~	��9ﺙ>J���)�#���3�N?~�b9�g�B��D䬗A#�� �h%l��4z	=����pY���R�JȆz�a[��pAs�Vy���P?1ɔ��<	\X1 /Cߚr�t�����	zp.qǼ���K��eW�}\S���R����\�V !Ȗ��Ji��|!�H��O_V�&,S^Vj���;�t˼��ʁ��8 r��	@�� �6�Fp������x�ӻB�""�$_����������M���9:��I���4�N/�슼ʓ�o�bB���X&խ�'O����v��3#�o
05�NL�~F�&��
�Mh�xR�II�ԛ`;�0N���\�k����n�xwFä�6����9��c�=(h���rB��� ��J��vbO���H��;#I�o�6�����G��	��o�����w�\����*�e���k��O�a�>������m��f�D���^�+����B�˙R�rK���)MLg9�T@}�!��\X�_�DmGY��U�c�>rBJT4i�B�I��#1B��}��.r.�#�f�!��7A�m���@�b�8a����H�!`M��'������r��l�,�È�*9�L�g[�G>0�y�^����e��=��L���lx*�u�X��s$W+�)LN֚�X˭��&��4;��C����`�������B�4$h4`��
�M5�7#"A��%Ӓ�
_�&�T8Q�hM�f�1�)aQ*/w����)6����6D��UO��p�z�H�+!@B��d��a�0�rFU�2:=/J0ʹ����QnzC0!4k�� Y��=�ȅw-��2ݷ'|�Sm)�eՓ	Z	���3Qj�����sJ��� [�q�*)A2f�\J���[q�w�zN�����08;�1���c�����h��)+L�A��R20�c&끫��G1�4��\j��b sO)	����>90Z��ł�3a*%���Ί'N=��;��!`���QOF�Enh�/���}ut�̾�@�G�O~�ԟ�<|u��Ͼ�'��5��v���z��W7�L����ȢKO YJL��u��ѣG}�=��8Yg��l>\ ɑ$���W�fr�G�w� ��]�ݵ��r��@Rmi�w�40~�!6A��J���M�~��9��kB���L��-큫��n�^�d���ex�䩛�k�o����B�ޭ��_ܻu�P�q*���Gk��[P�K����ve$�ir2�)[�JA��-���zu�Ӌ�P�2ِLӝ)�4���'�|bq{��������?����.g����0���{��I�<|���c�f&��R)ɼ���Pq����.#�+���5�y���Ν��7�u�������� �p|	2.>ƍ'�㕕�/y�;>�n��y����������7w��r���ڿ�~��������yCo��
��u��8�㑪��ܶ��$o;�/YP[�~RDC�q�D�=�+c���������駟~JiazDю�4S v/۟̔�:�)�4|qǳI�U�=w���vmۅ�':���������,=S��������#��-60)����"��|�м�������ߣס"S�����g�^�:>:8����.�t�)��w�o��X;ܸx�s�������{���)h4�ZA߯�g�\��5c#/������ݬ������2��5�×�|���'N��r�v����Tqy����"�$��r��Ȥϴ�0^z�ۮ�zx�zoO�B!Ը�i{(�Q�glʥڔ ��?��I��H{�wօ*�����d����J3Ү�Dӎ�d������JZ[�Qܝ���}4� ��p՝����?r`���������/^\�$�<aң�X	*�S�,N�JA�c���ո�&��ݿ��������M]����&�.�5���`�dG��&��vo����>���iϟ�替�c�l�<�{���xy~zq�:}�����^��ݿwg�h��<>���!�h!��0T���������xNN;��h�5PR�
�tA�1�<�}<+K.��.��Z9~���k�|���e�(N#��\��ڜY��B���ՌL |`Hٲ�nn���%O�h2�����Hn    IDAT��%(�mnS�դʥ�b�`F��oߺY�}�J�QH�y�A*s~�	�H6��G,��E�i
�iL dH*���L����#5)a�b�"I0��$���I�amln#(�[&v� �X�vq��r��z��� V�z�ވV��6��,B6g���jd�%���M�p絟~:=Q�vF��t^M��ek>��O$M�%Į����9��W��SML~�T�Ӏ���X!�&�4�̛H���#��"�_?fY�L�\)��cs�w��v��S^�ka�X�^x�r-��V��(���f��}�"�S{&^Ɔ�������|tw9?�k2��a����8n�uM;]���c��u�N
����nɯSW�ë�p�Fu�����g�J�~u�pU�]�`��<������|�΍��J��\�Hla������Ť��S-.�7M�=������8?h�^���ɯkHA �� ֘�'��Ԭ%LMr�%%�c���$��g��0xf���Fv4��.N7���8�Fj~�{C�h����p�1��*�^��ϻ��+N�V ����܋	5%
)�H!uk��F�y"{a����ç��A#��P� �JR54�7_��&R�L���u�B��51�ē��G}52�"����\pKz��9)��ah���Uu��;%���MuI+O���a:5n�:�������H#�Y�����O�*I<������{X�O�8��B�KSL#��̩�Ԭ\�B�p'��EH�f0����E��Z�@ $)7���*�$��L�GHf�*�0��9 ��ON�0B�JJa����bȊ>'^���hrPAV��ˈ252Wtq"Q1~J,���k3�
=�Q��"x�d��� F)�@
i�TR��~Q���&�e'�,��91+(K_���#�>�ˌ�0�d��-,#�\��B_�͜�$M���qyiX�[��e��8}��r���is�^1���z���pJLuHP:Iĸ�e 31���S� A*� I�i���uOβ�(�8M����$���%� ��*���dR�'�5sI�{L��d�o��1�S
�:8U3i"{g�|J��p�{��Fz�8�5׽t�1b)KaO=�����9tB���{w���W-��^�}�c�o�HEd�T�����C��P�d����=&&��PV�A�,	��1�d�L�8���B2a%pr��#J�� |�$�ġ�胣�V��T���qp��^�yA�X�T��vmD�Y�>�����j5���`ٕ�#�b�����>͒��a�Ƨ�i�u���Kb���,R '�أ Oe�\w�H0d��_�L�����u���	 F�.@/��`f��I<��2<`�GI8S*�P<m���Eiy�  55��X.�S#�r'��
kKB���|����~�8*�ҘI,/Lj�<�i�,N���R�a"/����a�ǔ�cz/_M2�)%o���)6��V��D�LĲ�x����v�I�*����N���::<��r:8��&BgRkX�tDh:����Gg�Z�Ժ���$��.w7[�1w���ve��1�u�m{�(6c9���(+�P�=�#FV_f�178�kH�>�@x@�O�>�gj�em2��
&AҤ��	��,��C"��d�3W�bI���x� Y.�з�=�`�ˤ�y��@TJ1M_l�}M�ܘ`*>��jo� ���8�݇.~�ԭ�f��>� ����q/D��#[�qWLѫ��O�i���4i�)W��WZ�Hi��Y�&�*�C��7�O��IX4	C*WHe�,23�e˅~-@��C��\�<�X�@b!�˒��EJrC��d�� ٹy�$Ȃ[J�l�JWY3$��+EB��)'b�)�8�؂3�?[��? )3�*{��H�C
�F�� U'2B�1���>b��BJS*�0!3��2�+q��h��R� �ES�iUq�Q��
���JK�`d
%�D�S��Ch�����E5��Z�>7V�{�"/��7��ʛh0r����!-=��T��9r��a<
Y: �"$@���*k�#X��e,o��АA����LPD�d�`(x��ɗ���]�K�s�D�7��c�4 ��^8
M� I4��!Kѫ) ���
����3�2�a���E�����p�T:zEc���(I.@�b�d��TY�8�	+"�� o���q�Pp
�Ύ8��-id�?s�#�*{�.8����P�L�J��Ǔ�F�)+�nm��X��3:�������lw6l�S�^p
�^y���<�$ ��Ν;J��c7?����B&��6�Kk0|��	o�&;�,B�v}��7Q\ͯ�k�>fhq`�㲐���6�� ��Ǐ!-�Xʁq��#bk4ʢ��G��?�CR��?0%����?' &F&.�D���q��`��G��$I��WL��Yb3m;���S���)�l;�hH�;@HU��?�ST���5��R�,))�@@_�RH!���XH]`�e'7I����d4Y���%���KT�y����7,�s���D�
x=��,c}���XT!��c���c���GpJ���r��#J*�́˒���y��^�V����jV8��6���P�������j�S��:|1���ی9ո���l��{`w�S/U�ճK��R�sT���ü�f%?�R��W+U0|N� �G.H#�U5k$����d��b���2<���,�hT|R`�4#�6T�E���G�����ȴI��a`e� ������D��嗹�R� ��@<��Z�|��g�S�鰥��T���$��֊� ��V��Kkd�?���H�`p�Νk�����`��������d�Z���r������MÄ��6�yL�%9g7�T���f�]m�-���r�W��K��G���ii1���E฀k��D-��(d)����ʪeI}�u�^?�d� �� ��L �GM������?��}��bҤA/ȋ��$�U��-=��6mLUj���	�pi'.ut��X3޻����?������w:�������3ͫU5ޮ��V�8_�j�:l5z��Z�ڝ�}T>z���d���`T���l�t.�1�����J�Ľ,���81z��~SEӅ<�$�	N-�÷S���s耞"���iI���ҪX�+�U0�zD��F�G�X<�QŪ�>q�I`�y�xj8Z���y/��ml��TY���Q<J��B�v��1���vyҋA�~|:ʋ>��"sXN�$���qxzb�N ��	�v�ov��Vq����������떓O���r11)��iDGFE�YH��F��O�\�%�,$CJE�!��$ ���.���b�!Ȱ����Z(ۋ@�Df[�ҍ8P��M=��6Q�����bb����^�Q/�7�K�e�+�zl��֛�:;{�V�t��֟ONN��g��/gn�d����_������Ye��^�|�8�̆��ꥼ�DV�&���/�[[�/ԧ�>` uؙ
t��Zf7Z��bI�^�x̘�2 ��,� ��lI�  (T ��{�&'yJUP���J�d�/Kb~h�^1>|x/�g�O�͒[ݹu��_~z��.��]2Qi��.�b-p�3�����֦��>�[��lq�wnv��t1{X�<��Y�}�Y�Z�O�g��w;�+��gǕ�n�$�Ui�Yi�(]Z�mu��ht����o�%}�9,��6*��V.󓓲y�x�sŴ!���tmdӰ�d���#���@ɆR׬Ҥ0i�L˒,ț�j�� KJ4Y�G���)'b�6���}���Ո�S�^1E&����9R������a���,�W�Т0�{��lX��z|�#��6Q
nQ���Rv2H���,F9���搏������)��d(��� �y��kV IB�%y�d��R�K����Hf��	�d�X>Ь����/���l4:,[v��r�m:�m��j�Z~���,wj�g���YTj.��!�Uբ���o̎b��<cx�{#|h�
߈�ǐ:�0�d�	����$n$a ���6���X���jE}E�Ȃ&u'&͛.���̕�d��0|Rf�I.��*��d%�e$�8;�J�ZN�`"�+�l���¹�v�7]b�������|.(���Y�8q1�-N{��"N��*��R���D d4���)sr�{��Z�+��r�O}0`v�ڡ�\A�f'IF��[j�vj�.>
����I)��4�L+��� B�����}�0��F<��G��IS��*�xv}

3��e�>z2�V�>mԼ�l��w� ���-�K0�
t|�ŧM��,u$�Ѿ
��i@d�;Mي^BA���B!p4�u��O��M20������ �a-a`��º �0�����IV��Xq�̸�7xH��$�����K�U�:!�Ë��>v��~��/��{K�o�9!iC}��9�bDb�\��7���[ƌ[i��<�,B :ιƍ��Q9�d#7qd�8$�@��O���0i!vQYbxę1�C&eb�i�u��� HXv�|� �	�rl �,�f]P���1	�@��HM������b�2:���-4��?���:�p���K&�ޯz�jH	o|AR�)H�f��dPb��G�T1�S1�G��I�℥��#�ء˛7�
�C0�GbYd$,/<��˕`0������q���[w����Ο�I"XƘ$� `+�a�x�\{$� @��Ɩ��H�b���,�j�g��I�o7���/e7��؊;�PD����Ս��Dɖ - S�)'bo_1V7�<y��4�p�E�$m��\&���aҪ��$�[z������)y�0�R�Y�ݻ���o愴>���)JIB Y���T�]�5⾤�ly1��F��W۟�6�ū��'���}�阜��F1T�\�u��z�Tow��v�<��m�z��z���;��V�\ůmr�J��7��c�j�<����t�ޓ/^���#QS��6��2�Ѥ� i+
� bę%��F�����8(!��98���� �z����}��3!&�~���+��Hb����͓qI0	]��ʷX�,�VL�6�M�aP���w��j�Dѐ���'��+4(	FHbЂ�łǔ�(.�((q��q��d�/h#5�$�F�]�D�F��t� ���L�8���f�y�XReY��P"H�<�ad��L!�-�G�x��,	R�T~��,�*�F��C2CʐSS���2	��H����LJzHE �Z$,Wr�*�$4�E慁G��\��H�	�W�-X� �(-���$� ��b{-dh�O�8��$I]G�?��b���f���&51`���(Af�+E��;%p�dZH����w�u�K��8ߋ�P!�b�Ä++�hs�i!`�1B�7���i= V��>�T��z�Y�,�xL�r�e�$��3 
Z#k��y�B�h;��L�dM�;yq��q���!�0`��&`>�\�	
�����������C���w�iqj�Xq�Ĥ�-�ɲh�%�(.)eG#���62id��.Y�XF1]��B�.N8�SH�,0h�76IV��K����E!�~e) �4ZL�8�`u����.�m�zqX�hm^�|n�O������^�Y:n,������a�h�$���]E~�xGf@B�T���mIk��R/8#@�F�G*�FfEc�^��dl=z$;>^��ͩ�1�n�H�&��D3̊x����4��")��f�q�JA2�M뉍O�HN a,G���-�!� ����b#e\�ٜ�!��`��)���+-��;�~��p�;P���0
��f0�@r���W
���b�I*�F;eIlX;��G	H�fF��"��]@�!����#����Y}R!Y��	U.2Y��|@�/݁f�4y�R���\��AI&u�5-s�2@)������GE�2��+����-�ι�'.>�2�qd���w/b�==ݼ�����"�{�g�*~\7]�|�Ng��`�\/]�]�����7�}>��M�U�.���ܱ���P���՝w�}��Ç���,�s2���/^B}*s8j��$���e�*���`ޜ���t�V�b* �$#_��~���qSL��g�V��H<s�<[�$L�߿���c��%Q-LJ��	#��?�i��e�D�(H�{��q}>�g����#>��DR��w��E#).;�5ږ8;����[�J��_��'����J/�@8s��8���۲Z��3rԚN��3Կ��.f�-a�|њ��f�V�	�������'���Ec����~es�]�&Ƶ~1��w�R�� 5fv�i|qx	KU(
�x��+f�TM �����-��(W��F^�e
�!���i���~�+�k�WS�ߌ�!�I�ݝK�n�|w���wn�l��[�L�O���U��!W���[��c�O�λ��Q��j�~�_����ŭ�z9<������og�����h�j��G��gG��;�.]�y��V����N��|C���[�(a�!�3Ѕ��������1 CT^[C�$���ś�����\�qH�)Y��$uUi.�8�"$q��L[6l��m��k��,�-�w��8�l���@j������Y�b�Q��d��ā��ܿe(3��'���|yXy����/9�ꦅOg����t��_<W՚u��޼{�Τ4i5�͈�,��������]��W^ih���.�qvX[23���4�����3���!�&1IC ��k �ӊ�`!e���.�CMޏ;.\�7�V�~�z�+���Z����������n�ؽzc{s��l�*ͭ��`ܻ\nl���j�������G�����y�eG�?|��x������]�vϛ����e�|�:4�[o���_d^��ݖ)�؄:^�)1 dfI�,� 	f�����&�O�l��V2
35���xH�i�I�p6��i,1'$2�Yn�Xa"�Q(�2�������G��=<z���7�7�]3����|��ի�/�q��,��Xq_��TW��s�et� J���#V��p�VyV�t���v����߼��ş��nN��/+��4y����[ǣ����l�vk�7j{���n{��Y��Am3��̆��r�l0���^������O��i�nuŢ-Ha=.�ʦ�3�0&!-�P0�)u])R��I�;bȬ�u,U�$��U�v��1�R`�;%�:�ԗnA�`7��k�vî�F��ܻ|iwgGMZ�4TՕ�:��ܰ�*r�O�?}�l<�y��������;��Z}:_�ɵO*&�b�H��]��'u)6	�#5� F@���B&iM�!Ӓ0 1	Ȓ���1��1S��ڇ��$�$71$�����+�H08c#O�+q�Ϛ�J���M���ؠ>sU�WW��m?�U;}X˥��8������`\��+~�`�k[h{5Y���V�Y�4���4y�|�Fꎉ����洌�"<�t�)9QYה!ah! Hɥ�Z,���I��) YhRe X,�ä�*1�=����Ii�y��`�
����̀G�,:�M~�mat�*�0�=��(M�Z���ض�v/Ǣgj\���,�q<B%�+�iն5�e�	���׶�eaӨ��l8��nJ�Se�).���zj� [�
�ːɓJAʋ2��$�T@")�� n��,�ȎO�a�eV(��$N2�R6� �f�ij�D���,�����س��A�o�������4��L��|9}�7�a��@0��f+�%��Lct��[��t�g�ްyx�ڔV��Ф�`�*3j�h��BC$��R�#N�:�^@&F 	1}��s ���4eO< �eO��:��[0C)4̛���N��чO��k�r�HI�WbxT��D�@y+�Ҽ�rL������l��-�X��8��a�jݶ�ň�Z4�kzg�6׶K�e`;��V<c�9V#4����"������	C�P.e2JK
&E���INJyѤ� � (Y���a�`M�Il��ɼ`��d!� �*�y��Z�I�R�I��QR�����W/g�N�}i�;�v	^43	�7�d@\��~VrM�|���[-.9����-ݗ]�s�q+��m    IDATV�2���� P�@���o�k�d�%K�^cCJJ�����O2��o���'�2�������rCA�>I|��Ѩ	(�!(Zv�.2l:�oy�s�?>-}#��F�y�#V�����%�~�Dlk�X�
������������(��u��~��5���Q��K�b�T�r��y�`�T �B�@�1~hD6��pP5�`):�HdNCI��� nbl!��*`7YdT����� �؜>���9+B,�Mn޼��b�YFh��S��8�a9C�Jyd�~�9/������ѣ��/��m�T28~qr�|8:u�&q'����?�5�˪m@�p;����c�}�3~ћֶN���\ٽ�u��S�����wnvg>�lҲ˭S�="~>�j��ܰ�I�hg�F���g
��A��6���ia4�� ���"IQ�&N8����02dzlg�I�p��!d���#eC�е����/$���Ќ5}� ����bEX�R��]~%B��N�zb7���<�����5�4�@��{?K!��Q��
^��ra�:�1�aXY����&�Hd!XtA�`Ȍa (�W
|@�3�8�����sp���A�����f]�aR0k ��ZA����^
Z�+O�`�`��&��	���$��c��e��0��2���d��(/���FHI �[q2&1��(����9�Ȓ�8<hh م�@ʒx�G�u�r���gYܺ�F�E)1�`��I��J�i=�G��.3�.��r�kG���%9-��]��@���LB ]�����|�9ċ�6-��ŇZ
�RxRJ�t/ny,�	���9u���Q�2J%X�,����LjfOa�`�	8	��Y�����z��3WnJ�E���Rq�B"S4�����,T�s�Q�!U-|����$�`���8�3�5�?�Bk���I����#h䑜d�
�Q��!G0x�ئ$�L�A��0�u�r�`.`Pf^��

"�I/� �Gȷ�-� ��b����$���0M�-�eK��tis��mw�lt��֫Oε���ə��(c՝��a־w���T���yQ�m�R��1#��<�	ef��&22�˂-$��7h1l���|`�K��671+�8�!Df3���.eG��;w\�I0���=��n$<���ٔh�:_Y�!�Nv��'0����\!�7%��5b4 0��� ݮ��Ҝ(�\�v6n^߲���W�Nkg��nZJ��0��ϚZ��)��x�x�[$�R�0�#�J�&�̅�d.0b�X��	�L�L-�+`Y��x"����^�C����|��������a�k���~�������Lo6V*.ح�9�J��X� �
�dKa�J�_O�L��"U���	��˓��^ks�30�t^}fh�m��Pp��}t�b𤰸�ԏQ�J�G�h�N8�&��ٰ��M��jXn�6�[�ew>�0��UG�iuZ�G�r͒]�Ӛ��s>��N|vr�������[��W-�q��?0[�Wv����^�$C��&\VR�PB����Lj������\�av�R�=x��eLya���h�"�E�<T �W_}�p?z�H*&��+-\Y�4���OI�%d����ƣa�<yz��m'$:͝����N�ݘ�=>w���L�ת��xaT��k���������Q�]ʢ��D���vn4�W�tz����i��N�	�k����(�.�#@���H�t-���"<*��	鮐��c�k��M7s��٤$�G��A/��ϲ9�𘈓���P�(7���ּ� ts���r�z��w'�/�~�{�|x�ݻwn����N;6{Og����'��.�1~q߲1�e�����r:����t�h�lLk�*W�֙�������,��~~2^t���2��7��z�}����~���W�=}�k�mLaI/`k�ES6����Rb��(W�_ ��$v`"0xL3J�%��IbI�W�F��� ��{�P�<�����}�D�ҟ}���?��7��OI���f	�c!=�B���W�>x��+ׯܺ�I��8��_���l������|�&�_>���lŋB˭��[f =���.���i�T��?s��ڪ	G�0�Fu6���4.����������m򽭭y�y��e͓vŸH}[�^Vk-}�B�A/��
�ʴ�AY�9�B��?���JZgm+U ums����%>��X� �1���°aJ��&gנ_Ĵ0Ec�
�:j��[���K;��\�ռ�����t�.w�.W�h�iq=�����mr����Eܾ�)�I���e��qnr����|�n_����������ӯ��O<^==o>̏�ˣ��Q9_8h�r��J�h�=�����t>�W��4�da�i�i@�tW�!�  �T���H
 ������<���z9��}��^WЫ��a�������"���L�̱��?��Ͽ��>p~vb��|jõ�^������������_� �٫Wͅ_؝���#�p��EM���W}LѨ3~oh�doV6�[evq�U;��^.߮T�^�.V�Q}�������髇?���ٿ��;{/nn��j�Tj7��s:P�󋪚�񓞱f�����j���OtP��cvwk�-b�7�%}o	z	���e�^:!���wƲ$ �:'O�G7�C	�رey$(%,_�O�::��ɴ��[�E�K�o���Z}ow�ڕ�����~��h�$:�F���m��^��F��ϢM����I���8u����g�ޞ���O��?�l5��:��fG�pR����������8hQs9�����l[Q-�b�p�J)/h}�ߴ��J���=nh���P:�����`	I_4�Դ��e�I����fF���#@��gpxo�#�o>�g�D=;���$d�����ק�,�����r�����~׵��޹��,�I��w�����-ӏ����#k��)��pzrd�s|����^|�}���|�>;.g����|^~6.5m�h��PF�ެ:#�]��N���Ĝ�4��*~Β�i�ʚ�ʸF�2�G�+IH�P<��i�ɧ�<2��X�P�!�g���9�-d���qN�� @����H���Ǩ��)�d66�bH��+�搚��%/����NQ�H7�i7��F�U/m�ۗ���Ǫ�IY�N�?j�:��[����χ�\�H|y2p�Pk��]Xf���ә���܆B�f�B7����!�Z�$T*u��}�Y�.A��� ?�S-ѵ�.�p�K5J1�~mI0��6Z�vZ�m�"�����"�BV���Ă��Fl��POd���N���R��.�̚cq6�
��9uVoU���f���*�^��F�ߙl��։[6b���xɪ씕�Ry�ɬ�W�g�ա�بx���ۍ��x�oC��b\��1���~sh�ZHh����~N-X`mCjR�
KJ��� )�	�G5������r�v�/�$�I�}`��?|`R 清{�1y��#��V���w�)�����(�A�J��n�bZl8p��4��m��5��7���n��ם�OK#�Aԫ�U�}��cC��hu�T����h�|g��h�\s�u\�`�b�#��x���|��I�e|q@��	�#u�ML40i*5�J���Y$1Q�u>�`��`�Q&��5��#���@��_')����:�~����Q�{��E�Ϸ�u�eWZY"3�iO9F����s��id�8c�fi��jW�ǝ5��M+�ќ���`���F�Kۯl��v̑���G�1��a"�xgh}�dÞd�Nb�S6�)Z1��äw����C&iüv{�X ��i%x��2&���㥖v���=�K�Sַ�/}��� �@ٱ/xD�++N�hY�?5<9yz����Sf<pD>����.ĪU|T޸~y9�حG��E��v1�QI�����V�ԫ�,E\R�=�<X���������t>Yu[��W�Y���v,_�-���N���Վ��f�8�,E�T��F}����9�3�P������0��6M*�m�4�,I��=V�\i���$��t��	����g�;�n���o�ץay��ʍ�X�m!�ޮ�0At>�^�V'�����u�����૯�Ӌ��x:9���?�:�z�ʵe'�m/k~�{�ɹKu�闒x���O^�ƶ���fpp�p��7���w���k�M��׻v��Q�v�_�l�!��"ΑWf�e}��7��6q�q���b��9�[q�2S�
�Z�A���Ҟ��P,yc[@���h�6{���I���x�R�,�3)��J.���~��T��~�g�QD�Bf7��0��i���Ԫ��,z��}h�{䋋$f1�hV�j��>��C�I�\���:���A%�%;�0&�6a��*���k�r�Q��7j���Sz�|�(�?�t�zL�]?R6M!5��%��3�W�d�FC�ceD/��$�0�� q�EfLֲ�� ����^���S�u���v�ї4H��h��bMI��F���HE���Ǹh]zj!���I�3�I�$�٣v�Py1��Tq�:s�$=$%�bH�R���I�dH��81� k$K�Ou��R���� �M<��.j?��s����S���L��o�}�/�F���>���9�-[�kq��!ܪlrԋ�O.��=�հ��ey�O�Ko��Sr:g :�����&S�-z��lj��Җ�F���P����x��1���i�m��:�
��5E_��1q�PTk�*B��,0`�$�c�'|���̮"��#C/A�ϼ0z�W?��Ѝ���c��;o��Z�a��ܴi�X9Eg���K�1�<jq��U<���1Tp���#�����q~�����ㆦz�����io��7�M��D�BZC,(P@�2�!�n��)��1a�D�� NeŅ:�ۀ�0r�<�1�tixd�0��g��m]wo��0yR���xh��&=���	��4����[���No�t:�j������E����]1���@f�)n��͞`(�05B� o@H 9��r��
R.���р���%)W(���!k�Sy��7��rMJ�O�����4V����Ƀ�Έ��-��h�74��钶���.�5��kb�[��C|�/�`�b>l���@Y��˲+�m�����
5sf���Z?6n�>;^L��6�.�;��3����W�Y��a,����U�.� �Ǭ_&�!�̒� 3IZ�B���$��`HvβX �������mfLآgO zp���:�]�P#���(�	�X� @�R���ӳ
��n8�GvG���QF�$�)���g��F�@��}�Nz��x:�t��[ŉ�9H_�ڞ�W��B���մ�~$;�0Ml��+��
d}U[,1S:�,z��F��~�1;��g�嵳��7�Ѫ�;�;X˪��t<4�ܴ�ׯ_�x~��_°;g��ެt����z���%P���=;�V��$L3z��Դ��(�OG���}�Xa�2ɰ�D��$��y��>��S�:����a|9�i��~��˛��*ɱʚ�V��i*�T0u����<�Ą����X��烋ɭ{����[��t�ܺs��Q��_����M%��-�^�a+�8���1��e�/f�S^`z%VwWW���f�U��z�����j��jy�o�zǪ��4�~�����=�������" u�@R�#}=�3�$��O:6�޹s�c0b�0O�(�`�
eX]��_m�������T~B;<�2�ͫ{�����G��{�v��$�btq|��������ppq�(�9�lU�X����0�Uc���g_M��[ǌd�����D�u�\̭K�/f������ϗ���X^�����Ѹ�|0�+ \�φ�ͮ��o��(�(��_��6�@�ƣMQ�Ap]]*�
�E�Di�yZ#M�#� �z;I�������ث��ݻ�~e	�G�L 2����?���u��V�����|]㾰��yyw�޽{���W��1�,��b8r���8��4R��(�+ضoUC�bW�=�?���qIT��밁
��{u_W���ָf��k	�ů��ߏ��N�����t<q��t<�zf�s�ޮ7��?z����ث5.TT�dp��wt~:Xi�P8_"# ���R_H;�&���>��I/	�U�U��I\޼r�	n0
B �S���:�/*!n���=
f���5V�vu�Q�w���>x��G����o�^kn�C\�������*�x:�k�̋�����s���."_��,~�w�������fe�ھ�ں�z�{���no��Q�?ٹ߼����p�R?1�3��鷴�5��e�5Z12�j�6YV�c�%S�tZ�R�:�*;xddik3��� ��ׁݤƉ&�YҀ�X���]<�3Q���jS�ܐ�h ɓ,��j���������o~��dq�[�������QZ֦����_|��������>��ݺ8:�9A�E��a�ץx��̉�,W]�W�:�Qf�u,޶����ʵ�]\��v{�����[���֍����gÙ�畧Ç��������n�����������n����4vZ��*w\l�����ðP�hnL��4z�������p��.�����ә�!�&N }2M
�D�d�zbx�j$�Y��@`4����ao01���Rd�nll�[�:�@�~�����Ļ��v������KW�Hps��_)=�K��������Z�V���8+��햺;7��zq�t6�/�ZN ��W�<:~�򉩟���Š\���a���K��֎���C��t���^x� �e�^���`$.D(fN�_O=�j�P$�LZ ���X�9�� aTMvG8���F���ѣV ���=	`�"�@r�d:�3�o?�b�֎�������e4�':��]-[����=��w>ػ~�����r����ջ{�&*����r�)Ff�<ML̠Mʫ����4;���nM�_��������d~:^�N��.�M���ݜ9�l�[w�.����4��!��3�_���8O+s�r
/�oNh��2� ���X�_7�||ۀ��P�̀�,�$7�0���H���#@�d�A^n	�b����\L���G�m����c�q��]��me�x���˻�/�Z���]�|�'��ȹ����ޜ��'��k�F&!磓���=��9�XLG���`>��x9j�7<v_L�t��ݤr2�+���,��6�]:ٮ�g~յ*�^bҠ�[���)]4Y�ڇ[R��ޛ2�OJ�2JM�e�$�̈�$�dI�#$R���48z� ���E(Gm C�����%��j�n=�jl�֚��1�0-ީ����;W6o]ݼre��m�Z�ޮr�Z�ed٨5u�\�.���|�j#˳��_<?y|P>�N����5��V��r�rӂ),M*&�t &rM�ĸNWg,m��чĺ�9��W�&�k��&������'��["^���L�8��S�˃�!2 �E ���3zl�R�$�M�Ru�Z�~���}�L�s���?-�\�@��[7uz{P*k1��vW�;�X�\��ٹ��*J+@Fw@��C7����_�^L���lCY>5�-�ڥW��e,\LJ�ܝ�M�ck��J[�o��ԡ�H]E��6�N�1q��	!~1�/�(X ")�Ik��^990KQLX,�P�$�@���Ӓi^̓@�Y�$�h�	#x!��\����7;�f�w$;$��]i�f5�`�O�����2�n����-І3�X���~5ֹ%x�E�i,=;���ۜ,*���ڜ�;�js���NІ;��{�+��hQ���c�8���>�5�����)�Gx��oB6pxM��$R,Wfç�`��Q 	˅?��`��}N��'��VH!ϵ���g��r�Jl�9>}����'���?�p�`0�z�m�.�e�̷-���uwɚB�p7�MZ%��caD��N�g�����g'/>z�9o}��Ry�����|5=>xq�k���I��y~8t���k{��(�
�;����:�&=\	�R�{��5��⃷8i��&ݞ<y⫍���8f��	���Wԥ��J2]Z2���2	}�$�*�j�gF�P2�$4����gML�d]ح�26�P!�$���Мy7/=�׎��W���/N��'Ϟ_>?fuƞ    IDAT~�`2<�z�����dǍ4uחƯ9h�����Ū<�T������t��ى����l_�K��;K����������W'��5�q��ݻ__۹s��S[mw�j��5�ꨯG����׉�X�q�B�V[�`F�ag�A&�ЧY� 0���y38��R�>ۅG�/}�@H4Br���Ș�gvٍIb��S]^ݼђfl��%���g�ޭ���2��u�Ƒ���(��&/�-d��v��rZ�E'��X-'z��w��\T���#MJ����9���R7�_@��Yl�2L���J�m��΍����T��[���� �g�A��qm��p�$R.BfQehXM6�5ϴX��N�9C����'[�,C�Z\��)A"ɜL�f-�C&�h��f�F^��G��x�>���`�juS�$'�B����R<l�&/��L�$qJ��
E�o�؋�� �aЀ	����Y��V��>�֥��n�@���k&�S_�&F���-��b4�	�x]��4Žu��5�����a|�����^3+>�=p畍��j�l)��H��竁������z�ڊe��I��n�
l�$�j:��D2ե�py�P��R͇�_@1�2��F�*�⢦h�.H4`R_�H���x��f	���LE�*��K�ݺ��	"@�$E�d�KJ8�(�DR�ejV89H�%CV�\h�^�����應)]*��/z�α�ʏpM��}��+d,d���j�x�����m��y�J� [��N"[�qv��i��*������'�Y�F����c�A��O�8�b騐*^�LD-���� �RtTn:d\868��&�!�uvy�	b�R*&�.�s2�$�:Kf��T &����8{�OH9Q������&��Ը�-~8ʚ	�6R����67:��W_?���g���������w���ED���_��|���^�AH��kZ�0�0�f�Ê����2�∌w��1]li6�������`|lZ�Q�u�u�(�$�d�xiyE.�o��߿�݊3�i������¤"'&������iC�f�pWog�ǘ[cX���7�-չ�$`��H^��X�A� �H�@�J�1��o������w�ɗ����W���;N���;�%o����DS���q�I���"(+�b��@ ���c*� z�$10J|�Y`��Uf,l�&�%f��2FH?g�̋O�X�0�$Y͏� 5�-��;�O�ڞj{����؝�Ȝ��H\d@����T|R�X��KMR�]I2�	�u�1-0�t�-��Z���O�K݆��Ⱥ�ɦ���K��PU��ybZ��6�F�o���1�45�����j����֍f�h�⺝�=k��Q�Ro�6�[;��<��)�k��.�e��I�)έ-��:��^�J� �.����<�>K�5$����h�_s@ϒRe�h9M�h��x���(��KΘ́�fƼ�N�] ڒ֋J�v8(�z$a�{R$��@L�^.��������o����M�#��R���W��ܮ�N������p�K�t�f���o^5U��8S>-�(�X[Y4��|YQO�#^�<��N�[���\eK��W}w.導k<� �V`X� xqQ��>�$q
���������M=2�Gu0h�4�E��.ȕ.��W_������"�66����o���;w��^�lLͳ�_�x8<��Ւ��q������w����ol3�"5�6,���`��V�����5>�:M��ݵݞ�B����������];���ʙ��}�����>Ǝ_�����e`����n�
��c�(K5�3�8��2JN�?�&� Y9-��*�;�9�� ��-J�,#U���j�J�x[j9yb�Z�eQ�ae�*�����Q�/�8����������}��FoSS9�O������rf|ۓ"45�}Z��4�������k���݊��N&Ϗ����Pf�����ݻr٧��/���%w����������G/*����N����HΏ_=z�3��b���+�V}�Vm��B|�����bx��	ю.���\�)�|����U䵝�DC��R^�x��d�^�.�����!Վ��y�Z��i��Fi��p�߼w�Ƨ���n�s�W�� �??4��:o��x��jt67�l�uHE��LQ��x�4Zg��pW�͍z�an��wݡP����s��?�<�����_�i��{�z�ʹt0�N��n����qQ��[(F�b)�+z �|̮��PL�0$S��|�#y4�
�ȅ2y���k��#��̋��d��G-���ق����s�)/A�I&\+Ë�Wz�����|z�ݏ�q�Z���z~vp��I�
�+���rQ�z��(�O�:,���
�
�jο���	Um�!anoy��~��(�{��;�ǃ���l��^�E�ۣϯ�Xv~X�lw�l6�n���k��e:؉­%��Kn���[�ʢ������ׯ�E՗��U6� �pe��N:~]r=�~Ϟ������	�ZH�Wi7�e=v�J� �&�{�=7�ĸ	h�Yq ��������;q�ׯU&��N�yy���[���;w�����N�TWǯ�����u1aTr���>xxQ\)ANoH�R���+m7lW����N��w�]���������~u���j��>�����l�r|�$�_��� �����3C>���J�Ҟݨ��z_�-���7�,�p3jr0��11bm<�S��&`!M!�\ٽCz�@�l�=fq��kz���Or!v��:�-�:����rnI�e�{��v��Z�t)���o^�ؽy��O�w�}��Wt)��,8�� ���y���/~�Q=�A	;&��[㴃�@�e)xU�����~���|`���>{�ŗ����ˏF��ά����,*��<lw6���ʹ�x+8F�9{����
�t���.o+�O�{�D�;ASY-+B� s��ziR�$��v4���ӫ�RיQj�ZI��9�ҏʫ��u_���Lj(�[��u��1�V���[n߹���~�C_P���1[�nn�p3�D��7�Z�U�h����+�z�Ӛ����(_���/���˗�z����w/���V������q����y��;��)��jq��e���H��������.�CA��S}~�.�`�ai�4>ʷ��X��S,�3� ���c�� ��c
 �Y�^�Yov.-���5s>w7{3Nf���{˳�V�SYݸ�}w璛 Z~��r��N��k�Tk���nu�v��f�lbs1��R�L灢:O��^|~q8X������W����K}����dR�kN��[ƈ[���n1�^:�/�/�������ͤF�-���2�+��F[+��$�0�!$Y�?(��!� BA��;����Y}�� ��2��$�(���$$��^o��%�s��W���=�}Tj;|�;f��r�U}���;;��3[�����7w���1~�[d�͔M[���G7���lz���+M*���<xz��tpZ;84��M����+?VS��_L�U]w��Xڛ9�m���"�.��i�8UI���ၩ�1^�6u�>M�� ��i�����h��2�r�����ijd�0i�x�&d�ed�d"F��h�}��'%�|lsۘ�f�j՗�z�������魚�;�^k�s��)�\�m��n������.Os�[6g�b�����~::���O��F�G�ǯF�����Ѩ��*�cW���vq;�-g������@�u:��&��T'_wi� (��4��ƀ�A�CS�>	���2i2U,���ǆ�j5��������os4�G�8ŀ���!���O-�jϞ��v��2E�rK���%?�����f�֔���߻�ѫ�ƃ�1sya�'���>�3�6F5���,ݶ9��β7yy^kt_z)�6�� �F�'��n4;��ˍ^���ūW�;ׯՇ[n�*o�{���I=C]�jddi�:,���\T��/�l�Ԅ�]��Ջ��P�dO'D�\,/<æ�ed:�Fg�W-�ci��L�_܎i�����b4�����wtH��d���g'��_~���>����h|��aik5���7�Z�xo����ƴ�42����~k�ewk�U�O\U�a�Z���e�ح=S�,�������lY'�.�:��d�`5�{rxع{�������������^�z���[�Y���Kc�֦�������(��|�}��jE7�,�c�kgF�b4��-���L@�Y�i䷉��.H�i��.�R��w!���l12v�Q���ql,��[���wR�4m��5.�<N��7���n�7��h)R��O�\���V�aL0y���Sӊᅽ�1�K]��<$	y�rH�`I�!��N�Ӆ�vKL�����3���ԴIZl��gϴIz)X`�T�8����!������ni�4)X�K�K�G.y{���HW��PB&et1B����$� ��6Y�CTV��.�ǻ��b��Wy(b�P�E����|��.Jk��5�)�}��R-�P�(������&`�oa4�@����Tjd�Z��2K,��ZC�*��yLI�&,c�{Lzr�$J��C�r�mՔ(�I�n�Z�~0��&9�`�8����%�)Ug�M�ڗ꺣�Wl+n}0�^�|K�yI��$����3Xu6���f��F��J�Ë���瓡Պ���g��7t�� rX��)�,�c�����l����jN����I^��S��V���]�k��r��Q�▚�k��*3bi��pѴ�8+Z��� ��!lQ�h Yk�����Y�����[�kQ��2�x��cXjי��u3w&Ya6�s[i�q�fq4|���6�2v�m��:r��	+����ͫ��2�{���֎��@�:V�]0�7=z�����6��x(Y�#�i-�Q�M�I�Dz��G*�Y��"H ���J����E$ �(��Q
�tiEC�I�@2��Ԍ=F��9��D�	��"<Р��ty���Z����>�ݱM�8\,��n���}�ltn��7�&�C�t��US�ј����������+��H[´c�2���+�:88 'ي^kef>=GRz��o�Z�7����$���C�1��1��I���}ȜW��q�2�֣���6M�����ZqVIue��i.�^�pd����|w{�M���J[ىgu��}-���*��DN�9�}V�X|��/�x������`���m�U��N.��������2ˋ�[�)8������c"I"$<$���
Ȍ���!�:b4b2��h �,F$�+VJa p�b|M㰃�˽����2�'U�?T�lB�+t-z�Bn,��TE�ܩ�Ԑ�	���9���egC'��ʫ��Fq��f�߮YC��Ok3�#6���U�6|����b�8��4C%*K�+?�^V[��3}S󀗪��}�q��r�^�jn�m�;�ڭΦ9�fl裂a7/���9"�01��|L�-���^���h6�f}���3<k0�BRYv��,�l�b𔑹��m�˘[{�Bdg-S�! �rq��`mU��YÖ++gژ���/#�]��� N�+�몔$�q�۬{%
���XXR.I��o��o|�4�jV�����'�wn���ul�@�������hL x�Do�R�PT��,���Y%jz>fͧ�n��Wl�E;��~"���W��ۚ;so�em8�n��OsB4|39`16ɂ�IK�?|A�/-F� ����KN�Kb�\M�)������c�̣� 	��Z��/��y���,.�5���π�Ν[?����#�>��MN/_O_^�>+-��u��]�=]��q�hqq^0�V�c�x�I��X��Q8�g,of��oy��\��W/�����f�����:��7?�Of���yk��o��}ŋ�G/�,��pu!-;p'���OwIk�vi[��El�{�8���P�0��.r��i�4�$HY ��>i��zjݺ�����@. �P�ć�����7,,.|*J���WC�~y���[���ڋB�燇/���3ϻ�aq���"�S�j�7cV� {���7uh�����϶[�m�jh_zct~6ho�.F����ަ�P��oTzW����褻9�n����[;_�8�}��\��7K�/�ߌ.*/�L96/�������ijq��P����E0/o��~V#�o��ыY(�Pz�0�FC�Ȍ3{rC
��pB֚r1dLA�(^-^.q��x9]���^��Ѯ��������{�|�;Wn�nm�����h<|>�v���L2�g���&��s�*#j�L��7�- �*kNrf����b�[�Ӟ���������*6nT�g��[Y�n���ާG������+/.w������rWJ�s?>k["myEh�3�t3����xd�0k��JM�4�T@���C�̅	@*3B�uu�b��.E�Beς�|����~��ѯ��?����W����T�ի����~��_���߹{���*n�R��_b�s����nD[�ep�U�$����D�ʍ��U켰i��hz���6�����w��ܪ����<y�������m~�Y�x8|�~�b>;}�������;����^@]�
��w���<���&�siG���V�G�s�Ê�B�%��!����jV�����p�û�n��*ԁB���#K���"+������̗/_��퍵��/..Wn��7��������'�^r������ti�����q����;�O��J�G��"A�v�'!h��W�$�'�����.I��0��5����RÃ��i�f��&S�Z�͝K�P�m~�י�^x�7�6�-/xt���w0�Z2<��]�+�e\�?)u�j07V�ʨ�#�%�ʶ�t�^�-��{!i}��zدhn���]xw�r�[j���~����p������3ڥ6]"�N�6U�犗�\ZxƏ��*f8AK`�Џ6ߩ�6r� 	����@~��9?�}���O��T¹L�X�`��%��@U��,Z�Ăw�G�(�>�,Ezp���腫w_޼v�����T�qZm��Pl�@}��� u�����dߘSE- *6��67�)���l՝�Jm�Z]�\�=[>���fejg����~��o���I����/����h/=��:��!f�$�uE�"��-�tӃ�j\5Js4Y�>��&S�*f��p�������;��(�&�� $��%J�.3)� BGf
��|`�Ny�D�z�]����ss�/�y~s�ڹ���A��-�>A��4�Vg1*CQ�C[�zlJ�,�������Lm<՟^�9�9�z��Y�\���x�7����>��6WԬ��g����l+9g���ʮ&;M�xH�u�U���xb�hw`#��?O��� ~r��/�"�L��O����9���,?%7�*+'_!��'�� x��R$�ۇ2G�k��i�!�f����R���:; s�L>�-�^t(�V�n[]�8g�����Bӹ���2�Nj>c���2�Wk�f�2�T�~�>vD�߸�[[����䫝���g�Nmiﴼ;�t�qgܧ�A�oFpgM�鿸B�b�9HHlh�FM�i�_��-	�L8� �N gO&�X?����J�J�	&�l�A��&i�G�ڋVN�p�Sqx��|;Tf2˨����s��[W[�.x������K�Ջ�1~�}tsZ���@f�28�^��+����~����L/_y�;<z:�<�}v�so�;����n�����n�Z�p�n�L<�K�*��[��Y�X<�I��D����90�&�L��v �<�GS����,9 ��LR8�&z3C�'��`2��������D	�
�Ў,��y�C?��3g��9���|���d�9�z����X\�����v�j�Rǒ�5ו�7c���O��6Ӣ=e�3��K������vУq|�ٗ���ן�������';�r�W?j֟tz{�3c�<�����օ
Q�۫���9��GӴZ�������v����ͷ�-$���'&��F��Ο� �)�'�3d�O��^x��ņ=����G��͡�5qA�{&�^��w��(?~fQ�    IDAT���J0w�j.�6Vf��2^ۺp�⺂D��|Vf���[[�u�0$�!�9��9?��t�/���:�6g�U��w�-g���hJ��([�����ֲ�}��w������*|�Z�=Y�Mæ#�����E����J
7���,�Ξ���V~9��'q���?��g�A"��Dl �'!�I�2�Bl�Y~��܄��gz4Ń>��kD6�Svbe����O���<�}�����������!EߙY�9��ɘ.���t~���Z��Q_[��hmf�彂��s��.TK����ز�w��}���N�T��n�s��Ϛ������}p��ݣ�J�ݓ�W���� g�;�˥{W��s��7ז��gs�,���z&.�´��Y,W)v�	����������%�O_���x�r���B��B� -�̭��v�����P/�����Y��8d�d�J�E��P:t7!�*�M�);��9�d�xn�:���^��Gjw6X]l���K���V^^X��Cw���kÓ�A�hwߖf����(�����S�e"�<s�?�� gg��@��
��i�AQUw*
}�����q��g�DK�
Z�4A��u� j�� DZ_�R�8� �-�O�@N����K;�ĭ�2��f����`$TC~5�SVb�+�}�@�b�RĐe�o5ݩ�L���,s��a�]%�=��l�D�=����S�o	F��Vm�R���UJ$PTR�̅+Qv� y��4�H��Ɋ��3�Lf�3CuȲD�YB!��B|�"P�*�����(!����$%%!Fm?�S ��8td����g���V��ٺ�*�*뀳�%5�P�1O���/qޏj����
K@TYc��}�\��9�����g��p�y����4�� Ψy�8FBzN'튨�X�I�!s���-\27<��ሻ�R����O�?V�V�d��i����A0������s�l$��
�Md
�W��2P��p�yID!B	30��
`"��~�;ǆ.�
�$�N�gj.U�gún9v
o�S;�o�5�4ӝ�M�����J~pr4������N�-��w#�VBc���� 2+���Ԏ�~B���6/1(�E$r&M֨DO�T�A~ Q�8��3Iq½��$��B����p~N\VLQ� l��SB��r�$=����)gQ��C9�ʁ�*ěc�d����A�ùY�>ή.1e����ȿt0�>�ܝ�a�yG��\�ckj��?����<='<�׿�����{�ԟ{��! rxk	5�F��gJv �z�T.�0o����\iq���{TBfK+rie�V��HeIC�'XR��e�z
R7�Y�1EKN.+�pcP�~:�UaRn�(Wԃ�Rs2^�w'����x�u�LB�����j�����h,h�&��v]��C�Ȯ������Jkvuye�13���>8���$���7�-N�Z��t��U�O�I��/
䊎b��@߄��&� 6�R$�eO�&����U�"� 9�,N���ׯ�0�q$�ou�NaPdF>0%�~�\�++����+�Z)�j ��M�)R*�Y���.Ġ �$�L�-�cا[�Ly����l/y����I���E6�d��@��A]�2R�D'��y��X3���O��;�^�9㌧~Ҝ���/�<�nJ�;5gv.O={�t�hie�T��!G,�88EFB��\	fωr}S� 5!�X!�'N|�i���qQ 89�B3�$��$�V�cHe)H)9`����� F�u�
˟���lu���srӻ��e.�����
��$�G`�]�&P�܌�̃2,7�:${�������fenuek��Z��Krs�����,ʌ�����S���vS?&VcEp�vDn7��l��m���{O�zp2<�;�-�N�^"�w=�U�щ'�0��Jn<�!�I�3P�
��d�E�VI�oԤp~B !*���g����w�I��@���<ԄI���E��ܞ���w>���ι��w7�����ḿ�U�Saip�F�%z4�=3�`���y�IgL(O���5���{[2P��k��1���q����~y�:�[�֚&����i�z��[��v�u�r���N�V�vg?��o(�<y��?�;6g�Z��9��j`��|��L�D��D)�h�w9���{�����O��	N��s�/7!�j~&����3'��,��r�m�oU3׬����?x�M�D�2�v���:��QvNC�ֲ3���Bo1�[�R(re�.�xі؂1u�ClOcUW��+��hUVR�|��S{��Ym4���\xY]��,����io��oK?����lu��q�b��x�������'ӏVn���W��B��&���~eX\� $k;r����)�.�"�D:1�gҼ�D���I���|�%}����>����B8zj���A�o��j�Fy�:5_}��{ｺy�F��@����l������v�fI�*���K�D�v�g��T�Q������ ��R�r�s�P۵�9#"�*nsSOc�bEԜ]�M/.l���+/������ͯ[���Ϫ���"�t\jx�u���2��`�3���~�K���0����Q�$�D���s�g׀+\'�m�˔��� L���89(��������pk�'��x߱>�9��F��;��z���_y�<Kbn�q���*�Ӟ>�W뱞`�-�]x*0�v.�)6�H^Wt�&��Q3�{6"��wwK�����L[�+��J��|��Ƌ��Ž�������{�__���1���z����������&��M; e��38T��UL�/��<S��~�Zh~~�U�}dؗۆ��	��$ǟ?���Z�Ü_�Z�X�^��I=�	��2*{����Р2BRW�mwn_}���~��������eR!�G)��� �;N����8rc��7h�t|��;�r�П:����au�����}�Es�\k}�)q��⍭K�N�w�^�?*����������̧�}��SW�h��k'Ą�E��Q}��N;��&}5Y۵Wx�'��3(��PL�����e<� 9Q�8�jB�B��3�,K��|'�9JaB,ۢ.-�V\}(�p�����_}����l�;V�0��v�=kr��(�xC=�Ġ�b�DGv~X�%�W�N)��wwwhB7�To�m\�D|^nL�����5U~��G����w�]X+?�� }f�t��5Y���6��Iܕ�i���s��L��{��,�SJ��1�˚�>y�?i~4��I�� �+�B5�N���0���/���$�C��'�-N�V1�לb�xJ1�Ν�����o����nmm鏐��yrvz���H����iXd�����i�7+Z��a�BA�������]��n,O�V�/�ʽ�sw��ݼ|��2n��������|��G'm\�q��J�nF�C*��Zd�m¡J+�x�)�bfT�V+,�XlF4�3ޓ&y���~~9��Wрb��gBʳ�/����1
3�:p�:��Dq��z ��\5��+���s���X�~�¹s�+k���Y����KK}��'�F�ì�9QM������~�17�����Ƞ��Ҍ�kR�zc�������炙���?<�?j|�?z�!�ʓ�D���DW0i�#�1)��7e�h��'!*�uQ��%�8:� ��Arr��� ��_T�jx$��Y�@!�f0�|xጪøqïχ��3��ى��sS����K/����7/՛K旆7�볬�w�,���4�KCeAT�������0${����˴,��;53ݸ4U]��ݜ}n\�����x�7_�}}�p��=8{�s�Y� �䜁�<���� �шMG�M͖�y�	!���X�@B��9�M�H"
|���T�JB���3S���Ow�@#��)?e"���L������d��;2�b� �:�~C뮟�7f��ܜ�s�ʥk+�+��O�6&b����R�V��[��އ�,��#k^�]����G������^�p|���o�n|���w[�?>{6���u�1�+v�.��g��L9�[fc����$*ǟM�@���&�%&AN�'��� �	b�~#��OlC��Z�𫌽$�X�]ց�;� ��$̬��0:���|��4�t<�@���2W�O�.\<����Յ���E�WK�K�k�֬m��gȿǧ!�3N��� �ZԲ��S�>�7\���m���?'���}��?��}�)se�B�f}ЯF�G��p/f��-P֙��xn�I
n�8�a"5'CEJ���J���(uḨG	����$���`���R��` ��O�/P0���;���Z~ϝ��
��VEV���'�����{���O۟?���S�� lanLYĸ�FV^[�gWK��ɵ�K�o,/�[�έ�gר�U��+U/�,�Z��ݵ���NFeO��f����e��G�/��<*=��a�I}�����ۖr=f�g��G�{V���g����[��O�skL��-���[/CW\X½�W�BoZJ�C0����m�� -)��@�pI�3��C�� �/P�2sQ`d�É�[`�8-�u��|7;�)ָ�ݙ�`'}��j��W���i�s����be�b�R�|~�+ޥ��+�7�.!mj�V�V�Φqz`a������Q�耐Ϻ�Ħk'�~��������G��}~��7�o9�������3qwӍ�*�5֨����Uг�TU}��ě�����I�B2L"�K�LxQ`�J�����. ��M�gV��x2��y?�O��J�3<�B8y���(��Inƅ0o�'gN�㮳� �zp�P�j-O.��è6 ��t��~zH��?Fu���{�Q�BMs!��n6�A��'m�ʨ҅I�ҺD&HQI�ي�^�&-�I`�l�R& B�}��'&ߌ#�@UU?�+��mvq�"$3��� �p_N�")U?��3�g�)s��W?�/6j3��36����m�7�.-�L�!q��ocfi�Rki�ڜ�M253g�~:��������a��{28�Q8:�����v�G��ް�;�vF'�N����K�Q`�׳	s���r�yZ:�=\Ml�u���I�:����e�/��Ɗ��s�"H�s��!�=��(��"�[�<��
��}˓%;�P�\W�*{'�-��k��&O�8�����Ka��d�M�
�J� �r2�<�|qq�|u�^�K�o�ӹP!Ŏ�3Ø��S�~�l�)�����A��`�{< ������Y %@ڿ6�a7'�9����#�u��"��xj���:�F��!<�?i��N��KF0h�'����X�.���AH�F�p���S/�nI��6;1��:�$;��f|�L'V=�����N�CY$������`�N�5��Ks�ln�ɬfmǥ/?�zan��戋��*�5�X��:�mu�f=@D��\Y/�v4H��N Gy�5�:85TCGW��jl �V%9!��������4�e�̹�#+�2!����
�gK�%W��P!r�����8qQ�	��/�9>�QM�fVIM���j��J�-H���N� Y�E�Le��hN�/_���pq��K�Ԍk$�,FX��@��L�q��Oq"��-R�@	9!�j�,�|�$� \7% �	50����\5��|����tRq�BWV����G�h����J�qx�6�tR&k�h�6H�*ؔ�2��ɯ�`V�q���&��V6R�+L-U��.U�
��XQ�������������j<����;F_r��Bp��08ײB;��_������G�xe�99��f�MR�K���7��z����q�a�~�s�3VЎ����<aY5NV`S�&o#��@3�N�Cnb �)�QR����B��' *�yBf�~�1����B��|9�	���JAߙA��l��(�e+$	���K�=��fY�z�\��`u&��榳�\�S
�W9h���H��0�gV�V7/\\ZXn.�\�v��Ŧ�~S4���-����q�f�u�'JT%��+�W��<��=b,����u�0N{̴;�B���p��߭�\����v�U>Òڐ9��OK�j��-s.ۥE��C~a)J�n���L�$�/2��X���_2�/���Q �Tbbۗ����P�O�#�O����Q-�я~t��U��t����}W'�S}�<lK���I�<�#��|�\�4�!�u�� �/i�ü�n�rRRFVBp�����I���3�}�ey���r�lz��+95x4���[�w��i�nc�������Ù{����b�WT5DK���'V�,�ï����M�D德vO�F��Q	�<Z_@5^�����d�b9�p��O����nAa���/������ʋ�b�[��!|w|lw�k���v�
����O(�	`.�{M�BK�!�
�6Jv�YbG��M���T=�pA|0��M��:Yۨ7=�\*�n}�/Z����/�~���׃���W��`����q���h��Cm�f�O^��0>^�WCZA�,z4fN5R�ο��+c�(�v�O�0!��*�hR����I��,;7��u��	L�r܋s0]`M�aQG^3��i'W~���/���ݹ������γ�A��s4���ŕ5vSNGr,��Y�'Bwp|\!�
���ܐ�p�x c�0H��|��U����^߮��qOf��6VW�j���L��.�P��}V?��o:G۞�h:#Pf��L]\�������$��R��or�D,<h;���ϓ<����<9�3*�-0� fb�È���A2�>���W}�Ϟ����OO�M�;�zwn]xﭗ^y�E��z��{�}����w�Wc�5^eq�(�Nxk�H2K�@��tC"��q�iG�qSаQp���߮Ya�Y>t痚e��^��Tix}�[>����o.ܟn|V��ޣ坓����Q�ak~�ڥO�g��X|}�~�Zsw�<��(F�3/�.m\���fw�����:��T�b���؆؆�����P8'�p���D���2J���tr�N�
u�>K>�e��!�������޿�އoomm���'�#��63�����'�,ܣ��Рp�:U0IJ�8*�L��"0��.D6L�9��O��Kqg��n���:�8�nL�,Ξ��ϿRn���_����j�=�ۯ��G��q�j�!���bc���Vv��젥䮚6AN��Vk;$dO"
�@f�3��	����$��o1Yhz��Q���� ��L�E�b{�U1�J�{�j��~��s/<7����i{x�ow�]�V}v��₊�e�t��*+y�0v#��CKv�!',d����3��F��캧�Ύ�v�:|��Es�Y��\�r�
zy�F�d�f�����7�~?�{x:?���}�R�Z&�����B�?��l+��AD)��ݩ�H��U�7�3��X�N��b�'D���	��9i!�G�Ķ/����@_iy2O�g�Y�@����;4P��[\��iqz#��7_�����k	�]�M�째��M�Ԗ�����a�TN`��]X��3�Q�S�RF5�F���ӳ�'�i��Ͷ�\.�����_*��Ow���O?�<�y��a׫��74C��Pq����g�͙����!ƵPOh5��'��|�	QB@&0�� �ρ�^�.��M%A��#��pI&N�� �
74�s�4�qG�����/���Ck��W�!iB@l]?Q\ſ�x��_�cJ�b	�7�2�{���rJQĜ�ǫ���}����K��X�R}�ui�Jm�{���w�~V�x��x<;����t�̸m���V&DY�5`qA�a"E��r@"6�0��@�VbP�#��`04
�Q��Ȕ�O�%$i^�$��˓N`0B�c-�d5���	�e���C��fc<3_\h\�:����o�~wq��VV���^���z�$�h5}<�D�ּ��Ih����\�J�atJV�,�Qgzє0�Z�[k�Vn�=_z����_�z��o�h��̃'S�ز�͔Ξ��r�x����ِRZ�7L&��5ƫ!A-6n��D�rbӁ��5�L� ����    IDAT�dB!��'`~Q x�$C`�'�ϕ<�^*y��RL|�# qil`R��s}��0x֚�ͭ�w޾y�v��y3>����}$��C��ڋw������������kNgO���<ЙӍ�0.~|:{���&�;�p���~l�����Aw\y|X9zY�D ʸCR26�ςajH�e?�r&H��(۞�+*�#JHT�p�j)D��"A&���=��klnn2?�kǍ�Axf��)�WՖD����������?����V+���������L}ci����7.mn]9w��J��5��o���q��`��Ld�N�V��Q͸��m�����t��|�mCg��k�g�孏K�{/����O�?��h�h��m�����3m;(7�0���q㹻W[�#�]P9��T�� �h��Ђ��u'Zl$j/M�j������d��8QP'*�E��~��i���l*�������1X+�%G�O���=���������W���R�V�������Uc���`k���y��j�����3��N�A��-��=�M��L\��䳩t����=4��%�L딩���ۀm]؝7�����?��5�����ޮ�+��?���Čj�������[[�	m.TO����a���x3[{5P�a	� ����=Qcb*��Dq"O�A,�ONB| ��I`Q�S��X��	2�����L�e�J��
>&1ʴ��	�����w�O�f�W�[���|n}��rsn�m�Zc�*'u7scy\oƘĠB�{���cP/9m��3��d(�/�Ϗ(M-]��i���ˣ�ON�5�;�Ή#K��T�uD�t@�P�-p4�G�1+��0�-�] )�����D�p �^ �5\"6�z����0a�u��2�G�ى���y$�T�SY��g�D�҉�$��LL�<�yx�G�K�k+�|�/�ٮ�-������(Hm���m*kqqY{`rF/
r�����=�S��;h����A��DVLAMj�-��ʠ���ۄ-LB��i��ď���?9m,����|U[l~y2VA�3~���
J>��ȗ$k(D%�)U&��M�	��ʑjt|bR�Ȕ�d�8/.ԚD���:��:{u���.=�5��YL�'��+�ꜣ+��ß��Kqd�R��e��n�줺1n㒥�G���?�/|����tin������u|}�x��y9�^m�G�І��iF�o�D�7���P1�� ��
���b�M�=��"�q'څ!W���$�1s��c��dU����S�#0r+F<�����*�� 	�r�儛>����v!��Ij�!�=	)��u�Y/{z���d�h��Ε7.��ϵ6ί�0kz�Fmaݩ����[����8�d���X�
:;:n;_������g�����n{��s�ߞ����ӣ��T��DSX�\���!��'���VAho򫹶�j��Q�F�& �-*6�~
��$pb2'i3�(!���o��(��-7�$
�E`���ͬ|U[r.=���r��Ʋ|�}�HR<�h#r�H����6{R���������O��{���k�,�!:E#B��ehsJb��QU3��e�:shI i�I�U1Q�A��i��C��������d%u&O�E��Lw4�`�V�hJ��1�r��B,`�J�կ~�]�/Ҕ9�D�;J�V檁�*˺N����a;ʲ��S�ĿRݺuˁ�0���(H�k��A��QV�_6����ͦ7�^[]Y|�ͣ�S�y��S\��i��з���'�K:A�:QJ
I7	Ixi�d �u�N`b���]<��`���W�}�%m��Z-�j�J������ 2�'�I��B)�8�GB	q��*EH Y�u�4Y�.ѻz%�.r�ƨ"�e�Br��̡���G�qX�2t�6�C�b���q{jC��8D�m�� -1,��v���M��Y�M%���I!}�m�҆�ҁ;���g;Yޜ:�da���Asj����>Cb���I�e��1�2��^�m���Č4�]�П���-Evc A%Q'� y饗��ԉ�Q4
��ļQ  �)2��I������,JN0��9�~��@�y��P�
@�T��z�A
�>�)� Dr (F���ɡ?y �s}m�v �E�dr�gW��Jcs�uz�?]:��C{�Db�!~�(����ʤ?(/8;&t���[r!K2Y�ۉ�S+�L@VY*�#&C�Uҝ�'n�H��Ԑ��c.߹lH�Z�������� 9�����O ~j�Qp��_x�3	cR�R@�&�t�CMo=bmB�T�]����|p�����>{p68jVN=a4���w�ݼ\U̬�	.���%��?n	��$t"��B1�@�"�ԁ�7��a�0�?��E�b:3f�:=�����QE��y�uas�|����oh{����/�Р��7�<�:t�ߡ8R1�'�T�i��-<H� ぜ�@4�OHĪg�ʓ�X {ss��� Q	36�|�9���M��#�d�&�s�ryuu���+�w����Fi�=��fg��e)&>�T%b�����]q�CFU�l�0�����4�����<ދ�X�[ą���z�ز:��7�Nj�A�A���fe�a=�t�óң�k�,?�~��ZgcnX�t4:8&�-��S;�VO�3��/�m�yb!z-l��@*�l�:5�65xS�$B��`�WC�B�.P>��'�� �#
k҃b!�O0Ћ�h6���i�@=��F<泰X��������_����Ύ'��jL�Hs�nб��!�b�m�)?9��R�ɶ-X3�YMG��<=�j�+a
h\�sMt�;5���=p�4��f��}<7;�>t�v��U��ͫ+�a�N{��~�{4�7��r��Ls��*�h�����
�^mW�����` s<Х/D	O
��K+.3�G$#o�@�&�:�
@���P���Z�4���c�另 ܯ���������KuVg���?y{�)q��͊����B#�X�Z�;���N����)ڂ$�86:S��	���8��՝%٧��SK��Me��[�_��3ݝ5�4m����e�ϥ��/�F��j�sTǻ����ċ��6m�\�?e�\k2E�r��bj���xag��
,7�A���d���_!�R`v�e�o��Ȅ����er?�\>�Q�"��!��q��|'A�_���x���Z�+����g�;��+����:k.;���b�<�����h�1�gf���*�	�q7x��L���I"�l@��G�Ѹ�u�uy����pu����ֹ�o}����~�q��Q����}��c(�Z���!N��C��B��cսX5zĭ�1��[��M.�!�
&�v~fV<`�T�8����J&�0|�8�e�&!�JV�8�=θ���8V��`����^�~cpZv����ǌ9 #��b?�5��/�{�4(Ƴ���4l�]�Q��&Td@fH����ݼt�?v�rܮbl'���p�{X���K?���������ս�_V*��.�?u��1Ә<B�$PMŊ���Y^�D�m�C�K-Q�'�ݠ� <-��P1T�#d��O��F�?x?Ŋ���?��	�?S	�g�D&�6縲j3��8G8��ШT[�.9��b��~����x��{������=�p�d߹����Dn�B�m=�}�٢�^�
a�Rp�)8PԈԤ���:O���h@
�r�2vey�^z~���[����E���bgv�������
�5j��Q��a	���0.⺋z:2�m/��r���pN۱hO��%?I���KT�;4&�}�
� ���������/Oyf�JO�L+JG�jt���$� g\�nΜ�8���;/����VP��p��!)!hF:n�s1��<�ǑaTb<@N)#s�=�޼?m&w:A�����=5B�'��}֮�]4�3��'����͗l\�������_��3t(R�?.Z�I[R�9�AbQYuI��޸���r��m�"ɒ��V3!g���a�-�K��~��h�1L>����j���gTv<�H+���U�l��.=��
���~�J�U+_�>���o�t�µS���n����^h:y?=���0����r�=P���0�f��ʲ"8Q�j޺:�P[@(~Ġ�#b6���4ue�v�͋/���_��5?ޟ�w���gΎ�~��+Q���1	K��!���.h؆��: �0�* N��H
,�dZY�'�y�9�*C|�̖g+�dS%�;��]:BA�_<H��	�S�*�V֔*ϼ)����^���^m�^����~�?@�ĺ�Ѹ��J�-qBg��Ґ�|��,]1�=¸�\Ƿ����� ��ˎ���է�/=w�z����{����_�ݳ�|N�knavv�w��#�_�T��R"gTf4'�g���rf��X �d �'z����$�e?�U�-?00­3).���K �\k�av�,T/�X���|��_}�ѯe%�Y:L�'��f���4{�|��s�Wol������;�a{4�c�.ׄ0�q๠�0wd�aY��DuӺFld,���E�T��ʠqִì,�j,o]il�v��o|l���G��K��f�.���;�B��l�|���?�.�-�~_oa{J��G+�Z>�D�U���ڵk�[w��i����Sp�x�^��[!��'�|��B������2m���V�P�޾�
<�۶j��&���1��;������ǻ�����?|����'�*U���,k���f����ϯ^������K���Y��H�{��x��w��V�e+ńE�hHV,H��T8�Wm*��i��$!K��֊�^Z���̷F��z����NϜ���L��a�x���df�}n�ܹ��f�
Tc_�f���IN�0L*E ��	{��D�b�����_Q��<�J�ߗ�GT§_�\� �׹b�C����y�	�%�"]�!�ae��ꔛ����ˍ6��o>�\ma�&}�UL��=���=�_��ҁ	���
1C�n�����f�X<�(;«������N���~3���=|l���~�4�G����be�sv���=�nw���B�U	2�l]R*R�jl�����O�œ�̈́B���P�[?�E�@`�M��$�����@�N�̞�'#�X��p~9L@!{���aIbnn�u��ׯ�;����j�^�z%9�����k�b�y���>�艑l*^x��<�zum�@��=�g�}�$~��O���|��Fj����ܲ�<��U�	iBQ� �Ey8I�H�/7?��$Bx�É	
J��,Ql��@�Y~�r5�Y ���N�"�/�G52[t�T�i����s�Ko�`�+3�����/m�]�q�ڍ��V}�R)N�հ�����,HR�[���E�'	���Q,ƫ�͆����u�唘@:�]��o������/~�,�>�Ͽ~�����YgXZ�ڣ*k�Ó~m��"-�6��glA���22���A8z��.01h�Nw������{b��K!����Y2���$&a#q!%�3�Ykx�F4Q<�$�'�R%2!�������(%�OB�)�SC=�,�4�����������թk�6���kk+���[��iNU��J�nEr��t��1�֖X[R�7æ�u:�4={�2=[�U+�k/~5>���O�k�t��_��`�\~p8�.��w�#Fk����bC�cl��Pp)a��>ި���M�i����NP��J���ĭ��I&�3��I`E��/8S�y5��l&���!و�뻄̴B䓵M��e�~iZ����/b/o"MZ�ƹ�k�����b����Pf~��atB�ʒ�L����U0�V����M�%�I�I�ϭ�-��A�A9(M��\���W_}�붞u��<�O���>�W.Ѵ� Ǔ�ͭ���Xi%�!Γ3�:<J4�T����)���hj"C�{��/_Vs�u�J�"x��]�tI�B�%�U@U%$`T�D���������v{K���5�Uu'wJ�ғI�qo�?H�"D=5D�|8-�Bx��'���u	���RYq�-JZ�_�}�k2�����L�E���ʢQ�e�� �9�?��?hl��$��zO&����9�S��2==
q�N� �!��h|bY�����]����P�ƈR{9 {M�%ҳ�E��0�I%��*<m:?W�8v��iuݘ�죩6����]X!�s�˘B&X�MTJj��l�GuTi�2�R9�������t�l�Ǣ�Q����k����h:N�5�h���'j|E�SyH�Q�v%�����IӨV*�B�(<�����{O���DI�P*�u����i��!�,~�W�����r����b���;ڜ�4���u�P�VV�1����UU�}��<0	��u��ͭVkn��i}�f������֭[o�ss��`a����k�qf���ޔ��
J��>�	ɨ�n7U⩺�p�l�F��`��7?~�3~�����$��Iq�+fZ�P]_4�7q��ಸ�FM�h�ب�w�Z�t���b���°K�!�X���0����_~�P��� @�?������xee��e_���?-���@���8�wf�دņ�$r�!Dp�9&U��>g� w�Q����5�$�J�BÚ+,�{��q�-nX��{��5��a[��V��O=KS��iw=HK�٨�iX����@d��D���IĢ�@9�B�T4G���c�d?3+ ��A���Q�^����6[0e����8s���]/�;����~���˗רŷ���;����g��*ih�?D��`˚1(ɺ͢-N�M���I����Ѫ0�
�~h���(�&HCc1hK)'f���n�`�!R�>t�7h������������ѓ�Fzgxd�\����H�^wjzc}�lx��o�$�ؙn�R�O=�3:l���� 8���M��KU,� 4
ԃ9N&:]*N�Q�k�/�A�ȧ�鎆]&Ǌ6�+˳o���O~��͛��X�<ھ�A2Ѯ��j�+*ځ�30�I6@X7��|��2�v��pyG�qs�OB�Кst�"y�&���訄]3k��>���k��Y�y�o������^u�f?B��"5Tm`#N�c�N�`�8��l��R� �y2D���'�yF<��3�Y�������M���Β�䜲L�nj�
��s:�Y�0���]��������?{��勶�g��Y�����T�5@,�ɶ��O�z����!n܏� ����]� TW����Ö�P�74��X�Վ{���	��8�$7���G]qPk�G�����z~~�{}�>|6]��Oi�z,/�l-7�ڗ���:S���ft9�O���I)a�[{O���*K@XJ��U&}5��؆�����`��	x����<�eo�n�s��/m������{��_�ܸ�\�9�r���������;z����k{Z8�v��fň���c��#B}��*�]��zO�x�uF
3B�����r���[���d�}���aS�x���h�i���}+Ri]��"��9�}L��pOii�F
a�! t%i�@���8x˟(9|f,<'b����<~b#��� O�B���,��L\�,֫oݽ���[?��څ+��i����K�h1CÞ����~;���Bq�X�d[p� ��$�І��A.6=,$�m9�|���T��c@�`���^wt����/\bv����w�폯^�ivO��SO;m:ō;��ʮ�'���7-Q��(!��$(��x��
�?t%�u3$=���^�bE�O!�I�"��|+F8��f����*�4sT�k0,��'7���W���?|����~g������a{ףU���m�u�\w�Y�cN��Y���q��z8��,�qD�D�hJûuD=�����P9����&6�"��:!5d�`u�v����S�_n�vڗY	�����`a!ӳnt���
L�g��9�t���'*�pP!�$ x�Z�\b�(�@
��/ ~0QR�t��Dn\&���`�Y����4�l��V�?��ͷߺu���_ƻ{۽�m�F�bШ�R�!K�Y�6��jD�M}���ک��9&RSЋ\��!~�tO�n��z��K+���V���7    IDAT�c�sS'�<�ZgGO��w h��co���h��,�(vXP !��~�0~�@�$Ѥ@��M|� ��r�d`<R��*���,Q�Q����X����Z��j+��������x�g���k/��Z��ۮ���L�g��mc� #�Pb���ӓ���*1�VP:��XG3(A����3�ݚ���qx4�503{:�4{����.\]x��B��>s�3S��2��R�bEp�������A��4�U (����$0%��.7��n3���G��~כ��K�ew��I��EXq.2�Qy�.R�Q~e���[�o}����)�Wݠ���!�%ŀ��<��c4�6\V�J����c3e�!�m��k��Y�Z�Px�.�+UD\%/~�k^��Z�3&F�����VWJ���u�N���A�Kl$uE
�
\%f4X�9�?��2IDžG��N���e8V����lnn�?�#+z}�t�.�r�UI/�����_��~�;��ϲc��h�v�����>���o����k�T|��bu�vݧ�?�A��I�i��Ϝ�H�D�a��l�����]�dX�G��7pdFY���u�d�-���~������������5z�n�S4�vN�������5���?<��S9:�?N�Մ'���!r��l8�O�C�T闊�a�� J�w�L�y2yE$�m�S�#9fV�AN�?�|���v���y��O?��?t�|1uvH���5�]hN_Y-����o������\��\�q�Tv{ f)�-�?�ŒjH3�8&���v��q��_lv�C����@�G{���؏�Eϗ�'չŋs�.][x�M����]����l�̳F�x��c����_i�R�����&��s�	��$
�В��5���D8O�$��@�o
���'�Q`v�,�'�t�lM����X��@k�m<��{Z�6����ժs���r��k��{����}��7�7���M��mN����B��@��ql����5�4�Q�&���,��	 }�Z}n�:;���\�2w����덽�W���C�͊���U���Q�6&�P��h��^�����D,�������I�0 Kl'2�]��O�?��#O_ Ǔ�˨�����8������\�l��Aш�{3�n�|�;?��ݻ/�p��s�#������������#&�m��=J۬p�,������Lb��~���C6h��[c)n���������˗.^�x�ʕ�^z�*�¢[��&s�z&~����kK�"������ �+*񓱉 <\F�[f��	�O��O�?�
U��z�YgL��Kw��H�k�Z�dqff�Y���1;����Ko\|�g�~�/�/\�*ϻc��m?}�M��|����{����N:����������{{L(�t�w�����.5B:)�U�{r�X(o\��___�]ذ��n�\�9��O�3L?���_S�b�Z,�b*�j��;�;��6�j$-_���pt9HA�P&��A�u��zJW� pi�L}Q�4Q�`�\u�̈́��L�~ XV��6�y晝+0+�����g����SW�foom�y�ʇ?��[o]�ֹ�j�U�U�!�=~����g��>y�����Ϟ<�~��c�ϼex��f��Qg��#i�ÝMy��T|���4�p����p���[���7�j'���b�1S��<��L蓆!rK�!YS^�9~�<Th��IH�Z��G�x���I4�.�7�gn��M��
���2+!�+��~�2+W=(Ϭ��3�
dTf+?'0�����2n����6je���Ii�Af
�ãc�����'�O��-��Z=��i�Wl䦈lW��<����#�K꾹��t��ǡ�ۍ�	�����vS��죏>b�UnD�y�q��E��v�^�z"9g���#��K5��}q6sn��D)�����OM��q]��5�TI>hU��Y��'
�IW��L|��ʀt���:�@	��O<�Gz�Y8�F�Y�F	�� �����O��t|Ի~�����W�eƧ�vv
a�E���K9 
BR=5Q7�h�/'��Or���u�?�k�/��쬤%���'0.s���U�������d~d�9*v#����"����*tee� �j��)ˋ�b����~����q)e!/�If�-M�Y{�5�-/ݠf���`�4#X+�gFlaS���1wi#��<�\m�P�3S�"�F��yI�ĵFq��X��q!k�X8�`�i��3�R��|���'��^R-����ۓ��I{v�3���z���,G��2�~�+�Ս�����"|6�a@�Q��F$�B�v��NIpK` Z �!5~x�7D!b�-"w݃����?~j`�7}a��*�Iߠr})C�)�0$熐����LBA`�UUe���K���<U��}E�E��n��"�ulMp��p������OveF���u���o�������W�O{��,�b��F��X;��1����9CɂY(R@�ft���H���P	:;z�퇕�Ϧ�n��haka1e�o�Ĝ*/�#���<�jT�����x��N�!���<a�$�2C����u}���yd�0�ٿP�������?��?ew�������g?{��w��[>��E��Im��^>e��a��Ӂ
1�fq�ʳUq�7�c�`7�0H���E��X�	�B:5%�#�Ȱ�wZg	�Bf�Ȗ�l"��b��P���d͆��>����I�y���R���ٚ�
���E|'}���DQڎz�ᙃ^!<�=H�N��H�$���E!�*K$0Q	�i����~�������ݎ'4Lo��c�ꥍ�����rqmy�;:z��a>��~��q\`�Ytw�bd���R[!a}-�\��8oSuȫ�E2=T����8�W��h������6�����~�gN�2h��|i����9��Ͼ����VeX�����!ES���Yo,��m�h�hҶx������Ǩ���$������	1gרN�����7��s���e�Q�e�i�uk�$X�N1ug�rr|B�}�yes�'?���?}C:������#�1�c߰-�\|$�8r�<d�<�R�ցn/8t�=#7-TT���f���{į�j���/�K�y�N��u�N��;w�a��$W�\��y������/��}<�j��2�aZ����ꙋ��[�`�J�!6�-AA��@���L$gB�hCz��/��!�K�.�XQ��Ŀ̋��4`_$Y�X�����s�ƌ}Acu�5s�~~�?}�G?����ٛݿ���ï��,0"�)���dqO�\���S6����**ݠ`�ٛ�e֘1c��*\d�E����X	�]f���L�ә6����zkc45ݯ���Ψ�Yuڒ�0�包��ij~j�hv�?m�LZ!��Z�m�̏�"�>�ݝ�;P��y����0��
>��="���(0(6�bq	?3D�:y����+��8�z��u���4����j�/��;��?Z;�4�x��çΆ]�"(D��3T�������<�8�����*��a,P��:�3��ev�i�6
HT)�<eN�������{�#�J�j����g/^��=Y���;�?���h�cRQ��<�40�j<��wQ6*�K!�A�0��$i_8�3��QQ�{'�3VH��{��	�y .'>x������#u��c�T
��Q���;��\�3}]Y_��_��?����dh!���[����`I���"HkG�m_!t
ň�Y3i�����f�=��p�(f��'�a����I�1A�N�-N+�0�Ye��T�<����n��Ro�YUc?�� ^�D�us�3d��1F�B
V�6�{�:��PϘ�+q���Xቷ���!��#�$�X�.�P�%ň�V�l0W���x���)�ʂ�xu�������ћo��~u�俳�t����^}��6G��E��d�o*r3b�6��l�'4�(��B`@�%!qm���T.�H�=Cx�'�=ZV��V��l�y�~�J��)aZ�ݩ7L��<E��d��p���L��FX��R]�8eVC̊�$��1Q���@/�@�u#M�p8 q�&>��G`5qLH&�g�(<Y���IdM�X�n)6=�2���֨�����+o���чϿ�ڝ����"��>��g��������&�P���B��	�!�5tL�޿v��:TU�!���XeQ;qbfR���L{.�?>���=Ev�V��^y�����9v�ڌi����ik�zec���;)2�Ĺ}��B a$F�����@W��N����.ћ|8��j�������XfQ��`���i�/̹Nɳ>��~�!�&�bg��Fs�^Y�V6�*.W���|���ߚ]�B�}tp��<�S{�Y��%2&G������-NG �g�$n�[!��z1��$a��c]bـ��9.�`�0��l�ͱ/;��0Ӻט)U���L唴�l����wtlظDL�|՛<��J�:�B�����N���E���g&���G	��$u~}!��?����,��XJ<}��o�F�%��|���*�����\y탗������e�c�Ãn{��)�q�EN�h{8VD0�ؖhm��bW����b�
��[��\��
�Mޖ`�}W��)��}�Ӎ�(}��W�[�r�֝�o��dQa�1;��(��/�^u�[�1	�g��¶Mq�'����x&��Idfx���g!�L��/*�K��EYrX��K^�~���O�Ɏ&9�����u�	Nr|���W�|�ۙ��?rf�����K7�{���y��m�qc��.kSV]�h�#�ؤXV%kט%�a� S��HGc�`�O�h��! C�|��Rl�\���[`��xi�-]���1�Xt��h�C��2�c�6�gG���'�¦�<mzr$�䩘Z� $<`��ms֕�[8�`bd/��T��3\0.�����ŋ��!�#?IiU<l[��:������ww�l(������W��O�<�z���c�������_l�൫���s7�:-�2�rx@����W�P}$��"�(���_�E�4E�0�^اA̎ze��
�fFiY�l�n�.^o.�.o�y���h���r��+�ޢ���h�h���ᨱh���18l?c�f�g��њ!3EF�u��}��ᓃF��['#<ǈ����Bd�I�c���i�t1��H\53�sزM3���r������q�r��^��?���ͻ��89� "@ݿ�^�a�$V�l�1I�yg�6t��b$��
��gGb"��d��Gt�/�aO��f�g�6����q�յ�����{O���3��2�y�b-�s�[s���Mچ����p	�GK�TZH���U+T���Dob8K�oQB�`�Y	Q���+=�KB�c�}݂ɄrW����Lm�i��v�G?|���oo^�L���:���C痮!�{6C2S'q�ލ6g�t\D�7Q�xҟ8������WTT�'��G[y�ܰ�	�	����r��5,��'R;u��@���T0�$�-��@_I��C~9Xr$�&6
<|�[�N�%�N0/*c}R���$����&!���K�8V����誃��(���b���R��ڜ�~��������<���.�>��:��GN1�y|�������ig��R'V5��>������L��K�z�Lay���9�����y�h���gO�;�#����Vn�����>s�f�4�%$��Y<������=��i)�` �z �}��#a�; D�a�Ŕo�����\��P����b� �Ȑ���o�"��?��+
6��£�8�q |!9��~�qA�IA���~�)��s��������<�{���̾0 3 Ap'��(Q۵,۱}羲����|�k;�NrmK2%QI��g_z����|O0�'E��z���թS�Ω��
��ӓӕ�������[}��^�୧^}cn�J��`rq��̀���ݶ�wn�z�ڷq�SD�V��٩��!-pH�ut��i�[G�V�3�G'��aϙ=��a���ꕅ�7V6Vm�߽�bo�c��DN-�u�yh�c.{���*�Y|�T��a՞�B4ʌ���yB@T�x�g '<��p$*m��S��|���E�?sn"p�i}�ۜ<]��-�B�+!~r��&��C�eFD�����5([��G�{�
��h�|���}֖n��ܡ[�B�P0�L�G4_�EO��1��M/L$��]f�_��7�|#�$�)yIۍ�d36������o��bw��!�d{58���X��٨�-��B��#O��HV�Sn�U BL�eK�Qj@i�p"������fw ��m3Sr&L�|�[�t���J���[����|%�]8[�������:�C�`pyeaqy~���z������>���� c���s���짒�@�L^e*�?��?;Ѹ�������U�d����.�y���� ���˩��4ސѬB`�ֹ!|�OdF� /��@�]%e��ڀښaY^�7��O��5�@��y�W�<�������OON`wP��k�Ö�a�~R�s�4����{*���j\*S�f5fwz����C�c��y�W���˙���QnL��9ѴR}n����ֽ���d��P7�#�)�q�q�1ye��m��d��C�F{� ˨�=��F�z�j��*�/P� O��FpAOZK 8h G&0dk�2S�)�L|H� �-'	�}�����C�SCj2��rW��VriE�\yP����C7�!�{�yMw�ޝN��9Q{�0na�ZT���׮<U�����{���qŭ���N-zq��2H5"�R
|>�E�I#_��-����"������G[�}���Ay�9Y�t�N���k�O�5:J��9��(��yR����8���x���+.'��p�/���	�H�)���sZ	�נ�����W_>zd%վO��siy����W(�O�G}ߎv��vT>q0:H��U^H~DP� �`�fC��s�'Zبz��q$G��9A�e�lV�J$�9H�!qP*�s��kq�9���n�}Gl�,,�{ӳ˓3��oO����WA��n�L	P5BR�I+ NcpUM���3��@�(V���"%E-��/���ʤ(��8�QS_K-���<G��Pn�P����`o���R�AP�^�t��O�����f'*G��<�;v����f��Z>�����394�a�>D�^&����.+��S#x�9m�&�	F��HH���E��W�J�vc2V��da\�ʦ�d��.���M9��=U���jg��T��ip8=(N����K����(�W���҅��\CiύD�{��=!	�S3�#���F��G��C��j��@���FJ��G(MlvtZxŊ�y����S�?��?|+�n�����C���F�Z>���fx��P{�x86>���������F�?n��˵Y�p����A,�m�=a�'���m�FgM-]ܔѐ��ԭ��l��9�l5'й�b�SM�?�g�u*"d����y2MB�?;��$'�_O��l�Q�D�-6r���M���՟ 󥑾���?���<�ﾴ^�].�<CGM�_�����ﭗ�����w�'�9�*����Q���/,�h2�I�b��w[��CCN�&��;a�υ0�Q�D3�Vkl�)��c��.,h������P��<?�ML/O,,:������5$�uN�Y���΃c���=p&���MI� \��	z�؝Y2s���N�{�����X�d\ ln<Z'#��������ʑ��qr��њ��-(0L�ό�tV�pe}��~�᧟}4�(������d��ΐuUD�@;MX2z�Q��U ��j!���c�Co�.<��4�xT ��c0nʌW��u�
�l,s��c";5뾏��A���}��ǳ��qN1�,
�E|2�.A���I��vN��� �S`~�b)���2�7N�魚��D����sN�#N��D��)���	��nv���/���w>xy��%��í[�0ޗ    IDATu�P�D�7$ú I8���C�j���N&C�1�����:K&��n)Ɵx��{bL��ȡ�%���*��;������x�b}�v��������u�+渂�؉n�m��R�+g�tÊ�+P�+�F�%��_?�2�yf�x ����!d?� ���D�'��h< 5�3�<�xI��%���Ŕ�=��V��qq�>��g������hN.u�U~t���ݱ�?t(Vӄ��4L�F,]"h;�K��Rt�LP�s��0�_�V�����"8���B�D�h��BW�Y�*����͹���7/X_�>;S܃$�z�v�b��v!��Wb�ilw�i�Z�(F�"[SLeԘ���<�g6��4��G3��\�/���m��Ӓx���B|1r�֬Ѡ���-����=U��6�����?���+�d;�Y]07g�Dr�q�N� ��� _�Ԟv�"l������ܩ�p�	q���R�"9�)��9S��5��S+�ћW�+�݃_--�G�v�m=ڹ|a����?���K_|��.,�7&0��J�ú�����!�2V��=e�	��s����8�T��Y�H�t=9!�x+�x2Α�^��������T�Z(-�Ӟ�\�ٴ��T�<_����O~�/ܲS�}||�v�iGv�T�MG�>�:f�ll PL�Y��5W�� ���o�#^�:�1����Ы����.{A⸐���ɓ�����\�����+��օ�f��K�l�`ݴj��=����j:�#�N�׃K�F� ��3>� �����*�s����\AOɽ�#䟞9��=��EPu�t�>6,�a�Rs]��T��hT����/��+�_�5;�fd�u]Uw�H�IL.�����w� [�����T�Z!Uc"�4� �)��R� �$b�2+��}*P�^X!V8�-�ξt4�.N���X�\�O�NϬ<��\ä�%n�e���PuT��O��'�����=���L��7ġu���t&��禓2G�h�9�FQ38=�����������?��Jq�P�Vy�/.�?���G�Gy�T�b!j��ώ@8 ���AS���0a	�.X^�M���#`@�?��'�WX]��5�`��Y�6�:��Ѐ=]�1ϯ����ՅK+W����U1wo��ʬɃ�����Zf��E�'̺?��]��` �����h{�:͜������.Z\H�47�]*�3�<��SxH���8冹|�i�7Ep���5GE'�m=:��_�������V�Ð`Ǟ�U�3���o��r�헮>�Jqb�oO���w�:Xѭ�&�hܲJ,%�]>tp�4�1n�9�	�	a[Lc~e��&^Ŋ�>�a��Hm������Ջ�/�������Y�Q9mw���;[_?R������a��XS|۰˵���2PB�&������M��{+DC�Bx�識sKe��9�8 ��1��OhC�zSsàgx��w�6vN�|�>7[����ǟ�p��Wg��9{�h�{�����گc�gf�h�2B�¸�*b0z7��P�X(�P�ŷ0���4��G�3ʤ��6���x�X�� �19�y��m�DGaM��_���bg�տ�?�2����Xe�}	J�i�	f�W�T���c��Y�Oos��-Y�Lri���̯`ۥ�M�$�Xv��S���e~��ť?x��7�X���� ��N�u�F^��nm�+n0�?��n������Jz������nbA�-VQ��\s��[�8�EL��[��&q��څ���k�����\�U�3����G�wUA�<[����Su��\"�=�?#v�\���r^e���}���y��$G�9���%�����FsҜ޸:���f���:f:������/LU�,Un�����{��w�E'���ݭ�����3k�Q����)^�Vgz9���I�"���0#`nA���٢��1;�I�ly����YsU�Q��8��̅ˋ��(�>Z8i��w�`����h��*fP����GN��w$SZ�ӘS��� 
O�r��g��%�%`�1� ˓^��C4Lr"���K�,!�D$�g����q�%:�7�aunz�Y��:���|��;?�����Sk��uK�ûw��~�����^�R���d����	��Ү�n�.�m�4�ꎖ��N��ݴ8�<�[�|�9;�K�a�m?mo0$�m7���U��\�11<��?����U'������^��0)�L�5׫����*�� �T����@�x2}f:as<^y�pO	�(	�pO�<N+$�|����\V�䜛���V�'�s�rVB�?'r�MV9�������@tBTd��6V��t4��T�����CK O���i�c�V(l����P�B��Qf
d6B�B�`�䧋fY__���766(�Qy�ݻ'�Rɍc���,�]�쩧��Tf��%s�/
G�>!7ëA֪5P<`�a�T$`*�%��C�.�HQ	�ᘖ�.2��믕_r�%W<$�"�bˍ�[��KA�d��Vəl�7ϙ��[~I�x�����ɅY��9��U�݃��q�B��x�^>��R�?V#;���7�S*?=��)\!9��~"��=sd��h��s�sZJ�+3TA57����j���-xB���4�P�Un�!�$�����-+,k���ҥKZ��,ժ*�p�lnn��[��r�hQrO�|2W����
i'~�z��>���K
�fmvbv���W�	~����(J�	S��3��
����=�!�@v	���w�f�17=�X4ޚ�7'G��k{���4Nkn=���&���ܼ�B����íG�x�"��vGe&(�	St�,�׮]Cg�Y�8��&:�4 >
Ö�(=��i�����r���l��^�Zz�T{�h-�7�q�m�iѮ_���!1�{+���"ir��
���GP�l�"���öN;�Q���6i���!��3�qύ�����_���gf�^ӫ���v)<nl�#�c�{8��Ƌ��B������-n���X��D�l=���o��.NGJ��i�R0�AHi��2���`z�>���q�'J��x%Du��1QH�e����-;D���sr9p>*؂KO��oP�:@R��b�|����w|��hxr�(�4f�4*�P�(��2�e� a("A��P
�|)tכ�Hl��C��`�+�M���=������ܩ����B]��0:��O��H���
ŕ�������Z��J�)LM��˨��Ӄ���R�����'(���y���L�Hj �|XjG�\�����B�
KU������}񻯿���Ja%(�m����[�^q0�h�����۸�}���=�$ri3,#�UV���Ǌ������͖ c�y�!� 8��d@M��?�CA]�^1rG��&N��֡X<�]SV�YYѨ��+S����v{ذb�X<.��-�s"��D�1u:3;3Y���?����4��8=,�����,&����̓�m����m�'v�"s~�?s	%�Sd�k~:t�l�z]��*[�(77o\�/��篭K������o=z7��c��m�0�����a3�p�����:$�+}�Fy���~�]4K'kj��EX=06zF��~�uz�8(�v����vTjYFN���|�Tک��O�A��>������� He@��
�
�f�P ��y����R~�+�ȃ�`˘ �fd�G���Qe��kp������_��˭G[�
�R4}�ƕ_���}���_�,d{x�p�Rk�I���뢐0���� ��]b^�bt�Ըh36dӗ5K�@mPR�(���hq@Jp$���	W#g�3�=�[e=��k�cI?0�����Ӆ���f*�������W��|��A�tҭ"���)`jL�(A��ic��	���M��{-��$9�N���BЃaA�?s�y����1�֔�C�L�(ƶ ��=�GGo���_���7^y�:�������4�c!�!�$x����/�S�� K�+%����
���^@���؃�#,�S��g0F���=s(��J"Dmb�7��^[�O��:��������/_����T�㾳ku�3
-U��7��95L�b�!h!����s �8�E���.�P�J%�3Ug�E�3�=e�����J+�G˥�-0Zz����(ǽ������|�O��� ��W3�C��M'�聂#�W�Z����)��p�H�,�a�ay����"�4mN�LV�� 46#Eؒ�&��<�2#e�ьkÝ$:���\�Zlm���ߵ�Ȩ=N��擪�\�?j]C�_Q �#b�F�`\�x?��R�(O�	��M��V�L�O��c���B8�������G�0�mg{����p���6^�0��^����/\ܰg�������0ZၟHH9�3�c�O�L�����yH�i	��N�ނ��_�f��1��N[ ��0V��1��au�͹:�^�\9����Gw��Mub�A�"aX`c�}(l �'�(m��G�8��(q�˄�@U퀖����a��=��ɠ�PK��N�Ȝ8zU��r��c��S��Di<;S}�������^�ٜ�k���!��(k]�0����a�c��FO�BYC�	5�݂@u 7zX� ����!��>��O2d�k��._Z��V���z�u8���܋7��o��v(�r���Y���Y�7��!+$ߓ!�(Z6Qk�<`	*J�-�����O~�E.O�"��µQ���t�	�S�P�൶��p�섀�V6{�&J�g�M����[������9���9��	QWM|:�v�$o�Al���ثд=>8 ���o�`���w�Z),��W}� �N�8����!uX��b��]�"خ휘)L�������A+$7�ƹ�(�Hk����LR��ȳH�7���?�={� �$!�#Q ��q��$�r��V��yYi��V��D��Y�	�f���҂��'Õ��_����~����D�}�:�V�H��"�ؒ2b�v���$H���]+ �uLG���%������@������R��L��1
��j=><<�� �k~ysqievv�:?��mk8=��"g%r�XC���e�2Y�r�H8Oz�s����T���s�q4��pD+D^�~�ڵk���T�	a�"�����X/}tp|�������������#s$�d�(?��ܟ��[o�49��V����^��������Hg��(rL"C� d��.4[iA>̆`��AV��WBLH�OO��.�Q+��Z�#�jmj~u��m�}p��ro�x�d]5�1�t�vdsi�?j�N+�������G0P lP�	�̐�!@�f��)6�E�SLO	� 1qiO��ȁ>�ƍ6k����埍�ijS�랝v��w�~�����o~w�_N���Css��\�~ey��g���ыW�y�1s��-�mo;P�Q���tD>x>��6�q\F-��Ca�,qG���ꃓD+7�<�x����c'��)t���A���NZ�Ӌ+t���������Q��?�s�oy�ho�Y�����$�{47a��\��<���Ć�ǶX!6P��Tv���9">q@�) �����G-2��Q������S4u�3O��4�^�,S��+�����7��W�6?x����yi���jm�}�9�v�ݙ�9LXnH*2-Ǯ�C��ak���W��&�HP�����Jb��ڪ���IDa9����8������ܳ/�rվ�i{���f� ̐i|:-yAP��UӖI���s���eĔ���[���Ѽg~%gI��*!IrCȐ_���<yr8|��$�����A�� �M�;�1�͵�W^���{o���s�J��3�J�����8e�FX1�٢(��cSNEM����L9���A�F[�B��h(2����͙�:!<Veb��I+����=PR���&��TW�Fxrh�K�9�����q<�q~�3ʛR	��8��'�W��̐����'��
p��t��7�+5�>�s��m����:-�م����-����>������a��:�}�how�oc��׭!�e!BĒw��b��	��
e�N4��B�|�[��be�ףt:h�n�8L��r�����ư�ټ����xc���b�]'��vl���'�E����>�i�-��hC[��(FU5j�����X��4 ���������'������rD��D�xs4��� ��D��aD�#��^���1�Ӯ�;�����L������}��|x����;lX��޾��ik�8`�8q��j靏OyA�*L[b�TL_p�5Lhr�Ҍ�x����� ���{-�)�Z�Nb�E��S��+/�XX��MU�߽;�X��ĺ��̒کkA˓n_#*R��r��=�r\s5���!�D.�H�h�Gx�����9B�0�=%�IrK��[���JH�)	'\D>/�p��'?���9P�S�A�1ʇرF���~�=֯OXۧ�������{ؘ�Z[�dRÚa��o�e�©I%�� `>�tss�mRH~`�Qr1�+�vY$!H�%4�È��U�B-X�����l,#���Ɂ�[9���G���'��PS3��dlR*�V:!w�ޕ��c������RD}�s��T
�+��׮]˒��]����hgL����y�"�D���[��tl�hb��~y�����������]"MGۇ�x�4C�!FQ�j��j��~�{|�?�H���J�����+q�{�z	������E�N�9y�����u`���A4���7����oA$$�����P8o#�! Ġ�˲Ӝ�����c��ꫯ�c�����^�u-��GNʅι�74W�>1ŉ
[�m&⮘�"��#۩�]>�<�'KP\�<�?�Xq�r�é�ܔO��|�+�2����*Ӛ�Z#G9N~
a�֏fJ��<���-�5�'���+�^���r������������|������WH뙉Ue�"$�/��b�6�>��x�y}�*�K+ħ}����*�hv ���.�	��"k��UnZZi5������(�
㭬d⋚���Ν�@��jvz�IK4�Ʉ��śW_|���>s�b\iwt�����q�d��k�"�!ޘ��f@Y��H���w����-�[���x��ߵc��޾��N�
G�鲛�PE( BUj�ˤ%���t6!�Ad����+��剒�9��Ҫ��<~BOd~��b������\~� �͍C[��T��5���O?���go:�ھ��~��l��.��:�g��K��a�<Dl�פ�+����g:�۶�[㝔*�a�7pye\k�ã��nԵ��̥E��ɒZ��3]q�'Y?��~R
�54D}�����puj�n��8���m��򜻗�����jU5E�`4�h�,X�dL�H��|�:oy2t"H�9�h�:�|݄_�lŗJ�9�$�uy޿�׿����v�H�xp�Ҹ~����+o?M�ܹ�]��#↯�ǆ����4��+/c.
Y��(fB��PJ�&����"F�@(�<�#[Ǩ���M)%��r��b��	-�lc��c���T�Z٣��0�t���������(~1NĹ�g��A}<��O�.�OM6�n}���?5
��z��u��(�>n��E�Ө�H�.
�\&�� ����xd�#xr�1mQ�P��e0*�R�Zeb����?���E��M뗭+v
MjbH��ݓ�x8�> �C�Y0|�졥���_':�FC��^#����4=b�K�W1Y�B��.4'q`��õ�L� ���ӕ�o�wN��9ӳ`y�!6��jM��6�s�!��(d�4��89\�ym3a�pe�䃯:��:
�K5'fԋ3L����~�o����o���l�6Qy���������<;�o?z8��E�+BPv����+��)hP���/����#N@4�=���cg�Z(Â�cN��kl<���r�R�YhZ��re����9sus���b�=uZoYF�R:s6Y���]�L,���<�    IDATK��)�8�ʺO��c�2�Ã����8]�E��6"���JS�z`�3èu��M `�L���1��Y9�D>���!��e�����������Ͻ��[ou�u0�I;�P� [g6|�(����j���`კ[m�H�e��O;.I�i����RX��(�\HN����O���6S���2c�j%�-�g��8S�g�z�ЫL:�������=ת���b�D�c�QuT1����49�A)ts�og�2t���O\\8$�\%~��x��| ,\N��KxvB"��
��5w��D�v���_�?{�է������C���Q��� /uO���کH�v@՞Z<8���4�c�)��u���ɕ��1�yب�C0��e�Yl�7x�F�Ч���(�{*3=w����չ�B��V�S:���ܐ�2p��T���8�;��T���8���p!Q��U���T������J.N��ĩ�\�U�%&�O\-�!�
��i���٥�+?�����F�6�; g����3rU�K�i�Jw���A[+Y�0�*VAG	�x��
`���:�>��PYѕ;%U|�U�1(�4:�cEV /���+�O��Z�/Y���H���ɥ9��-OUv�v�D�q��� �hg��qlيC>� ���@�Q3V��g�n0O�1���P9qX�/	�E��1)�y�� ������@�,(���n��c;�h@����_���7�9�m�3�`5I��Ô�3�#m\=!u�N��I�$��5FA
1L��$�Γ7Lh��6�+R$��12!�c����	AFq����jĐ���B�fyq�����q����x�{���5�Q� 	<�d�"�%�5�ꢐ�2n�L��'�^��+M�C����'�n��r�̜EˮV�N�4���UW1j�� <�����f��7�}���/�skzr��֝Tv��P����50��D8v	��J�	D���G޶����6�Nq�մ��C�)�BD_ ��b�*�`9��@�b��i�H��˭g��ۜ_���|vi�6���G*��8�K�C��D�3��Џ�q�L�$�A��SH��d?��
���#���O��-On���i�b�T I2g�7���j��R�%W�L��߼��ۯ��.8U���l�8y2�:���u|�i1ӿ��K�4K�����ٖ=�;���<�V�~7��t���dфMpKUG��MT��84/��U
�˦�xmer��L������.8���w�G��sD��������рX|$� b$�<3����p� ���Y�%�c�\rss�d�>�I�Ň|œ���t,������ů~�2�sZlS-&F}r�g?}mc}�-�n��/مjN�P�$FUFwu�`��p4B����\�(���P|#���o0��	�}2S����Gv���ѺT��<sq�9ӛ�?=�n��d�ܟlT�������n9�󘚵2nn�N�S��VТ�	�ex�gڈνRbL@�ppeT�pm�.D4.'$fS�П\��pF[��!�Tt:'��;;_��W_�˯��)��PDM�V��/<]z��^��ٕ&���m����k
��צ��c�!�����i#>�`�ئ��c9�o
	�F\1d�b�N@[�B���ކp��?.�1_,4�g�.]��X/�-�f���a�2d��ON{��3��nML5I;Frx�lNĮP|�e��	18��]���W��@R�9�j?�'����9�h<����
?s�zv�rn�2�������.��Ըp�r��7��z�ś�=7�V����������}�d�<�c�����y��!���B0�kI�O�j�'��33h���l���Q�%*3�������)=�Y�[����~�4�aU����]�Ses�y�į<�W~f�Ο�%�2�9!n���8~f�dRW ��X�
�r��$�F]�cmD�f�i�T����~��w_x����E������}�!��9�j][��X��7bSB`
�X��h`|HAA���Y�,�z�t���a�G�!tǩ�'Q��͐yl���I5���7776p�ťE��5	�������/Z?m��Ҥ	�j����C�uF8�&'���ό����%"'\�?�x��\ߕ��=ː��5��QH��74��F�8?1q���o]|��7מz�ԧ}x���kmo�ȁ8�����N�rY?���9+�8cYZ�\JF���_ybR���z[��������"�r�a{V,[dvkLM_�\�0��;Z{�6�G= �ġԅu�%,:W,sq��E0?�K0F�(WE�h�(d�O<�`R�U+7�*������+?%3��2��4%�[$d��t�,�_+g��KS˳��_����ϼZmNaG;��{�r�g�MjRg5��\���5��o�t�����*n̂�T@���p�S$��K�|�t����ۃ�����V�^��L-]���t�����i߉�Ds=�?(.��I�z��5�
�4"�0�95F�'J������@�D;��=B��osZ~�rz��ɐ淹���Gd��i��E���p"� 0���=�x+�����	�26�И����]�`�h�&�i��;>=vÃ�H�fKw�ߛ�h���+.�jY��)Ƶk�>��çҁ�D]����4� b|��AQ����:��E4jg�1�$|��J81�1��[8'so�޽K�Fy����O��F�JaDS�Z%!�����+dK=.�O�)�/��W�W�߾}[!��!M�R�AE���R�F$ �{����)P]Tjfj����9�������ꚳL�E����1��,�&���q�4�4e���S�sa��O��?y��!Jc�/\�^44��p��I�B8���u!����9�e��߲kj�\�L]�sbBRO��5�$ld���4em&1�����	����4t-Ğ�14�}&�\�����9�g.��<U$v8H(��ciL�b�؜]���'�1�y��QR��^���H���/2	�B
�zT���HF�8�h��� cR1Qs&m�)�׫{�����U�	�[�e>���������mn��8�T�#Y�䐎����ڀq1۷�ƣK��@
�x��!Sq�1�o��3��JK��	��ښ��u9��Je���SQ	�I*�;w��\��l9+�|�W��ho����\�1�@r>'\&س��B�8[G��{���\�\{����|��i�ȼ��h�m�Ɇe���B�b�S�Ђi+����w��P��4�E*�c`�;��k;��ݫLN[�J�J�}P����*�W}M \�:z
G����y2\�
�i���,������M�kA�$<�����O �z������e��?��O_{�E����°C�_��<J,�7��#���?V|è������=����9)w�[���G��v��������CX��i��z��p�x�9-�+������z�:�[j�(���O�w0E�@�,�t�H�m�k�K�J��A*�Pɩ�~ �2ٯ90q�G{�u2�7�����2��6�sn2�'<sm �嗿���@�h#�����⇟�����8�t���� {`��u�Ō�ZN�'*�[RH�56i��6Ӥ.o�5O��P��o� W
A>��S�4Z���<���Q�����>����L^I7!4�Γ��g[��#g����f�͋���;��3Y��g嶕�cob�0���s��Z���MP����*e�l��A��ЊA����A�1��F�Tkx�p?9e����q8]_Lm�调3gP�MLNM�����/���[�m؄����������]Y�RQ]��@.�u���3H| �ݜ�����0�J���ZD!+ө�ZQ���P��=dR-�@�* �pa�G�j��t��k�'�Z��:���013����G���^���$�	i�8��Ʈ���|��������S��	�?�I�(D2'�MP���Qy����'�g'�T#:��m������7�6I���`U��?��O.]Y�1��Vkg�T"F�P�E��}A��M��|�퀫Q<E����Yl�Q��V�M�Q�^Ub��!�6��:�yeF�ǀS�Qd���NjkN�u�#죡���aԬ�k��kT�����	�{߽���
:���X��85Q��yaZS�d&��H����N�8>:�K��=��t�'�Zs�����gO�"���Q�'?1������Д�AI�(
��믾�_~|�ʂ�w��<� -��g<uc��O����4�1��r*S�X&U�@��Z�9��-Xǰ�P&7���=j�7��
����Ő����cibM�]-o$)Piu����k����������6!���5(MЙ�|����P���,�|��j��/�=��$\��6�^��T�L�~�+*��E��*���񊃶�:Ht�''y+Pn���R���ک���W��W^�9�������߱�8C6��'&��r�<�%�=s����1I�Y�?Qt�['�p��M������jb��%.�ET�6wCU׋6ļh��z+[���XJ�z�<�o�����d&��J���íXo�=u	|��|,:Dqhpd�G��6A�>�`������r��?�s<���	��@΁�o���+@�7��Ǉf�8bVg��Nn�jkW?��_y��f��v���;Σ��G�
SE��掀PZ��p5n�#���]B�P	M+��%�@!��J^��D碬�
�J�s�p��D+Ɓ�
H8r�"��QT�B�BG�.��ĲN�w�-����job�ݵz�a�ap��Ԟޫ<Ř{�XO�#t$'mXM�4��R�N:��Q��'�]�W��
�����!�����O�/j-o&,��q�\��V����?����������3���r$�'��ʟ�0����X�!z Yڗ쌰~@/�O{|�Ш�����
I%��j�jAcd"M��a�м5�F�B�&6*ss��G+����廽��8l؀bP����u��&�K����ej� ��YKD7��o�`*]�U����!���3�^	��=�.&pr5m�B3�
�-�J�i�V"�ԪＵ񓟾������Tw�Y�Z�p�Pa���c�����"��Q0�%�E�������P"��\ y���i��UZ�hu�* I�䃭���՝oS��Ro�Z���;��uw��J�j|��X,�25>��e���3��	����2����є�?�ɟ�yHn,Oyf"�3J '@ؿ��h�1�cX�Я���D�bR���K���>x��sg��Ӯu ��\+��G4�lM�d�t�/�ڇL�!X:��Į��&�`-FuE��z��ɢ���j�h?f4�HM�Y�̂�C�D������(���לY�Y�kwf~bp��G�h���A�`r6�*K�E��"rQ3Jٟ�T�L�e�3��'�%��M��I��'������'g���َ���3ͧw�w�������W_o߿7�@�Aߤfss��7�y祕��Z�$8���5��Sg}٬3�.�^��K�c7N��X�`�$���,9�@��̴b1�{��/�-�c��fB#î9�d�� O� �褒0�Q�N�L��	{o�:o��n���֚��Yycgx6���gSap��q`l,���'X�Z�2 >}N�~f�T�?�%�<�����/T1��^y���YI�+	�<�d��L���-k���W��ÿ��?��=;=p5)�bƱ2?x�����{������ww��v4��>�5��
.�X��8V3�%t�P�8e=�4����N��boP��Ŝ�$���ȡ&b�	�G��BG�L���.���^�Q�1;�\8l�^^vwz���#$���{c�*��Sgn�si���t
k�mf�f���� ��Q\x�:S�@�L�lʕ��?x=��� �4�m$aFB�>ǔ����[�mD5�8�s�X�.�n^k����k��v����8�X�b�'W+u�ѹ�pa�,�Dib�	�H��u����9$ ~i�ƻ�$��������];!����k%m�J���Bmry����K��˵����$�&�PF��J��ɓq6k@${eQF~��?�'��{�� ��ejP�)�<!~J�#K��I��<�$� �[!�W-7m	í�~��s?�������5_��v�G'��j(�g:с��H��#��/�B7!�h�������z��9$AQT���cS��a-�5d6Sw�� M(�Ƴ��ڨaȐdb�/�������*���
��@��Q%������u���8wv�<q9Pd�\F�3�,D��V
?������r�b�y��Z�FX�)�����.�ť�G?z�_�/��{�������w@�ɯq?�A/qi��m�}
��F���	d�՞נa�����h�g�4���"QY��Ğ�w�d�����ڕ��R}v��f}���׮���WH���$V9}�*CJ`[�I��N,s&Z+&JG]+�L�+F��O�a>��?	T��6�4`U�~�6��`�h����q����́\,�萞,�:k6���ƕ����������o-,n��m�����3k�����m���q,3)���h��Qm*wH��ۆ3�j�7�S�B�3�R3(i���"�X_eU6�;b�k��d7��!�.L?����ѝ�>k��y�}Bgf"��PkM55GT �[��D	���y/�t��y�SA���A3i#D�@1y���N4��Wٝ�''A4~!��{���C����sa<�>*$u�880)U�������[G;�̚�ٹ�$�F-~8f�x������w|Z}�ɾx���_��W�,)����~M�r2[+	�1C��7��@�U"d�r��YCTDi�v��m�4�gI|���'$q��D����S?1�	�y����r�[�n)0}��x�l��M�0sK���)�8�2���S���*=�ƍ����Y�f���K��y���T�~y}������ŉ�9���o���]����R>�UZ��^���"J�v����^\���|���Px���ĜN|�p�sq�gT�����3��ɟk��u�n`�;�V ��l[�Y���T
���\� �As;J�
6;'CZc(%�&S'r�oN���)�4�x��k]EWVN��G���N��|���6��S�R�&�ul�i7x	bv��L�BIe�-%b
d���H�ԭ�MR���Q\���X!�p �u����r�Y[�z������2ݿ>�N�\�Z��C�|��m���/��;<��ȝ�PUVE����N��/8�A�Λϐ :�@.�7Iډ-G���8�b���E?�dxׄyK�͍�ͼ�2@2�����ׅ��#-33M�2`�JI�E��
�9���2�������ީ{7-r5Kt���SHlbf��[��͏���b{��}�y���-�b�5�(��Q�Cw��]c^��4V��ri�г�W�8ŋ���uo�޽��������e�2H�Q�LTʯ����)����ux\���r�x
<�N������"��Z:[X3I+\_�6?eC������}� n�K�N��?���ܦ{��B;�0G�J�fM?uI_�� ��q�%��m<8>m�N\��>l���`���޷�m}o�����w�߹��{�=|����{[G��;���w�:�ΰ���r���e��� �&F"�mφdc_�/AS)��������E����b�93;7=Y>>��f������`��׌�\���+`�SV�� zf0qy�gĄ@2G��2���l��f�#xz��BB$C˝�-���o��zp���G�v�9���������d����{Y�1`:��@k�)���Cj�>a2&�IT��=��0��C�θ2������Q��+������z�V�9�q�no:v4�ړc��R���3� @��#�c(
U�/l���}'��l����ң��UGe���$�m���V�������5��Y#Is����hra���Ϭs&��
ef�3�g��Dؙ���U&f'���R� x�!�[nb 8/��~y����kϭ��'��;���>u�[��?�X+�Cލ���H��m�T��k��    IDAT����k4��$7��a�[��a������`<���?P��t
!��壁`,dN��Q� �)�=��
��wb���Y�zxPenq;�4e�������Q���v�$I%���Lb�Ё(3R!�`��|�Spy
��;�W�y��h�r��K"O����noQf��_���?~��i�\zꙧ>����|�-��w���=��ӝ}2�c1�^�����'ߥ�8X�B���S�uPs|��N���)=ڨ3(tO����{Z8q�c�~R(aL��,��1G�|�W)���7�y��G��Y;h'NP7��p[۸pc���c�3}Aϲ����k���G�Ņj)N��Ա�Ʉ��̭!������g��I����z*j����!TSCd0=!|�S���a��	?}+#�`)6�T�O��ȈO��_~|�Ɗ-������~5m�� %R�jw�����/T�E�	g��B��]Y%B����KT��"P��O�~�7<ru��3����%��{jU��wa�:c�Ro&�e�c<s���b[��4�ܝ+TNv�I��B�6�NX��tZ0� �B�8:(򆏏��8��_	?�y~����?���H(�ۜ�_�9y���d&_!�X�tq��×��Z��l�[��SS�(U�ɴ�{���~RX��P?�Tah�M�� ��% ӄw�ޘ�9��?[K�5���5��EAy&�WR<���1qN2�������Ifӓ���T�F��݉��dj�ɐ��Y��Wԫ4�S��b"��&}%~�	��5}�a��XJ�Q�� :��#�8A�2	ۢ�	j?SL�FSb1��v��3sنy���;����ǯ�Ǖ���I�wr��9ւ�P�%bw �����2l��7x}Y�	���DiʹS01'@ǁ�1�2����_6�1�_�^YA-t�S��2�����	s���M���g�/ݘ�~�6U?z��ѩB�6²6jH�@ر�"(�.1���1T����8�2���-Ġ��'�ѰW�bOm�r^͉ �8?�k�<.��|��RՋ�?��|����jב�4�킷���(�}����rM�m�i�?����m�������Sɔ�����*[#&§�f�@z��!/����F� ���b�x�iG��I� �2W2�::!�2h>h�{{�n��l�;a�!'�K�y%�BǕ8r����fy#`�C��EN-�8F��ON4%ӓg'f@���"xk��Λ�� ,5��@|֨�Tdf��֫W?���+�O��-�]�3b�DV*���&ӡ��!>V2����2׋;��p�R���[��N��-v��~�E<+w��'+�y3ɧv2��aڪ+�9cyZ�̉nl�h��[��pae}fa�������G�F�̩��c�1��0���T����2���qA�Ii�x�D����r�$7��y����ɬ;r��ZKD�dؚh�n���˿����g�f��]^F�^ȼ��Α�$U�����ѡZ��%��,����qst�ɘU�Պ��=CƛB��0�I�ĩC��'�=:�M0����P�q�
a�i���=�����j�~yb�5l3����M\ F$l�hRp�C	(��`������OЩ)H9~�m�k~M�~��� ~����y��:2�����?����o���ho�²�����K����}�8�쒖��}�a�F=_��Vp]*�Z��EQ�˅�<q@��"K�S��,�;��@�q-�~_��ɽd��P�����D��X��ě�QF�v�;�}�L��%7�f.՚������p����⽃G�b�#jZjeq�hf�8Y�4=E�KGc6n���@���p���sT��^�e��hB�u��_ �蕫7o>��&�i�nW�:DY��E�*���������W����[��9�bȺ� ���b���]�o._z�n����q뀨 �`!�qF���+~4��c���'ə���	fc>�f�XQH1RI�aB>��McJ�R7���wE*��6-�4zv�}}	�̮,�?�������v��}{�)$�G�f�tca�mS�2�[p����"IG�ȸ0���	g_��@�?u�%�!<�Tv%!<*�����C*&�ş��fDT*���܇?z��ko�.������h׸(7��JLE�R�'�3� X.��wR��+�@��٨b5J��/�V!1WDmuV,2�
��Uj�F��Ⱥ�jSO���Ox�M4[����#��ىM��M�t5�%�B�2�)Ǜ�ԓ�*��t��WJ�-?'���sP͹��9�:
�3�>���L�D�rm�h2����`}e��?y��^�YX�v[݃#gr��D�4��0����h>�!t��kȬh<���/CJ��RУZ!�`8����xtH�2P'�\~dƳ
c7l���˨i���l�p׺����+W֟����Kl�l�k�=��[yvvw�펩Q�u����
�1�T��2~���e�2D9t9f��E;̞�6'��Yd����XB�����1kڌ�`|�2��wp���Ks|��ի�Ɠ�{;����!j�A��5��Ip���C�R2�ʰʇ�:A�B�h��48�EFZV�Z8�\�æ�uG�YP�`G�Fi}�V<�]��gS���L��ɥ��S���1���W���Z��5��h�>�<}WV0	t����B �����Jj�D��:��83�j�D=��.E�jf�Q#6j��Z�H*alԌ�A2O����>??�b��e��6������>y�������T��B�ހ�Q6�t��	���-Ʈ�^�lR�␺$PǬ�k�e��zK䍋�t�i�{�}��@.���]E}xt���]�� �g������<)�I,��R�dFs&��Q$yVo���31K���?c������sO�Ad����-1yr�9�MZ1��|���O?9o�������I��E�Y��ѼrJ�:bX���/Z!]E�C
w����Ă��"n=�����t�>�6�߿�.Hɖ ���O�ɲī��j��G.��(��"��Xp��Y�O�f+x���J�]O�qG-���ۯ����F�<acc�6[Vʣ0di��P!!)&Ғ��,��R��5,�Bȁ�GbT$9�
��ڵk�ʯ��*�'u���[5|�S��uP�Q���������2�zy������ٹe�3��D�9,w2��0��h/�D9}K��w�9Q�����/��D��`s���#�'Ӏ���{*���ϙ�R�ȍ���(	� (� �F�S�W2�JMyD�V��2���`gÆ�8y�|�ҥ�P{M�����!!��Pm��bI��2�J�D�!�r5��I.�9
�D��P/�6��x�D�3����b����deX��N2B���g0|'�Ɗ\5�-)�wC�A�!I���NQ����ރa�9(Ϥ�B&F�K��Ǔ�ɕ���s��B�؊%ũ�}�５����5].��3UCsB`�pm�QwTw��MO �h��.��R��#䎄��4
ی��h	}N���d�!�x����8�0�D����t���O���P�8:��r�\O���XD s5���΁p4"�X����Y�����?�zq�n�r���a�v�^����5j(����-Z$�5O��Cl��HL�y��Q�������h�HNT8VyE��p�(��2�28Bti�`�"9�U\ 'r|19?��V ��+��zs��ē��J4�sZOX������4 �z"�"���;����ɵk{;����v�l���
��:��X~I�pL�����muO]��B�ݽN����nH݇,���m:&E�c��ݫX�i���}119��9��mX 7�5*����!��H����y��%��Ť� l�*�l:0�X�T����twnw��T]�FC�8hlww�._�4�M+#�!P��"O��p��q�P�!��sz�$�sLH�k�`�z�������<|�Q������+�>w��l��5h9�5nYeW���i��>�H�Z�YofƏ*�(�0��v��S'�v{�9y���N�w[_�)�G�B�=8f]��̄3Y7��3�2�BÞE'�8fSh�bQ9�������%���E[;X�\��8S_m��ҕW��sS�߲��|m�l�}Z|4��;�۫ͅ�+e�����fL_��hznzeuaogk�Q�#Ӿ��[F2?U?7�~4�^�s|����1�;�����gp����ſ���z�b���{t�ک�b��cg�Z��d�4�s�<�iO=F<S?��l#�N�t��T�N/6A��t�>w�P�ı���k6m��|�<�W����Ά�T�%�/�{����*6;V�'�=X]��o��K�k����?������ot���8x����r���j�L��)Ob�Ɍ"#&P��A'�W~J����[�Ȉ���f��WR�̳�����������W_��S�����ُ߼���=><������9���v1���0g��Q�Fv`F�5b��!�)�Mf\(m�ʡ��FU�80r��GQŬU��0�Z�G�����,MZ���V�M�s�8#N|4�j���AY��F��R�V�uH�Ye�X��-�+3�fyr���g�N6f�4�G�Փ���bm�Yn��ae�d�[l^/֚��������Rsa�S<v	tl(�H��=�y�]T>U'��kOI�dԎ�N;�씲�����ʏ>{��ق]��N�I&�h�l�N3e�qLu�Xp=E�F��ф��G����S����@i&��1!�lZ�:b}jf�a��D�e=�Z�����q�������MS#2��B��\�����jת'K�U�����`��n�����و~h׾	Sٳ�J3N���M�BN�
 4f;S�� '�x
3�SH�'�d=91=�s���x0�s:����y�?�S� r���������Vv�㣭��t�PV���������q�j| f���Cb8b.��:���b�P�	�P���v�GC���ٰ�YZP푘6(��FN�k�B��֒k"�lt=��'��'��f����>����,?U���W���ٯK����6^�)��R�R#��!�6d��[M�Nu� >�:@|B�^e`3����<�s|����*��j�Ss����a70��TV�&������P�Z{l�/ך�F��9uԘ��1WZ�_�Y���Fbg�q��M��
���8�ٵ���EM����0�j.5@f��(� 9��o�Q�!�N���{=L�)_��O�I7��Zw��ܬ_���X���/��\����^'ݲ�EKD��y�T�Y�="���Ѭ"��̓S��9�����E�G���D��i������s��ѕ���c�0)�g+����7߽ٜ�<u?��>5������>:pXW�OH8�h��j_
NF"�Q%�۝A˙�M*V��5A�a���>ر-v�t�ԝ�W��	Q��@�Ny��: ��DC�4�� �0H�˪=y�-xOΖ~�)��g��}vW�q��yfh����-�X��4@����_ G[?!��A��Y ��S�L�9�W"����6��� �gP�Z�ۍ�n��TGo�z�ǟ�rD������q^l���W�;����|i��4�v �l]�
'.�A�B9��j\k��cj��|rz������9,چMM<U��Y-��5�*G�Y/�t��kt.�&�St����%��)gu'/�\?�|�r������Kw9l�\4F�%4q�Q՝�NjA ��KR!	T���}5���"�dT�SONjo���!p.��@���=h�l�ҧ_z�����K�=�?��u�g�<�b�BB���)j�øS \P�kKH{��A���戉�����-��PCu�T�� a��:Fe�@q4YN5��N�	�In��éUݏBgۣ�����gtk��0�/.���>���������Cv�B���]�@�>:�����3�~f秢���L�';� �S"���S���Ƴ�>ke!P�A8;�d"�/rZ��������΃��	�ig�Q^�:��'��z�EO��8�󴯫'�
�v G��`Q���d�Cprj-�����㺳��C��|%�K'F����b��TP�}mު�`:��8�R���嚱����λ$;�İge��^�+�n ��	4 $H7p���cKG�[_�_����JǶ4����4���C�4��K�Rk�{fe�w_ e?4^EƋ/�ƍ7�g�R��y�dv8^9:f{�׸�y��O^�����Z;wޙ� B��Fg�ݭb���VA(^�+�L@3�8 �?�r����JH�� ��H_��tU��	�]�z�Y�ޕ˛��\T�d�)2�K=�Z�N��>x�����--G���|`}��_���5֯�R�O�Y<���b�cU���a�!�9?��X(m`����G��Ǳf��X��E�.^EA���`5_s�������A�+��,1N�` �;�n�u�2X{��֥�7�����Z\�ng��}�%^;��O��Y���%���,�5铽�g�}��6My��҄�	W�w��MH+3Ṓ���--T	JO�SU�X�*1�g`8����{���+Wn�U�^j���A�}F�l�l�_�)����~�^'�D��
�"�$
;�EQ�|�k6fq��Wn�������<�ݐ��+�h��ᚘ&�[�ekr�+�m4on�s����o���lC�FC�yth�DD���h��a�DYfĠU҉�V2������]^q)��H��)�
{�L�	�}���钟�������r���~����ƫ[ǧ��@Ģ!� ��w�PPLU��`C��#c&��8������60�dkgC��Z��n>�X��a�?�γ�fo[!g��\��
�kS�,.'6�Pĭ����'�y���}|	M�s7bJEs�t_��2��"u�]��.r�8���*�*|q�ʣ�&0�I�
����Q�X�kxj[��'M�7V�BA�|c�������7��<����=3g��SѢ8;[x���.7���ub�|����dER�w�a'�g�P�΂�@@��7�d�������ڧ����8������W��õ|��,�?�r_��P��Q`�Y����7�i�hHl���Ћ�fw������LAp�P�qGF�n6쁐��Op@���4��/r�px���2F9��)5��J<�	^,���1��r	��+�k�������l^~C�N�I�3pVA^h� ~9'ဃ��S	���#�[�P�٬-rE����ɺc5�G�8$�9���y�#=/ڨ2)�X6�cۣ���bn�St���.n�8eug��_���x�����ӂ�z�����:�J �]1�b�ȀF��&)\��S��G�ލ���c�	��S��T�t�$���E��OS1?=Mi�4F*I�$,_זJ*�Ju^<RR嫙x)��sl42�R�?�,�Kk�Bκ���E�6�"���@������Z�i+�I�ym�ؽ{��ܼy�O����	���>���م�~�����#w/zJ'b��C��QA�2�z�!eb�u��[�M�A9��:Qy��<��~z�QP���mJM}�v���C���'���;�U����MR�����7���C��8>O`
��P({{��Ig��v�aK6y	r ��дt��]��W�7bo�h�4;ڦa*O%�&����.ȑ���L�u\f*���#i���V&�r��[�~����\�Q�bI{�F��%�)���Q!��;��D��&ڠ�L�c�|+\�l���d�7
���@#�Lϩ%|U��_�$<u��O��1�*�c2-H �.�`6���̊u/��,�bdL'��l�n�ş���+ܸcV�v( ���.�'hl�j�K��vW�l֟��$���\�����)����o�Ϲ�����v��]'�v��k�F������۰ufCV]�U�a@��N��d����Z���  �PR&�䎩��m>��j�������*�����%S3|�X�4�i~�~h��ųz%U���s��{1Mc�ʄZH��;w��!{��Q�{�g3O    IDAT&�bc�v�O�����*�疣B�}�j�Gr� I�>����L?v�1�jռlvDY���x�`Qj0!����'����bFB�)ϱ�!����P�ֈ���zT�5;������Ү���#ǋ2H��!s�)���Ivy�%�1x���; U��X�~���8!f>-FTRB�bhD4�$��6\��M-�K�fӪi�=9��ۓ[t��q��[D����<�œ��=v�����d�>9>\y^\���ؾ�����Y�ݭU��F��a�#W���� �N���c��������޵+g��W^��ig����X/������K`4(`h.hxJ�l4)��P	�����[1�θ]_7�ˋ �Jc�(�� �~F����?}�Nb���������;����ٰO�_Z��&�<+d~H��Q����,�p���}�B2ˠX�Ug�v��t8���x�O���\<�W삆i&N�R]�������ݵ⚸ގ&O<���:ΰu�1Ν�Oc��l�A��u���'�#�Ze����>����O����R�-������Ϯ��vy�Z�!�$g�0��RGZj�s��Xw.v���^��{��4x&�B��H����N��E��;���ЫE�9��rsc�/�՟�y�Re:��r�e�ɂ3X9`�&A�E�ʜ��+��f�u-GV)����u�e�?���{ܓŠ�X9�V�pY�J���Z�Qo҆��A�5������3&D�8�*�ų-�)^1��i�:b\�����/(**��+�Ǔ�N��'/��[|޿:.=�2�q���Zk� P�JوfF˲NI{�
 e���
�|0T�F�<Q�ې<զ�:SUF�e�|����?����N�mW�a����z������ɳ��g4GG��&i�U�
�0�S��sa1	��K/e�Y�\YA,ǥΤ�w�Q���#�qr����r���Đ��0���z�$5+m|��E�(f�9�R5� w��d#�~��T?���qnD=�w`����~ug�׸V�W�������{�����/r�G�����z�����rX�7)�!=�c��/]��;�~�H-�2*LZ_q���Y|�tJi	tF��(%�S��1Y���T�by2]�����;}���h8�qwt�B�
���&T9�g ��M��.C�}�c������g���Oڽy�=r�6޳���LMc��Y&�t!�x��c�^k�	ʷçw��b`e�FU�L<���&#���.�|bee�����z��7�W�C���4�B+"	�c`�}<�"�1q�� �_V`8��&�N���P�\2�=�SwR�T@�@����f@�jGP"ۋ񿾹����Ν�%��Nh~���`��*����1�bǫf�.;2ԅ[���IbEt��*�Nodm24\��-��c�4�5!٨;+|�X��(#��F�__VƓF�P#�_����!b4ĸ�m�n�D��� z�k\[�q��ޝ�k�������K!��49��8	/Ĭ��"��@աVp��J�~��X.0l})��W{���=� ���*Iܝ|9��j���ڶ����K����O~��/�M���q���Џ*��oq~� �e�V	ͻi�8�Id�-V)�9J$mơӻ�9���͙�z0�|��0;���@{�|h�P�
M�R��ř(&�֙�d�hD��Ng^��1W͌2	��v�{��7�ͽw~������pZ����&;�Jic������S~p�

��@��%��(�1!�}�Bлi�Sb(��/�[�AFr�T3m.��{�^��w���i���FhI�P%b,j�L�����\qf[P-�G����\�d����|<"J*&��0�pً��Z�V�J�6'!b%/v�S�F�<�:�&��3q_�d�E�y��R��i���|:��jlo�rݕ��6_~��˟-�ٳ��#�xLa�ͤ�A�|�"�GWHB�ڲ&XG�L0�1M���'Ё�^�2��.?ᛱ��2�%�H�4L�^�,�Vi�t�k13���O����v#��="U^-a���);|�m��QД �a��ǰO�4#�a��E��	���l"���� ���m�;\�D��d�����ޜ4+��j�����������Hrk�ש*��Jљ����}n��b��?yt�����.��}Y��8��z�ȯ6�f�	��M�"%$ݕ�L	�	��-?��5(��@���ǋ��t��Ի���N��+[?���o�p3?a�x����W2�$�S�{E�L���0���# b:&��t�c�P�?��������4#S�#h[���@M`��Z��V�o��׊���s�QZ�xTdHu� ���gJ���!�:r8/�8��6?��w��^jl����v��o���ZĤC}B��2�B r��}+?X�]	�	J@���E�[邟6�7nܰ鶩4v�:0O��^T����[ݽ{�q��k��؛�Z�����?z��۷j�9:���܇"�?��a��D_{�̼��S�#�x��T�c1�"� �KM�î@�؇Pf���6��
�:��x^)�k�?w&p!?-��q=�r8?<&�af^�In��7
�����d6�O6/]\��{߹v���G_<nNNG�ļ_=���x���V��Mo�ا�-�`�.|2X������-�]���<RƋ�����h_���&w*+p�p>�AH�\�O�|z�?}~����8��r��^������������F�Pv���ba�C��+��
BspDqp�m1k��8��'���d�� A�caq�Z�P���Y^S6�m����ӝ�d(��:Zl2*Ĕ�N��J���OW��}v�/-��˵����po�����{�q~�����������z�r��Z)�`yѼ�'�^�6��P��:�*~����� ��#��C)'z�]r�(a� �tz$-�*�H~��V����;�����o]�������@�e��8cGM��NH���{!�f}v��02�I�H�b_i?�sτȮ��S��v��q�UO��[U�Q�����!���W�86����G�S�U�~�Ő[�v^齵+��җ��Y�[vv�fs?V�����e�	Z"SN�b~�R��	�^� c��UI��TB�OH��j�����3_)�Vv��۷v��;o��R,���d"���z�6o�.J��"M���A�^t�j���^l\ͬ�LGc��k,������y$�q<�C�Cf��Ub�����0kXY�����y�������)�Wj�����O�!����!o�Yg�3-g��z� (y�'|�#��
����ӣ����G�.��D�T��+U�o��h~�G��g��s�"�R��̯�.mT���+o��ە���ӣѠ�7U�m�W�x�:A��[(x�r�]=��1P�m=��i1C��k��%��J3tID�%�`�y�8e�Pa�E+f�Y��z'���1mq��R�U���/]��{��o�˻���p�g)�G�|}#�� T`�<�/��1����F�F^�)����?3�}E% -���|iw���L�2(}�x��9|�F��b��"X,�yk����ww�\-�v{�Q��t�>��r��4��¨a�?�*}.� ��d�����JjB �;_������l���W��^�p�2����k���!��&�g��5����om����޻|5�������i�o�X�O�p�"�&�a!�T�L��j�L �	22���~ꅴ+z�GRلϞ^P> ��T��(�ً)��br.���N��V���x+U�ǫ�:e*�j��T�H@�C��0����%��qA�6ϛ��g�y��`�zis���Pey���
i�E9�-��`9���?����Q�h����������i�� ��L�fr������<y"Syu��'�$�h����ｮ���w������zMAc��u�����~TP13�ZZ7j#��p�T�IDN���T�E����~zK;=LMuW9��� ��uO�|����G�����;� �����a��$M\���eCb����k	�/�ޒ�E-��)��GB����
����ݔ���]��2ڬ�jS ����YG����.
/g�&��2�J�ZU`�L��O�js��[o�ES	t��m(4sjO�	�ӈ�U	����A��,X� �2i˴��Z���$ ���3@���4�ƹ	�7]0b�GPnk?�{��Z�<--�� 6�Gw�)aD�J׌*ۻF��z^�j�E-F�7��g���<Yv��b-�X_��U>_�5nZ��_8:?��ʸ��lg��d�93oųbi0����'*����P!}�"ܡ;�/p�e������ި��;P ��^��B� F7Fm�Ֆ�L����CSS6����W�+���}�O�[�`ìܪ�T�'T"�j�"�0@�@#��k8dlcNG�9�-�����ѳ֌��WM����|���r�Vq�=}���$����5�>[�`�*���L39�c�B�l�%�%Q�?G|��b���X-n�V7OXh����f�L����X6g�)�׌��u�%G1؟�"���ԣT��VS��(n�
k��W]��؋@m,�ݻ�F�P��2��Y<��NŔ��'l	[[z��j�t�"{��8�#�&B����>>�DD�3l&?�l�wF���&�Q���������X�=���a4`�	j�V�����f���I����̭4�dln��v�CcAD�L�/#n���¤�m�1�@|[�˛�*v>y| �]����(��J�8�!�	���7�
Z8�-a5�&xjd��N��pU%.���B��=�ܽ�i�u"^�l�cЙ�m^ݾ�����y�t���:b�C���GȽ���v�E�MR� A-<	��v����q���IdϏ1ī��U��;u����D�L�,��y��y:����r�ZY[��m��ݮ琪*���I�X�`V�
/O|�}�|��{I����Ѳ��vV���Vs列����Q���+~ypc��N��R��/;`B=�"t�
���+�8;��*(蜙�i\$�]9���� �~����vy6��C��r�	g#V����G~�zqu��w�ݶ��8����!��"9x#{�0W9e>�������Q@������h�,�R4��2��lH��9a?*F����~���<vw��q�M�\+���z)Wc�����%��Ԉ-��2\g��`>�/#:k����С���;/|p^�����_-zAms	q $@ۿCG���D�h	�v���۬��PBf")�^f�3���b�����,p!��DU�&�-�^��O�G����}���G��T������7������Ѵ{2=އ0h�W�*�!B�f�K�%��O�Y{�1��Ƥ7;��=:;m��;۟�����R�N����.(lt��x�I�ƕm}m�����z�Y\o'���rv�@$L"Ǵ�hHQlV���c<�(��'N[͎ͭ�����������k�������jy������{ww&�K�-q�R4Ȭ���ʊfs���b��wTͭV����[�L�ct0�C a��%dN��(2]�)S1�?��x4����l66����n�~��?'���z�DY���p�$L��oM�P�#�AK`�C���p�j�N0ٓ'�[\��I�$��|P�Ҋ�-/�c�xr�
��<�+�R�?E�w������FaX��++k��5���]���J�.�ȴ�vh��ͭ�ʍ��>�^�|r�o�\�ˍj{�&�+�)`'t��4&��!���� �
Hf���7�A�#��
����2�W�0�%2�'�7��%��h���ȋx��j����w��f}�|pz0�5E\L�_�Ò�C�Z��x9�S�27Y�;`�d1�O����a�3v�հO=!@�f�9%+1/Y9t��O�nW�-�U��m66�ON7�6h�p�Z+��˥&iZ�'xN�"E� �,�؜�n���d�>��X켺�s���>m|Y�w�w˕�'gr�����)��ie^j�q��Q�M�p%L2HF>iMXpNi	04ӡ+�rbQ���@������#N^�bN�Cf�R�B�Zz��k/��(Κ�N��e7��[�;<rbc7�4TI�f��Y牥�38��g�Pwf�m��9����$�LR�Ɓiz,�պ�X�QX�6��Z��*��yue�,��7�>���7�c~�z�9��& �}�Aw?Wn��.m��͝w�?���֧�/��=M{�OT����-U)� i�ʯr��/"!^�i�"� )��2�i0<A^�2�e�<��aF��]�#q�"�1�,��ب�������#��''ǡ.��`����H�xv�E�.��+�M�<p��{�>�L�w��a�}:m�G�G������1��FfR��?$����z���Xk��j�^lV#^h�6��Vxyh=y�rĊ�*�v���pkeY�a�8�ә-����/�9o]������'#�v�Q�%��Vv��d�	)�Y����.�5V��sN��b���9��BHC�.��^&�
{�P4�v����&3�&7�k�X�goܺ�Ï_���f�F^��=<^�ņ)�G�8-$�8̋���p�M��q�p�?yz(2��|��s�He����"�����3���Z��Ia���jpc���U�Z�o!'5��E�$V�Ô�y�\�R2��>',',�xm�q^ح_�S.~q��Q���Γ�HԂ���2��1���!�{d&�@� ��d�k����=��@��le�����?���Q�~P�1|YlD R����L��oZYm��l ^���G/�#���S���P{�~<Q���~VE����`�Hz�1xv7��i���N;c�'���=V��n�/(({:�갴
V ���J�_�p�+|�5��d���c<A���bVŭ�VY��O��/ lϻ���qywu}���y���>O�/�m��=B��xǢ�x%�?.}���]	QY��!�VCC��]�4�\7o�Lv�8@����K�%� �on'~��>{���^�nc�Z\�l��|x��n��T8ڢ@�y�b�eęx/��|���B6�؀Hۈ����vt�<�N�=l����\�c�#�x�{$_\'��2GY6�������TcUE�8����q���l@�AL��yt՜�Ч��o�_ؾ��{�x���Yo�ʧ��?}���U��o���2ň�"|��9�v�;��lP��9>}�l�>�����u��(u����@���K�n�x������+�X��L�	���y;���_~����?����H� �b��z����.���w����yi�V�0�8��<P���v0蘒��x�l�	�3�9��ɔe֚��(ld��iVǌ���̅謱���M].T�s<vuu^/9�m�Vp�/�GnVb�<XXVڂc!Xn�i=ջJ�2�Ra�ƥ��+w��v�Nۮ��fLZ/���nn7
ճs%�L��AA��K�d{�aӋ����v���f��,'�T/�$��)'I�[�����~�sk�����gj�|����Ε7���X+sJF0��2b�,~[�����a����>��B3	�6����ۖ��l>2�Sf��J@)ma���CU&�)R�� ���JET	s�r[Z�7�h�6����K��W"�k�j�;����V��>9
�[�����!�
�H �V�l�7F�]Z�  f�I�������F!U��-���!��L8�CaJwn+ҷXKCj��Ja�V����?~�֫��^�N���0������XR4�b�C�c����*�@f���`���|�xm0�@�XCmd2��/GT���̑L��1��sg����V,��"dV����m,�࿵⥫��O�g��ѱ3;���32���?��A��A8��og�[�N���tO0L�$V��Q��q������Js�(�˳�c2&�2w��4��� ��ͯ_�x���+��(��w��:'�`aG��[�`�#&L8�ŧU�� �L�
¢[�M�V�� )�A1o�N)� K�@�o�˰��,�l��?A$�    IDAT`�	��P�|��Ql�Y��<{2(�n]ݩpx\�y��U����C��w��F���U�aXb��UHL��&�+�e�Ϡ�ŲkU�_f$�Z#?�	�z� ��c��IϜÌ9�:�}FoA�G����
�m�w�/�x��g�~���ߜ�W������A	aHXU�V�A��z�g�0(KAM�<�E�;F���Ar�tT��V�`%q屿"���=taՉ5j�̌�1ĳa��䍶�'"�r+�����<Z���ow6�
��w~����7�������F�Vc�˕'̐�8�YL x����00��qZJx$���2t�-����ҩL����ʧJ��t����Sf�<Րj����PFZ��ti���^�����yL��<2�G�q���m��apHS^[�W��+�V弱����"�����9�V��pH�gEϹ��*���r�E	�"��_Gh�|ѥ�&�ֆR����G��VX;	�q�7nܠX��L�J����|�`�z���(9R�|c*M���Ppd�(�+��r�W�}�'�P1��
�Gگ|ZOլ��z����0�8��@�v��[��&�)������wjբ������@rzN�Go���� "a�e�a�b۲�A����"_�K��݄�$HO���nM��ws?SNʔ��&��.u�_���F
���/ �1�*?=�
�\�ǋ>�]Г ��93�7o�T�⋔a.�AYu��e \U'/{'j�ԥ�iE�5zQ�.Z/SZ��yхN:�$Y��˓�U��$BI١"��~g4\/N�+C"�S�|��	�X�M�L�l���m&V ��p{�n��P��x�-��O�z���:F�Ш��ս��O�>=����y���p\q�M�Ɖ�8S���Z��`�Q����������PU&���Qa������F�ݕ�\��ICn&�� �	8ʻ�+�N%u�O��m��^1�2�����nD|Kc�f�f55��0�㝹C���vp����N�%���w����?����{F�98=}4��b��Z$<!;��d>1�@�$�h$����[h%9v��'=�̚q,-���������!�D%+4�!xJT��PH$��SZ?=������d��|	����{�	�Q�[����7@ib�jӻ��2S�s@�^��o9:�����^���@�Ê��]��^1�OM�摾��{탮sm���N^�|����ڃRLPW��-����h3>�TB~�]��8Z'JƲ��	����H
9��{���������C"����+���	Ts)���B�D�QZ%�;<�|�vi��K�S??z��\��q94@�����N�Ѽr%<�H/�E�@>��=JJ_%ӈ���6^q��
$��R ��W���w?i?z�����Ѭ�>��.���?z��y��~��1�gÅ_�='�)y��v�:�؊:P�i*�N�tx�|p�S"z�;�v�$m3"�S;����CQ�<I�[='N>���B��>m��n�l7w�K��qi�����Y��9(x�!���Ya�ò�Bӏx��ڠ�sl���.��ǲ�í�nc��wpo�w��u���b
�zy��vٮ/���C���b��^�����o�)���)6�Gf���Ϧ�L�Jd�[(Ӏj���0lG���/��������!�ӻ�Qv7�nۤ��U\�x7�ma"0V�^
��lz��N�O�����i��`��d���ڐ�h�|?t�<����3$����e[�^w��d����ƚ��
U+Y�fu�gFDu��)H�!���|�lP)�<��J�f~��Y�y�;ӕ�����>\�T��A�X��~�l���P�f�G㲥�Fw3��.�mψ�����FI��G�/0�b�.(�#can���k���V��̫pW��?���2>}�kڳ��I�S�Ɛm�Ƞ�EPۇ�=��K۫Щ-���������iK���x�I������Ģ@�U��a�l���
l�l�:��k��{�w���&6j�IiV/El_`d�|�c��%5����F��InQ?�z���K���'����Ѱ�`RX�Vzﯦ��W6��l��昰��E���֥k\o�Z.>����(��Bc��i��֥_�%����A^��H��U	���.�&������_����yg�9���8�A?�e(�B�j������b�jw=;r�찻h��8��W�� 6vJٮ'P�#J����qi3R&(V������ɐ]�vk}��Fc��tx�ʼ昭�^��$��>f��!ԍ]�X|�'M��t�8��/�.]Y�����~�.�5u�� ��A�Ф�=kl�2!�E��6�ܒ%�+ܖ	�H�7���4�F�zZ���V��(��y�
��V���(�
���Ê�^�����V�p!���uV?r���J?ԓ�`�C����.sp|��|з�O�Q��r�{�PY�Bh���g2s|��]E��A�v��iko{cg}ks���[��g�-�k��t�<������> M�JDS˭���{TK�����3{v���M�XX����mV
uB��5�Б������yt46�`b�����L?�\�tyՄ�	��~z�����ؤ*��t���@y�3�aO3=�[���/>db�F(, n-���/�P�R��g��
!y���1���[����9c5��H��^�gJ�cJ�Z9�:$�CGZͮ۷�+�hۆ����Bqo��_ܨ�8)�9�a�)�̞��"^I(gD{B�=�VV��d�͗>�|����?�C�?�_%X��+�Z���lZ�)3D+��q3� �@n�1���KZ�r$�S" �񓉞x��EI�qq�TX����XKƅ���>��������Wgk���&d<!�v�g�fPD F��{M�m�N>?>霜:��N��%a֣���䊆0?3N�5�۠�J鴵Zbc� ����F�1�趶VXc"� ��ω��|i��"��]�b�kDL(^ǈU��j�,W�6�7on��k�����V���0+��z�䠷Xo,��/& [��S`f@;�3icfD��G gD����J��
�)3�=\%��'��b�W�8R{�ŗw~��7_����@(���0i �$�1����!��Sj
�q���&�;�����kX�ΰ#�6�D�5ZQ�4.f��,��Ʃ��wj���\��[��/��V7�M����71����*­kR�: i����k������l�ʕ���]�]{�ˢ�
.�R^2.�y��`h���:�It/��+5�V�%���W����J�p�2(���tr���@T��[�
Ӊݽ��v��W_�Nh?C[$t�-Lxj#��"�J��ě��`�����~�8������n{}_���3��bX��C��J#ͳ�y^4��0��
E�{VVeg.��$��@Y'@�s2�E��՝mm mka�_̫ە��n��Wk�^~�;�s2+Ć���}�|���B�3�d���]=	n~���C�$@/-�@*G��3i�͛7�p����b*�*|�Z�x0�?z|��O�?�g�1�`������z��[�q��㡹ǓBI� j�N�rJ Ka�Q��\DX6���i��O��������x0(�gM�LB�4fh��@b0I�W0�R�k��[¯mT/�(�l��
'��Z��L��OLv_2��,�T"�P�Ei������;�9\�.�f6Clʪ�G����o������a9���h[A(�\��*t�I{{Z�I���1
q���'�_>B\-	Z����o\yẕ�N1��=�����?�������@�R�B���o���sgkw4 )�h�0�-R�J�2�!�P���0-������A���n��{z©l�f������0��$�>B�ȴ�F] ���f�Z+7vj�;��;�Fuqy[�`\لK���QDT{3��u��Mj�~c������w������?+7����������f��Q�uJ�ʌ������hh�ꓫ��1���&�*�D�V: ������h�L�"�'lW^�4/RU�R����e!A�R\����ǿ���[��ɦ�k�,�+�z4�J\��m�e�o��|G��o9��d`h���g~���J�ij��
jFO��J�nk)NG�Qh���B#�y�eք%��(�m��|*ſ0�"{6u��$b�i�7��������}ܲ�i(�y����Y ���\z�)|�wW���M� 鞽0w��2���P�H�d6.7��1� ��40E����\�ş~�ڕ�a��*�}`?B�i&�3h_ȧH�l*�Sr�,��q�&++���N��srH� 9!���$������ �9̂�D��R���!��F�]�JeN?�����$�A�7(N����?�k����h�n�r}ϑ���o���Zv�EF�g��2��%\��������%,HSBT���%h &���F�4(�aŔI��)3ᶟ�cz�Sg� �  �����-姯������n~�u#�>>�vN2���ǰ��I�:jS��.��1�D!t&�h���������ȕ���a5��X�;\D��h^9 �¢��&�͘5�,6��{*�l�����a�v�g��U>�W��s��s�����������Ҡ�lS.��!J!��2��h��dV# �pdd>a�>�n��Q���� �]
$�E�J+��܃�f�"T J
<��1#l�,���-�� U���]*������o����{|z���b��:c�L��h���L@^BmY�ic�C���!W�qxsp����K;Ô�TD��`j=�_��Vy��:���
D�-_8��� �2��,����x��Ji��������L�8�՘����\b��<���d�"au�.����i�DNoy`[2W��i*������w	��E�
�D>j/�bR�!�#ӥ��\jv��%ᒣ��f{7^1����bJ���A$��F}�~�|m��u��ݶ��\ �2�P�Z��z��*�_|�h7�����0*��&}d�q&����g9�R�����"��0��H��/���SB�>��.U��s�k�J�j��F�7o��5G0:@�0��&�����S�z�駟��5s���Kӣ�OK��@�=���F�����'�|�]����r!��IC���|O�n���������2
��k�gHT��1�Hf�M$��O��>�@z�Kk (��y1�25(�N5{������e��T^�S�t�R ^��Tg�L�|�P�6}���H�S���E@H9�e�E�
���E#�|/U�^������!��r�˳�T�>+`\���G�1�X1M����8��+�o)'ļ�:�� f
 �Γ��̖��{�>m�v�x�;�n��A5Ϣ�X�K|��*��Y�/�l�K'���=p�X������&˦���;ͳ�K�o�W^���?��[������E=֝Wr��z%�V��!�kׯ^�z�B�����G� ���S�P�+�`���c����Py
��l��(@�/�<�
x8<v%�3PF�T�*�� ��˴gc�QT��y��R&l0�.�E-IS��wZm��I�F��m�������|��^�l_�{���~����"���VG|M�ևhUȐb�ar��e��]�e��}e���4F�4�I(�C��l������|?E4K�e� ����ɣ������U�{��®hL6���Siw�G^d�T�[��rPx]T�we\�~�!5�.���QP�22)�o�z�~���p9���ȶ���nKm�3��1R�����4��O���=���29?e�E��BjI0oϦN��Ə�c��q�Ш���9��"�ʗ���2���[��q������ᥭ�{�X���lԨ��c����6��a�U�q�����՝��h��U\���JP���`�P��e��j0�Ӡ$0z
{�hz���@�03��d`|B��=�cW�'mbq�՗ߺ�ҍ�zu6=>S˘�!"׊@�&�)s&�3t�^�����P��V���I��xpx��|nsD���0� p%���P���6�W®?A�0�R..�L�&��V�۽�;��ȗv��ΧM��(Qf�L�
���l%�s�,gS�^i�w���'��k�Zov�8�������ғ��˵���Bȸ�1\��qD�Pƿ׮l{�-Vq�B�UI��L4��-�7f��4L�BڽH�m�2l��ib��)V��|�����^���2m?^
�WB/Ko�W|��1�|8Dӎ�'�8w�����p,���zm�IXp��aΔ�ᙫ!�����6�L�U��+''OڝR�dcg�r����V�y����|�y.<o9ζ[��~6a��*��P	���Y��~�O�]�l�/�٥�k�N7p��8 j8.��
��C�L
9i��^�ͺ���[W�t��;���֧���ua8[Ϟ�?6�D�l��ucs��o~����s��X�ڜ��ь%,.����Տa`2�O{�n�5��{v�9$��q��
�|����g�	,Q���J�\h�k'c" R#^_n�枑M�;u¢+�w�7�;���E�F(}�5 ߰WA5I��y�K�F���F^9o.�v�φΚt��5�gG'+ͫ&g�d7vZ�d����0���X��m��[�a�$H6b��T�`�@���Mi9 �8�K���{� s�ܾT0�7�x�;�}��Fq�]���8l&�L6��|%D�&�ݴ�s��a�ĉ]����'��`��/�d�
`<r6ۄ�f"�X��Y�d����,�fC���PM�'���g��k7^�teoz�>m��7հ�u~��,3�&x�?���
�ƉYîs��	n\}o���G����ڹ?0�s���q+�$��(Y���4#�6faw�0$q.�_ 3%.��)��K=�pP>�{W%�שL]ٗw�~��}E��Iwd$b߆�jBc����[��5,��HMh�>�#�N��O�����&ހ Lt=4#�ڦX�/�#�a�j�̆���
�MtS�+�t�v�r��������j�ٷ��/���TyX�
���IY�X�O�k߽z��7�?,�~��0�0�ˆA]d�Ut��WM�L�[bk�Ǆ����Ut	�	�2��ݥ%��	��F�fM	��~���gb��� ��޺��_�������;��X,��K�"3�/1��p����C� �Nk�Ϲ�ɳ����ჴ�]r�8�:�c�����ِ5�0�I�%����|r>Z��[��?]_��ܼ��X�^����^\��k"��w$��/�g�߱�Ex�X_�ג9^�'��K�k[��������rwV�c1:�ѣf�G̈c�>�P��>� c�#C�c	((��׬����0�ٞE}Dm��1Ӌa��ϗ}�p��j��K���'o����w:t;��ؤ�+?��EX	둽}v��E��u��L�C���G�q�Ah��
l�0���^��ƾ���Aʅɀ�[�$+/
3<�i�R^����xf.n����u.�b���rͱ��.tw��A�#���C2��_�N�����S%�X=ħ#}��pMP�zu�3���SLP���Ϙ}U��\�J旡.�&��b�����B�?��ў�0���S���1�en��<++ۗ7~�g��5� 5�K� �g#f�9���r6F��$�e1��5�O�-l�[���qg0>��@-��%�=RO�/29�u� �rl0���$+�"-�t��pC~�����r/�pi��t�G���i\��{������"�P8��k������+{��鞘΢uz;JA��"�^^���OF(@�O����l)a�L 8�$�(�g6S�RZ��Gf��q�ټ3��&v��P��Z��ӟ���w�t�A�%��jD��S��0�De$"pm�R�v��	��GXǐH�tpL��)�.��p$��I��
o KC�V��Aӝ3�ik��Z�7\l4ϖ�B�N�(7�5]���X��H����b��*�G�j������O�N�b    IDATvZ�s�z���ҒH�@M(����e���(My� .��pIx�H'�c��H�֭[�FV�4@C` ������ptp���ݗ_���F�
����W�����Ͳ3����j�r��cƬAlM|51ʨ��+�P�t��������Y��x�?9�uB_D�*�P%����&�O�FXfU�Z��ݎ�N�7�z��-��&rs�Y3��թ6F +	檕ɣ�clI�Z촆|���;o���Χ�U���g+�U�cG��/v����+��D��`[��H0"t[�"����O@F%Q0���-fk���߸��˯�7�v4�a���c*��qk���ct�lڛ�J�N��t�λ��|�����^t�Ѩ���v�<>��m>��-���;�<f�
�g���<8h?;�w[�No@o�Aܐ]�lu�BAM1�7�L�	B5̷;��J�|,�%jW�naGN���B�3ɣ�LڎZޜ�P�t�4��=���n�����§��Iw���$�e�t����սz��\ݬb���,rxjd����2�J� �g�=�!�g"8��!����^�3�d̈́�2���� �R�����H�|�֋[�����W^D�&�P�}��̾�c�Ζ�g���������j�L�G�8��=<j�{���d��#d X���*�E��;��N�^i��Xߐ(�mUך���u��
2��j�9$�!��3�V�|�띭47�o\�������^�����9Ɍ�8�V
�OpH@� ���� Q��G	��|Bl������x�A4'p9� ��|�d��Q:�<��q�k�� �7nm���|����i���)�S��#d��4�����[uX�ס`���I�nN �n��("sӇ�p�i5�~��#B�R�X�@�䎕t�|�����
k��f1ob��p���Y��F�MF��f�����l��jsg��.��zΑ��e|�\h���u�e�
���dm�!7!��.?�PҦ�̄����T8%��l(���:��]���81�}jn�����o���7�.z�7Q�"bD@�V&���L�F�``l?�WG����^�u*z���e���Yq���X�i��&h	W͝ݦ��ެ�����Nb��S�:f]�0m�.�z| X�;�'��5������7g���������=��g:*2׮�]c�M�ڂC�� 3h<`������ �	�.(,�H� ���g�RsMh'<F��fP�0Vf�o�R~VX�^�\����������Ǐ���<qv	/L)ENvY��)�����D��Th_sauE7�3Fᱹ���tM�P���u�>쫜Ƚj�+���������Nx��PD�,���w����X�>��V�\�mh%����;?ȷNN�0�����͎�X�̢�%�wt<㫁�t�O���ר.-�<� ��2��b*���:�r�Vy9^O��姟.5x=՜~�2E�إO��T��\�)'����K����T�а F�PQ�mCd]3*�/��Fm���v�	��'|�W��)0�4��D�XU��Xh	�B������}�5�����RFK��a64ҥ���(k�l��л�)�W*��駟���eh@S��5�+��V��1t+Y�XPJ�/��L��8�%��ZKd��E���.M��hҵi�6+���#O����Q���Og*��Q��q�n���Fy絗�6�L2A�2��b�VXJ��טG.��Gܳ�%կڄf)�O��^ ��:��^L��yKZ~�F��d�J��%�r��K��i��Ź�e�fԒ����4���_�mS�����U�1���W������(�ҶG������8��*�3��=�yU��ٕ> i�Ԯݩ���3f	�XH�B�T��2hb�3
Yb����.d3Og��(?��'M�j����A�1ݲ�$��$Y]@<bay��Q�Z&�m��4�+'��AI��Y���Kz&d���X����������{�El���8G�t�L!:P
��>}
tJ�5�[�� P��U�����Z���08��؟g괛7o^�v�:�}�(О�h�?�PK���ٻf���6���m�č�7._�����d�B�����j��ޥ����?��?�~�5[����|����!�0Sgo�d� ��CkU��r`k���VO1��>gU9�'�,����~��
w] ?/c�����xB�����qWm|+�������ǽ��
H{ݻ�
�
�8��Cn@՜Q@%鮼�.�lL�z���/A���:V�i ��xh�sH
c>�9�a%�l>J͠A �B��Q�{��������՟���`�vg��d`C{��6M�1��L:�!$dF���h�_��> �,N[2�"�_ht��hY����~��5��N2�4��`@�w'�ć�#�U�ʂ�V���0�c�<<$��q&"/^wr^�4L���Cm���
�4c���N#(�����"� ������@�%���g?yt��������H���^���we��2�N��@��?�c�0��.9|I�E%Yc�7����t���g�ۃY�hz�&������[�@� $�7�*
��3+J?��G�M�8��N�^ع�	4�eL����}�2�� ��$��N�%�nR�MRb&���Y)�a6G��?���xf�[]��5k@*��Q�d��2�96��gq�5�$�E�2_�k�|5�Z3R�6uL
t�m�г,����{㭷?�֛۵y�{|>2�֙�
�$졀ce�Cȅ8��YXL��>�?����'��ϏG-G��0
z ��@��I�H F���Y�'�Y���o�e��6r2��b�Kko`ɥ�"�߲�,�e��M�8=2t�Ar���	f1z���F�*"�i��-���%᱙Șq��D<�`c�Xh��r 3x�w`��2Zo޼����	���ٺ_�	"y��o~�y�G�0C�|�w��n5
��5���jև�F�b�Z���2��@+B�B���Z�gON~yt�#x�O��Dq�
�jK���%1X�A�!��>:����
IA���zuO�S�/��W��llTb0���Wb �y�ؼ�ǆ�6���\�͆���Ӛ�~�7�-n=�V��nڲ�tCz���=8��sP�/=�|�څ�h�W�D6 q�6LhQ5�Gmdjx8㋌,/���?��_޾}�l�Z�9袒5I�'�g z�m.�S�%&s����˓�w:L�2>aEB]�)V�Y漕Ǽ�i8�2(Xڦa�c7��@"�D�+J�~a����PY;�i5_�3X�8��g�x3땏�e@κS�F��P�r��/��I��D@����N���?��i��8���ܖm=T"�  ���LTB�G^"\m
+�5����1wp}14���������xy��y0�����1"��F���v�������ҝO���N�=9�{�����G�^��K�K���Ŏ�u��#���H�wJ{X�f����|��)��g#�w��$7�Dx"��l��`�x�(��ۦzĝYd'K���k��y��V�����|���j����g�-ҷL��d�U�-D��� "��^'��օUK�X��� ؀OV��!����?���Cb-��]{�_����W����+Bz2%�ꠣ�{�/tu��!��]�b򳘍�b�����飇��|��>{~����Vs��ر�H%�j�[7��y�bQBfj�"��h�$ ��I46 E��a�1�F�Q`�G6�c#�s��].Ʋ�1�j�`x��͛�g,G�'����s!��5�:�i�)�\�8�����l�姴{J )�I'�2FA�T�*Mba��Au�%_>����|�V���w�{�0[��(}���lݷ�;5S�gY��1�"�wg����;x����q�i�o{�n��w*�o͡:h`�ʚJ������6�B7���D�Ӹ	�a5��@4>&�V��T솢Ǧj��9���w}lLgO��'��I�ʟ�V��0�y'h�p^�A�OX�#ª�ɘf�"�!�p�q d��$�OKg�B�r��PXNl3%k�q2SD0�3�O�Y��g���7��R��Tut�le��'aF��f���XWM��'ϟ>{����G�Ó9�mI����XC�[8#lX2Kػ�ß�f9���:��_�IA�><�s}'�Ӟ�@IH�d@tt ��V_18��qf)���q��ܸ�}�Rn��t�yk�������Han�$y�iN������@݋L�d�q����H�~*#&r<R�m��6� �$���\�e��z�^��������.��}~eƂ-,�⻤����ϗ�ꑈ�~�O=>�����ɸ�U0��p>9��p��7y8&[�y|&�_aV���2�5��J�r�
�&�ψ�XA�V�!�<`GL��7�-�ŬbqVA1w��<w��Q����@��%R�x
�~����
�����"���ӊL�c�t��꫄ �� .�+��� ̘��bΐ�O?��O�+���b�R~�֋?�ỗwטUٷ!�7<�����WZ�?�5b����~��>y���'w<?d�cD�*&�L;�����83]��@{���I��i@l_�|�$�:6q�7j��<����d��|Ʀ3ñ��ɴ$�b�1����j}�p~P8�G��4C߇s 2D�I���G�c�F���>����u,�٥�� p��P���q����~�Ν���B��+Ɂu1Ё�V��<���7�y����߶%�a��y����?�s��X%PH�,a�X��6~q9����,",s����=i?~|r������'� ��]<�形�lsI�C�m��`�8�N���8&�r&�VSo�za~�� ��r�,��F�&v0��Z�-��C��{a�Y?]���2�܆��o+k�˥��͵b��)!�X7~�VAE��ɓ"�K�B̄�� %�_�L#̄3i�x��$�֩��w����N�?}��;��jD �M��� �P+��K��`9�Κă���q���w�~���G�NO����qz�ЙUbq�f��Sx�a�	?b�t���p0:9ju���I^�nx�f�۞����k�21D
I@�} ^��9��?r^y7�-�eg;�z� �u�� 3聉�+A�Ӡ��,��{�2󮴒`��?�Q��SU��`�n���?[�K���WJ?��;�x��q{�=9���V�98�(+�#�oGlڏc�/O 1@ο�_���>yx��ƨu: ɸ8�K�Y�"������pd��u(�~"�MŠ����=�!f����yx�Ұ�����aRcR�μ	�*U�כۻk�*��I�pz&�pFPDx��1Ԡ� (��Ke�w���J%/�,�F�⮘L?w�#�ӣNbs�Pg9Ƿ�~��~��7����9:	&PD&�	!I��v��z����J�JqI_�^p0^��O�z��{�߿�����G��?}�����}D�lǂL�N�b@�[m{�?>�d���8���[tٖ��0��d�·[!99�������#6w)B�7g'�;F�E�@��1�]�-ɛB2='�f�\fv$?����q�{�W�u1:�4M� [��i���
dt�!?8V0�G4`�7���������������lԱ���b~b;� ��'Pob
_��M����3�C����5z���������G�?<|�����O�>o?�?z��}�=���g,�.D�F�t#�oi��L���4�F8�_������0�*�Z����_E���Ǆg+�*{�2��������$
PW��e����7���x���F�3<�y�Q!w��:�bjvO�xE��I���ݥ�b�1�]SF�]�tOo�O�:�w_S�l��B�bQR�$� A�W#��(&��~qyw��	�}
����*�PN����;���-���d!0iR>�裤L���%t��O�_��;���<
@U�� )�"Eq�d-��ŋܒ-�n��^���,�n>��'�s�9sfƧ߳ۋ6�$��PԆ����3d��$��ʌ���q��qcm���bn*ϰ�E��xX��S� ��jB�C��,�{����Ɔ������������c��p|�x�e�yuu�M���4z�=�3�t��U))*NI�Vq��V���H���#rQ�p�9��K�����ڱ �����|(�=N\��<d���HȆ)���z��l5(Z7��O0���(�wvS=*�(�����MwJa�9�tV��R���̄�j(8I%���m�<bvx����5ט��⦟ʨPy%��|� �0Ȩ�z\�|��I8�Q��ޗ��oh�vV�;^��[S�P���Q���.y�Q�*��t��F���W����V���F���aa����j�̸pX��������B5!"0 ʸԛ�`ar�o4��&gV�Q:���|��d��8uѿ?�k�df �R����U2����R!0�+ׯ�~펦���|TmH{��p��0^7t��o�è��7���r9�?������J�ijP�u9@O�����̅��aL�.R�+�ex݋�:��C���ҥ���_�}���+���~� o$;�,,\Z����H=���~z�;�SE���?Z&��**Io�H�A@�] �J�6�<�A��ĭD�6{5Ԅ���B"�L ��'6�F��FE�ez�����z�
��f���׎�\�|
��꾒�Y��וw���Jv4l�ʯ�8D�2��SQU��H�!64*4������߈� @s�K�i�tY:�&lXm��	�6
k	s�hpi�����n�J�w��;�w����x!{Æ��� s�<"ݻ� F�6+����3Q&$9%y���V�O�O�J�%+	5��1��ZS'J�V�[b<1�5Xi'J����޵�!�Ƈ�q�#4�o�gZP i�`>Ё���&��+� ����b9��M�2jK/�z��W[OWۻ;L�|(�3+w�{�ڵ����lp@ێT�LlvY�D�e���L#���B\��ۛ����:��@�4[��->3s��!�P��u'���z�<�J�=F�I��`�f*�V�s�s ������!��њ3�B����[&2e�@�T�dD����3+L�f�g��~�;�{:�N��L��&^�1{u����"~��]�34Xꑣ�]�D$������U0wj�� !�e����2F�"2�&�&�G"?�:��+�n��?���������-�;rqŴ��P��"$�ר�c�1���o�nn�u�?�\��o���1q��.b�}i��Bsqi��Ǌm��Ṁ���_+��JP�D�ĄEkJ�DT̬lIܵ.4��Ż�	� 4����{*
E��]��gP���BKRăΓ��x���'�<�>�ǠEE�XY[����];
zi�^�GL�|��:B��7)_-��m<{v�O��}I5�U6��K/��?z�>ڛM4�Z-������T�`JM�d���z��aw������O,�=�<lw��bi��J�7��n��31=����ɻd�*'����0�2/+Y�tG�TX/g�eΊ�UjY�)����FS&rh ����Q�A=�6jsv��(�X�������%�F�kK�rS�~؜�����?��9��D���ã�^?j�%� �����}���U7���["T`;�(˘�6��z1��?����5���C��L�:ʆ����|眅QH��t,��������n�l:OVT/d&e[���!������#�cKREs�4��!C��/.�3�������ݘ�;�`uk���|au��L?J*�߸�p+�i���4�����09^�|e��~+	�@�����n�}Ǝ��d6q v\m��2y�CUCiO�P��.B	�*�Bi��jt�EAr7��=A��*Ɯi�����>���Fmt���a"�xy'��`��I˷�X�9��Ȏ�������lp�m젋��QSX����hh�ZN9�    IDAT�Yc<`/~oD����ߊ�;�q�%-��ŗ�f -��7�oɭq���L�Ƚf!��`*�3�R���x�&:��ͭ'�����{��Y��o+�^�mBaϧ�aqZ]I#Z[�����vJ�U`���:ڃ���t��	6J>������7��2ot/#. ���J��R��R ��~�!e���i��ǻ[��}����`4@a��l&)/C�H�����Js	�����D#�i,���Ȧl���(��h�UO|��ٌ:�Dh!,�*K:���Ƶpv�R�{�ߝ��/�e�a3�ZRY����:�.TZ���"���B����Y�j,��~����k �4�X���8IB|�"P���vx�����?�̺��^'����͈�Q�A^��*� }�C���Ƨ77���m��I��h �Ė��B��	����eMJ��v2s�%�L\!�����x	��AH�l�u󪖸
#�-L�������0'�����ߥKW������:P�ufF"�<�0B��f���	|�zE�"�
��1@�)� p�Ƀ"��j�j�R���w�G	=j�1Ā,�Yk?��G��w���1mu�0A��P��]�1�	`,��֙ŰV����_=[�<z�3�aݱm���x˳�B����8ߵ�> _AR]�.��n$=Ag\�Y��A*��$���O����:�B�#� �9�qm��� ���g����Zh�}9=������z��9Aodw�s������P�B���m��&�w�3��+���[�Цj�	억� �[6����o�ݯ~,��(��ꪠ�����(bD���>_��||p��1x�d����vW�oh��m�D)F��|zX&���h���p[��Q�2~��0��T��U�Ý5��!'N,�G���@X!�W��%�K��r��+K�[V�5z���88���#�&��~b�_8�$;��X�����L��TQ�,����Y?(5�Q��R$�����+�G��lt���ٿ��w�O����+�����ӟ�{�Ʋ �j��#, �;!r|����l�D�D�;�;���߮�p}���P��fŉT�������IT:|3)�2�4�D�"M�;1.���7�*k$�p������O��;�tB��4O�N�YC[#j6����Fw|pxq<�cu���B���Ek�Ҽ���X� ����d� dh	��W(����iC�>؜����~�ͷnܹmm����\�)(�_:e"���~��7Oݏ�Bҟ�����o>�}ﲅ7�V
ƙ�a�8�8� H��{�ck���ݯq�p8������Hܬ��&�/O��1��h��Ve�&�\$�J/��}���9)z}���J�W�&�M4��L$��J%������bsfi8�;|9�L�+ٟ��!%�O.-�\�eɨ��"��5�Px���%��`�t{9ԅ�~*��*�N��~�:�1������Q�;J׍K����÷?x�>N�$��(aرg�b�����������J0�ѳ�[�������9�%���!��F��R���R3V�@E��D�Y�>S6
u�:���u���Uj�H��I%�!�w�4��q�q3G���&�����+��֮`6�N�����~0�:Jmd�w�9�,gw�y7e\�^ar&�&]+U9�TNF�	$vd`E����+/����������;m�I�V���HL(Fl36&� 
�P��Ս�G϶?f�g;<��W�
�6�Py�(�dyWx�vB����C��Á�#���;���6aH�:22�����&��&d,���eQ,���\��om���U2O�U�D��Dc� ����n��]�G
�.�
2����.�,��be�äH%J����7�'o��-�����O��E��ٓ,sOd]E�dUG��!Ը�sc1L��H�]"���nw$U��g;�m<~��g_y����0��@�Ԕ�Ҽ��	�<��qG#�+'���A���G�gcCC��(>(�*� �Ci�G�bК��?������^�y���j�>��1aA�8������n�o���s\V�9��:@3!���0��ՄH�q��HS�Š��$��g��y���4����������?��9soc{ws�L�:��"l�$��H��1B̔DmUN�����<&^v�ymc���~;�7��\�"d���f}���L��T��������!�Z*mBdvz�vg�	C��㩣�WRq��lon�ꕻ߻~���uz'��1���K�B���%�H@��`��N��z�s�� �����2���Mw��}U9g����TN����g��E)�.�����ʸ_�r�?��~��X�����@29��N����`m��8!S�[۲s�x��Iy��'g��Y�_m��k�$�#��m�����ɓ'l�|U�r��%�ouu�Ǫ`�/j*)�ش�H��޽{�H�,�����D<r��ݻ��8���� ����K�-�a N�QOU[��s����������<;�uS{|W��K~j3��k��"k:vi&�RB_����۷��\H�L�"��ppq8䮊 Qe4Ak��ʕl�Mw�O;��׵�\�c�����0�jS�uA��l��,��yq������驛�u8��U$�ȀB��� .mP��` F���ļ*$�(�>~��O���w��}�]w���2�@������U�2~Z��Cyv���b���z[���{�O��Ä'b���Ԡ�ߙ�ن��8q�S�ͦeK����U�9r�`���J#T&h�?&���I,�G2'%i�_����KdA��=��l6�]ј�����/��+fK�I��:����W�:���K�u��y./-YPh��9+����LG;��:������/���'���Q�y�A��;��'(������w FUl��OHyO�ф氳{��mg�@�V%�@fv�\UJ`5pj���������Vwo�7FL�[o�'��K�^�����{?�byqP�9���IT��Aڤ��z̸g�� ����:����9��a�j-,��V���q}X����~m��»@ނ������'�P ���� N%�x�g��|�"�����U��������͛7�ܹc��G��T� �`���#�H3<��?����X�f��T"���GB6�G�l��J/b����d;������}η��A0�� z#��h5�R�q+�TM�s�䆒%�,����#b����rL<1�ؼZO�4	�b�������W��N6�1�x�/,��27��?Y-�m12f�����N{�~�p 9�T��Ы�惒s��(|A\�j�6\��� T�(�J�:��U����?o<{�=<���]�s��_~��0AS#X��cbZ��JMp� �	�����h�6�����g����tI��S놤�A���S��*�xa�F�Ȓ�EB�\D%������<�yD��"3Z~,>��E����$/�� ����
��5���",��p��Y�S������������ّ,"�C��]��V��Ks���g- � ��&�q�L�D58��J݌3+|���	I� �6 W�%����F�EB�k�����>�Q?۾�.Άd�d3�#�!�~Fu��8&���n�����jg�= ��s�f��*o�g�ۀJ�!���B�T	�M���@s��D��5�߿�:+s���f��0lr�.��`+��W�(3-c*��z8�{<%�*K���w��rRo�xn�:U��\|!Yj�������}��Y�D3l��Z2�PȈ��#!D�Jc)f�������a���IR˿��;?x���dw��g��t ��y*"f�T��qX���'6B�z����aݞ�I)�����������jɻ�����g�NRT����BY��I֊�ëCjK����|s��`6���i��T΂@�R8l�tL��b!�2��ZKWVg�._}���6�K�%ݲ��W�f���s٭3��4����G#؟}�j,� �.�+��l�2(΅z�@�=��1w��̊�)���o��/>{�72FaLZ+��@�a�&�d���uo�����'�o?;�o���'3Mf,�����p�k�y�3T|�����85�e�m)7<v���#��FE����\K�3n�EsG�$/;�h�=����!bEg#��I�*G>�0�ycv�k�Z�|x����`���?[��Y/���
hf"@���y2x��2f*��mZ��#~xzŝ��*���͡L8H-�=L�O7^}��?�����ɓ��a���̮ޤ�.�S�5vdmS1�q:�m<�x�`{u�p�7<H��Q(�|5�%�Zc
�%�4�u�1�`�9X
8�5&����8��I��䪴��dD
B)ۈ�h#�mt���VMʵh��3|��̆�b��B�����D�`���Ϥt<Df���e��1��^��.�)8c�\Aյ�:�a��3������Y�H�*�K�_�I4!���w�����������`@+47��8���  G�e�:6�k�^���?�k�k������d��dsW�19��F�D���t�����L����'dp7�(�'�J&)r���٤���!����`���1��rzu�@"[e�~�&S��<��D���8��<�<���+iX�#[�GQ���]� A�* m������5fw�w���i�T�*T�ܫ���Z�y�[�~���߸<uJ�u}T���!v��H��ǽz��l��#�v�ߪ���vz�\��\�V����cA��J��!�V���Z��1n�l�L�U�.��	w�0|�p���e".���)����f� �����v�N�O �w�7z��:����ES����)|	���`7d�k����G�2. $��"a5����]�j�&�M˄X����S�n�|�׿��ͻ�N����6�K�U��7���f����L������7:�;�';�α�YS�aP��y�̸�l֕��%D��:�ʃ�x�a!�e��ĥ7<��R&.��5l5��}3m�!p��ګ�8m��2���O_��꥛�����~c09E���#pE�6�Zݫ�#c;�,`qS�A��BgP-OKI��9#/���щ�3�����{7���|���)�j��F���`K�t��,���F\3���:���~��I)�U�>��ٛ>�"�E�p���Q'��*��8�g����ݐ(�Y������X��;iq�Ҋ��I*o+J�1���/������:!%z֞��t�	�u�f�,Ӈ4M�T^Ð�_m!P ������>�	z�i��)��5��j_g4�R�+��J��Wp�������͟�x�i#T����[������������*&LO�Q�A�8��b��'�t���{[��O��nn�z���T��%�%��#! "j�4t����-x�i8�ւs(��f�1�END����k8���`0#��T5�	���v��psa���Ώ����w䇟����ļ�N���˲l�o&7�
aC�C� E�F�v�~�\M���X�pAY/�����o�{���KWV�&$f��Do'����qz�����i�!�}&g��>����s��/Aş|'8���L�r�ғƺ���`u��dko?�T:Vƶd)z	 ��ř�*�01
�ɛY�$����c"ɚ:�T`�.��R�<�#�0ǋ��B ��G���Q�c�,/���nޯ���#u���q�t��Q{in��1b�L`32ی- X��������"�~���
{���0d������ނMihd�@�Z�wj���s�~���|��MÕF�0Ű�D�"UG�^`����K�A�~����o�}������oI�'M��[r�*t	��Wd?�����&���Q#�w�${�K<��-̮,(���V\�+㝘M�����ʔ�h��&���G��������iw�h�7wy����L�L\����u)�*ΎR��r�k-%���:�.�$:���y/���S[�2枷������?��O�߼X�o���\��R���l�0(i�*7Y���X��?����Bg�����|�"wc��e2d�1k����l=�"�ɄMg-%���2@�4���]��<��iI�iJ'��҇*- �N�2ib�@���,k�.߼u��������__�h:j��>�J��D���
+�t:��� ��tߝ�2(`���d��T���M>=��z�KO"���	ժO���O�������_���>���j�y�H �jgn#��	�8��m��=~@��X_�a�eɞQ#x�I��א�S$W&S��v�m�d�0Վ���Q"�á���>
g �"	p�(��=�-Ѵf���uA@�w�56��/���䋬I֔�&l�����Veo��	�$�P�����}w�x�!���( �~�v��+"�f��?���i@X_!�lB�f}l����?���s˯ʣ��ؾ89D>��T�ǈ�Z-̛dH[���;���������ڏ��?{�����~rL���1H�M5z)YiJd�VcaP��n�ݝ��^���8>�k�=qFTC����j��҈̀�ŘD+h-,5y��X���(��,��wM4���'��!�TPѻ�:?}�\;�!h���H�;����" ~: ���b:Q�g��+���(O�����z���s��O���R�W^4�|���C)f���L�Kּ����J4�<*�w0d�x�ի�y�}�+��	
�����;O�<f�'0�</��>y���G�]�������Yd�U k�ܟ��.t�|�8��R���t6=������>���/�����۔�W^yEt٧=�o��QMU�pX��|�GF3Lmp���v�S=Yw���T�S�tD�T�n b!ӄ1�t��]j���+R�fC����Ϻ �3����Y	(�DA��Є���GV���2pnj��;�L3(C�f�2֥��r�����B�O���A�K�t�HԀ���_�&��@^y}:7�8���	�jS����UÀw���Ei�A��Du�yGS��쮐��%��D-s_� ��J;J�K*yљ�`U ��T�AY�SNP:�S���x'q0�vx��ԡLS��pJ�#���J�Q���y º�.��m�`B�B��.-7%y�-�+���y{s|д��dZ���z�n�x}�ִKM�����]��lN�B���ar � P�e��0R�@�	��5�T�P���q?��Ƙ���j3�dS��P��
���D2����*���c�\h���k����C��'��k����zc��˗����x��Ť��qm��h}��O�N�Q�ll�(��g���t\qfb�j���N\V����𠿶5\�;�9� �#���������[n.
�S����M����o��\ʘ9��g)��2nz�p��Q%T��ͤr�4pV�|�E�E��Q{��
�`޽{�����h����e���Wt4V�H'V��NS{��aw�����|�#�[��K��I�\���C+�ॅ+�hb��"��F�c���f��,��V���ۦ<-IJ+ �r�
��&P/��Rt�ui���g�UeDΡ��+sE��8���]:!Ō�l�� vGLn��niD�!8Y�p2�b
�!��1
ȓ3߮���?�QFͻ.�W 5kzmc�r�/_���e8/C}�{����׮�Gv��JV����3S5>I2�K���{�l�Z���3��r	1�	4�$����b|	��#.R�O[�J�|�S��8T �~H4�P0�*�~^g�e��ǅy7�ãnK���.����l��k���Yt{^oY�Kq:<���������ʓ�|v��µƥ���ɍIϖ!fn e������:��|b�wƫX��Z�ҍJ�����hG��n ��6xh��o\��������V�X��#K����� "����3��{ku�у���Í���k��S��    IDAT���4S�GD�jh���`����gY�.�%�+i���T;jc"buN��!�4V���7y��;� +ш�A��q�v��f5@�Ux�i�Е�������pi��!@P���	�%V$��JEB_pnz ���!Q��D���8	���(�Cs�U�(�ݍo�|���YE]F�x���|���I}�/�.O��2":TUW�U�޺�G5g���:;��Ov�6���~�T2L!��AI�>K���fkzʖG��Ƙ��{)-\"��|0�_0%?���)3Y�;�2*qc|����G�;��$i	[��v$ç� ט�hE�3KWi������ӯ���cN9��)F����7��-�f�|	���c4�[,�]I�d3b#����q9~ƨ:�+��]E��H��6����'|�Zk�'���wc�A�!cfB�SũuE�&U���y�>�y����v_k��k�`,)6�c|	ʝKdZ��6Ѱ.U�͙��G��7���@�Pl�k�c�sdK8��f��J��d�>i��rVވ8W������m#����^sr�n�O���]v=��z˨�|��H0!��6�#��]��)U��p�����Uv8�ԼP��x5S���p�d}�7����p�b�w:�G7�fTo ���c݃g����8�m�n���Nw�u0�Y�+�yr��FZfZQ}%t�����T�?a�����ژ�'k�;0��������,5H�qg�7V:u!w1�e��}e0F���'E�d��d%�������d�q�W�4�V&_���P`��i:$ux����\�gu�k��>`bz:X�vF�P��MtT��R� b���䜢�ů�������5y2D(`r�D^��'$��u�Ŕ��P��ph�_�>z������X�N�qC�=k|*���$��>�U�	I7a4�� ��'38��65�l������5ܩ�"d�s��Ǭf%{T�(�h�
s�y�2Mr!#Pa�獥Źei�[ۻ���]aC�@#���3�08<�IP��
h^�LE@� �P�@4�#��U�m/�ly��溥_�fk�Cw<�������V?�V����G�0ޙ2AM����Qgo�����#�?Z�l���D�{L�Q&�|�e���l�9=q�jX'q�q��o�N���R�$w|ܗ���E3�h1?טo6$Y��>!,���~vӌ��t��10��XU�h�%Q�af�����������#�l$*�<3��"T�[1����HP :�5����QpǑ��v�>#r|+H�Yi��0��������>�����8����44njm?�I
!���lYʩi�6��/=JoO��j�Slf���4�;�nn�=�(�uaI�&�*E�6�FLk[�T���+  7JT~��F��SL��� ��~p�T�`d���㋳�a�<��ھ��q��]��X:MĔ�q3T2`(E J%�(w �O����g��G�f�'�4�t������k�)�g��R���wv�4��Ͽ���\���z��*%�ѯ����9�����������I��^[D-� HM]���며h+���%eQR/���цKȄ�/Ox���12p�C�,��u��^�0&߷�d]�PT}0O#�U�*M˛��)p�>o��K�^���=8=hl���&5����B�*�U3���
V��@��
�堞5��͋^�l�� ���"Tp]dF�~����:;;l��ַ����xiE��O9!��I�Ll�Aʓ��D�b�;���Z�˯�?z�~�ݱ�������Z�GB��	���ۈ���'��1֦bTv�@UA��M��z�1?H��s��I�v�X��l�dz?�7|�)a0�gg��/�5��Nڛ�����/&�g$��$���/-�k���l�0�ɡ#jFx���6�`��`��Q#0NO/�_�u���_����-Ġ�	i�I&��8;{���G�K7U�x��7��受��d$M��a!��B��ҿ� .k�;�����>�[��_ۗ�*P!�X��LF�F�l��<�6��� >��
2~Y�,�s�ޖ�(-R�,�6+E`��P=���k���15*���U�{�s(T�[���#'(����1�N�ag����%ir~(�~nnI
UX�,M�H� �nKI�
ݬ��XXd,��*�G��f�P���$�;�_=�V����/~�ѕ�T�ژ1��)'����쳐��Ө�8�l�ҭ������˓g[mMD��H8�$΢��ńAM�˰�S�/Q�NҬmwX�Ľ���Jm�ޓ=�N�z�+J��;_R'K��ϸ~긿��a.��PC��e����K+w��:�o���K�M���P@T�U����(���jg��LҊP;�.���Q~*�? m�
��s��r:{��.���O?{����s��H�Co�h�!EJb�&�B�@�,g�lo���������׷�̗�����d�h�?��(44Y�'[ċf�����i�M�)rg���
׋9����)v}�B�~KT�_]P&<���� ���I���/\go_��t�cwo��U23�ԁ�nP��䍔�R�ۀ\rU6tQ�y����G�vP�ʛ��D������uRk�e�r}�W��n�����^�l�Y�,a`�����^�m>��>�x�twmuogk_���F�Q��u>ɰ$_`�%�]������Л���͞��� !�kGCN�D��g�*���ږZ}o�ѷL��y��͹K+W^�r��tН����1Yq�	D�1�#Zӑ޲��*�q/��`H�����,]{�S�N9�9�Īޘ8�@O+-G����{i���˿����v�{VLn����;�4����Dׂ���vI� �'����N�������ƣGk�k�{r��2u��0^U9���}	?�v��)֤���8�F�"�D�i�g��[��	�ۉna��g8�D�N���Ϝ����%k�"K+�ͩ��ӝ�Q=F�g��6Tt c� ��
t�=r�i��R��L�.�(�>h�	�Ԧ��=}Am�����i��}g5g�*LPF=�������S�.�+�̻�i��@EO��85ՙ}�2�(䄑3QnXQӜ�}��e59�5�_�RG�:}�*��k�2���@>G��TO:L�9��Ǐ�<y����� ���-�����=�/�8���ͽ���������o�8x��b��L���k�x:WWW��8ˎ�I�2�`�+jS����S5{� Ib�҅b3W����z���V��i���OO�\���rY[`ʥ��޹�ڭ+���$��@qGVj���bs�n��!�Q!J�~~V�F2u�_����`/F�M�)f4~��W�����b9s�Q^W�! 6���;� mmm���E8Q�͛7ޖ�0Mn�qG�`RjV�Ou2g�ܹc�����{��mw�P�����}���w���W�ϒet��i"���� H��g�G`��A�EL�Ί0��Q�� t����M�k.�W��L�(\Hģ�zD(�[�Wi�#C&�
q�ŉ��4ɋ̆��c(8؝��ٱ����4�z���,���f�6�cx����Ĥ,X��D�!�1�����Y���7)�A�_����k�5��ˤ2r� 2.�Ѐ^���p�(�QO9&��&�<΀YppT�& �0T�X_�W�!`C7~�� (�]w��[P�P:|�O��7�$�����ᒳL^L���=]�^�{�������Ť�P������G�-HB�ӱa�02lz2a�G�׸��_�"<3A<�Ɍۑ��1:1V�+���q(��1����r3�PBg�sqǪ�X}'����; VU�̷���&���i�駒��~���qQJ�	���ݻw�%`ش�BW�����M����\� `�T���w�ݻ<?�O�����D\��Z(,�5Ğ�fۢ0��o�no��n�
g><�
Un��ȃ.5Nj&a�"?�M�ǲ��ʂda	���D�@�h1=�r�
G�rLO,-7���`-�d&\��:׾,eIq�j���۱Y�i*F$ �:(Z(�]@Y��|s�#X�c׆��W���~��������� �6���W��WЩ�`ɡ:*K�
?5ދ/�¸�:�x������x{��j�������zu�~��D��#H��Ӥ�Q�C"�D����v�����+{��U�yP#� ;l�"3��X���˶M�A�� ��5��ω��{(��$�^��6�6��"Fz����#0e�X�dnΎk�M!�5	�u,���S�2�b?̀6f��3�ͮU)lV�6������n^_X�ߠ�N��|�2�Hq1@؇��t����g}V�=��=�76��R
Wݍ\R����3Zqb�F��1���G?x��[K��ڈ�O�Ÿ������0U#��Mj�z><�Y������vg���&8<�n�'7
�L�p	�e���C:*`�$��%�&��^�}<]�E�KZ)��+r������X͖}��m�0;5N:0/��Ib41�H�P�jZgܲ	�]o���[;\X�==k�� ��
��,	����˅��q(d��נ����C�	��#�q�ԀC氳�����o����D��$7���>��\c�C��V���!5>C8�q
ۆc	y�����o��>�h���qp�a_=xo�2�:T��9M�p�6�h��8����G�>�$g�Cu{���@�Zx��6��a��M��9+!���lLLbd+��c���&a}�\&כ�|�זkÝ���v���q��8��^���\�~e�"N�*Â6�do&�J����f�S�'i�Q
`�sd��j0ReDp�rv+����������'�@�w�Jgc2H�$W��H��S�N�?���{{��<X]�쎎�1�u�.䏅(���PW�Đ��\4V�Ro ��0π����%�3ӭ떣W3i�TU����$G�y@�3l ����
�	����4���*�]B^���>�<��6�� Z�j4d�g���?)�;�]	�Q��3���͂��60�CL�O����z�s�Ғ�Zv9f�[��|�ُff�/��Q?NAd3����
�� y�����@fom��]�w���l�cQÈ�*{�Xws�Y��rv��m9J`� J� ic�e^�w��N��WKQ\��t6���VB �t�S�ꢑ��!q)��$��]�<Г�ǘz����<Nx���]:]���@(���B �#}�������݁�;�	�΀t`X Y�8���P=}�zꢑ�a=/����u��k����o�<6=ړ�! @�XH���ȷ+��/i|I$,Q�G�!K{�`����տ|E�>��}�]��D$��WfF�|(0B�	�b��l��'[^a�F���G�{#,[�auDK%}'��Fݲ�$����,� y�+��bbF��yd��ڠ������g�{2�����-�@�m�����e�`(?�
ߩl@W$:�w�����D�%��G ��險��1	9壋�9u�{_|�������1���1�z=�%�hFe�b�"p'#j�૯7�}v�#5�4bfq2+�<�����-�N9�-��p��`S���k�.n����Y�C����k�!�>̖����)=���[8�x�5�EtP�3�\V %J :��*p��EY+�9y����X�����-�E'�B�H@WYc���&}�y l���AH�X*���;�<EU@+У���a�nV����<V{��/>��R+b&�Q1���4���6r!ODgQ�6�{�`��G;�;���w��{Y.��~�<�૳Q}�,j��m�'8"�i�) bP,�I��F�"hxN���)��z��(k�L��D�샐�}�����L�Wm�yijb�vT�nO��G�	��aZ�ౌ�M#���z��g�@�AYvG?�����O�@8]���Ś��=�2��n���5��9�����~������g������v�͊�l��P=�Yߊ�=y�����`o �z�n�����ƂY3l5>�y�1��{#�UR_�sU��H5Z�������2-�U�`%�նo�\���/�_�{�R��c��C���;�5���1�}�
ٱf&��;3;L�+�gF���@D�	M������/��~��*����G�����"Y^�� @zj�~�����o���-n��n�|��W^�J<[�P��t��!�8��>?E� ���4k������~�pW�-�gQdoR?�S³�'�IR/�!�	���@p������K���Z�z�l	Ů��)��Im�;+W.ql�u
I��J���gj�A�/���7{x�k���Z�\�V�̮��,M�,�.$`+v����j��� �X��S|���Zј������}��ݻ/[�Y��S����,l���%����G�~�'9Wm�Ưb�_���wo^�8:DK�BR��wJC`Q�n�*Yd�\����Y{�����󝝑�]�������NLَ�d4��E:E��yŴ2Q'��#<evyi���ۮ��8�M�u⒏���f�>&˳C�n����P$ӷ`$S �Ԃ�Y����_\^����<:�Zwtzl�"�a�5�x�9;q	�>O��&@Vn	t�� �G�𐠊� �i�%�<r���9j��Ѿ���?��Ɲ���a]�QkX��B�ɤ�zЇ&��C�ͺmN���ǻ��Z��}+��GUT�)"p�>Ed���A�!}PU�5XJ,)ً
Ϣ3��BN����C	�5�@cu�x���Z\;��֐�����0I���8�3��:-J�Z����n���0< Q�FA�rD�,�t�(�I?�9\x�E9�be\��me�X����;�F0�ݼy����ve�J_��m"��F*ॿC!�*����t�����;m���xFvӆ�Q��T�T����[Wfh3r�#�h� {_Q>樬�c��0yH	�kO�cj��]ə��*R�I}�UuS�`.cm�2S�r�	�U��;U�����c�5���U�[~g	�f���CTe����ѻ��TC�V̅�T��3�$�u�h$��t�
��?~r�{0���=��ʲ��
���JǒW�?��>$������[=kw�;}�(�0�Q2+BO�?K�< ,!?q�R�qW�
���W��&��zhR�=�	p_��T�VY���Ȝf%Ί9��s���	�����hw�/���6a����3ZV1�$���3�0��
�`}*��8Q��p��Px7]�?�.��v��"��hd�Bq���+��_���7~�}}�5:�4�dNC��,��:��� ��o���]�Y����f[jY�fi �d�Ī�;� ���zg�+���.Vwb"�p�'���I)e˘��}Lz#��Ƌl�#�E*E؝��'D���F>J��-Of��k뇛Cf����c��	5
&{�z;d���WPu�����rT�/o|v����
�İ�(�����ᣪ��Ņ2���HU�Q)��~�;�y/fV�h��
K%}7��)ϣM��*j��Fg�ћ#�=��|v��xc��٘z��-��`�Uӌo��6�]��Z��l���>�����1�������(<��}�ٽ{������ZH~���1�nW)0��x���u
��ϕ�J����I����~�;>��ɓ'�z��Ƀ���o{Q��W�w�ܹ��߮���������K�\����a��Qˮ�W��i�1���]S�+W^��y��������[�߼�Rka޺��wF賉�hl�k��	�3s"S8b�$7$U�����*إ���M�/Ʊ��^u�p�����qӻ���}e��q�P�������Z���T��?���I>�u�7
h�� kXy�կ���[Qg��w�X�X@S/�p�K	�tI]/�9[qQ ��y��nL�2B�v��-|�4Tߴ�SgT��M�1��VH�?k��m��������G`���������{����&�{��Y9h�g$���P��C 6��P<�tH�g��!����E���y5Ύ����zc|�ՋD�Ѵ?    IDAT���Q��A:6��E((�?,YX�o5�KK�/]�F����`@+Zz�vv2ow{k���h6���%�!��j3[����1� Ш��Q7"�M�rm0"Ҫ�}���PN8^��0���@��hɄ:888�,[����.��X���O~�_���y�m��#�G���G�AU�� ��BcQk���ρ8��%!�p�D������b^Nz�k'Lʵ'��������[�4y�h��TLE�a�~��(�>�gA*Q��O���P���.g7UR����/
�[�x�. ��̣inloo&	C����gYsGYY7uq��5kg�E5�	5�>�P;�<���v6�Y�yr`����m)k�ķIy�%�J⵬ d|�^
�ˋ�W/k2�ɯ@
�è;!M� W\��M
/�\�|���@RG��pb��DWf�[pג�2��,��۬D1)"SȬ�rp$'b��^'��'���5,��:����y�W5����~XZ95�tFR�����"���0��5ĹC��D�ϓ���o�����z���2��d�(�o][����bCp&+XrڊRF�>���x��b=���w���:�;�G�#�61Gy�QO-��,x��f��FD%��� E7�S�q�bт��}N�(�=�2��I����8�l�W%���sn!y=�VxϷ��ȉ�QL>�n�%n���(wv�9x����9�/�)���Wn��^m�jM�B�l	�����D_�>��Up;���*�T6�R��vM::T�F]��^�`��K�7>��'o]g�޶sRHe���Vfk6�Uc}6-�4����Xx�ɣ�=��!d<�*L()�p�\�r�Q��N�s�E�1h1��:0��	�nN,���//�V^�X�-�Xj�O�Nk��1��o�4��aq�#ef�� C<�D�w���,���H��>��-]��];?���$K��D��wU۬�AB���[\h����ݻw�^�R�=*��EbE+��O����]�i�c�?=}��_���z�|ر9)~�T�PF0��X�te���5qt��Y���9X��v<`��b)-���:;�fK�B��NR͕+s��&/Bٚk�/ԇ#���\[P�<��D玑s	m�������Ҡ�����Ͱ�)l�i�8�2�g��^�xa��y6��%���2{�hw{fث�}3ӚKP����Wf_b���a���X�z� @����ݎ��;:���m�[����{��E��&
 �p��?
)�=���o~��{��g��;�CbN��C��*�'j�	��?��:[{�ݵ�hCP;��n�HhE��uq�f`L&Ѯ8���|}�Y�N�p�~x���Ķ1�G�b�D?��[XZ^dk(*F"F5"O�V���m~i��pb��s�7�̾�G���16d����f}a�J��������\?���m����d
���u�
�0��U��@
�]WO�[�?�G)�=R� ���L�������^���O!���6-F�>�2��BkyI����A;����L�v�ZfЌ``��d��j�T�l��X�},��|3�L5?G$�3�XUs�%�MR!6*pv1a���Y�=Lb�b�-><1�-N�L�)���:��.d�~֚ۅ��`�jƿRΞm��j0�n�K��KJ:%����f�MG*��΀e� ��Y���;p]�o�L��L��:�x	~#��?���s�~�!ڑ��a�����0�����af$��´��Y��'zVb�NF�2
҃3�Ř3���a�(h�J�)��'��A��EL5y� W%&PYyk#X��Rf����~v�%��BD�j@��o����-�C����9�����6�֌��wZ��'C�&fbC%�I`�^G��|�TIQ=�N�#	��b�ҵ�p�^@.����(|��ƒ��=���p6<"�M�7����sa|�'����N��8'U��D��Q��>9�u��?ݻ�xg����l�cl7��!_�xN%A�1/���k >���1��r�C����%e=�:��]�]�̂�6r�K��L��=S��5~����b���-�$��%� ���ԥ�������ʖ��YcC����g�`ߏ���,��`�4{�3�1QA�ʑ��263Z0
w*�, �zXa8����@$#�+���-|����yc��h�o��G���"FJ:pqf��a��]���ڃG����ђu���X�#F��Y4_c0�|�� ��R��_�rQ���pF�'e}�!�_~e�͊%UScR��bh�IWg5�`fA�V��"1b�#����.(��҄~�x��ޛ��Z$A�aK�='Fo-z4��U�����L.$�@T�q_�r��B�xA��v�
&^C po����|���� oV��Z$]<v��DP���{h�o�~=�~V:C+��EiN:&@���@���@%��N6�Њ�zΥ���zg��-���F�HkA�6��-C�����2�_si��6�3+�湈�9{%W�����7ٚ[ �s��_��[r<7��4)��`
V4��n��g7� d�'�O�X�E�,@V�
i�?L-Xl.�?�-����x ������Ϳ����J�����O~����^ZYhR1���ɛ)�@�Ǹ�T�c��9���>C���N����� ��J�B�Q �!�6�CР���8.õ���dnD�V���L���D�L��aMS��C=8̜P�O�f���C�0k��o:����Ӎ��8Fg��斖��O��ݡ`�,��c��R[��)��2:��թ�Ca�j�)� ��k=�FZ��:06�����+���G�o]^�������B���sf=���o����m}}�h@�4�O?��G?���l�S�nCm	u�س�K��	r�o\�&f�p���q���ݭN�f�t�������g6J`[�(�XmI�J���9̑��ڝ�8yqd�����zF��	��C��؏]��V)�Y�,C�}7>:@J�Od0]� ��,,6f8�����Ϻ�L�͛`����ڕ���+��bg�!��?�&�ol�*a�$7�����Ź��J���k�MH|�=���@��r+�ך3��[?���0;J;��i�ɼ�=431Y^�>��'�$?�lw0ʯ�mna��L�p�1�jU�_�
5$Iyp4��	��8�9b�m���R�)�Z߂���?��&,�JK�p��AO'�)	^j��9�]�5"�H3R&T�ꇽ����\��W�
E�$Y PJ;�����9=G����~G�����~���.I�n/h�0�Ӻv���������|��2�ou_t@�m4�9���*�-��,^�׻����f{φ(��qH�
G�򼫁$j8���"�*f��̠�(����XP�9�� �`�r*�S3��X�	薥�R�
��6�h[�s	�9I�4�Q�l5b|�d������hb�ي���e�q<�#?�׎�/*?�ͻ`B�a� �@]�.��/p.c�Za7=E���x�W9��o�NF�[���>z�G�į��ݖ��x��B�X�BD�3���8����G���G�?~��|k���WfE�I���	�2�cXB�f��L0;F���)\ޘ�&�J�`b�x����N�iYDh�p�d¢���L�Y��Wq#���,�fԳ�˙4�6*��Iw~�Ѷ��/�0 �'j�%ٓ������*AŔ�\�3��R���a�_���p�}�wX}bW�C��N�����1������ha�Rg�����K�G"���zJOG���$�6��χIw�{����������t�y���3�U�E�;�9���u&����F��Ť��� ��f�^�.Aqc��R�MR7T��!����\AF�I�+sw�hbDv^h.������&t�Ehh{���Ӏ�_��R��B%��\8����4p�+J^�I�������rv��Q� W��*q߹��Ha���]��ы�jP�|N�R�Mw��z����rǹ��7�gf~��kZ����'`��+��n��v�}����|ocm]d����z�ݏ?���[�W._}��	��k��
T{m�����m	5�vw�9_g���y@Y��>^F��z�s�{5�Ԫ��U<��%�YxF���\s��@��gE����� Y�tY�T.����\�2x{咼q��[75F%B�^��q}��]�R�P�GR�����W�\}���CU���ٖLe�ӱW�;w�޽qy~�)��#`�V ��Egt�
�����(ڙ�Ȣc��D��Yd�e�����)�U��年V@�O�UʔG�݌c�0ή=��	n�d?�nL����e����/���kPP�X|���~�g�F��+�j��9\m�OǍ�<��0�O����fy���L��I�FNa�s;�(��8��@�ꤚ5��ʹF�(,�W3��A����F���C��ݪ��֘���t���^�@L猚�r�w�Nf&��{�����nYa������-"pD��C6��HƯ.�K��X������M���6�g��I�	7/<"�f��,M?{�5'ɉ������}]�S�.�X��f���B��L���9Q�NO���5��5p9�.����/� �5�x�#��P�j>��(���j�jCc�����1�2�aq��ɰ��DH�Ⱦ+�-vw7g'-����������l^}�أj�������H���Ȁ{�42��}_'�8`�kh^���I}�Hl��D�L-q97�n�l�}�;�d�rh9ߒs*�VR�N���� �*�}M����.~�xŅ��ñ��oq��o��T��J~���S�#G�_t�*������.jU��M ����X��IQ5��xl;_�����~�]���x0>�ַ))P]G��΁�`Dx)'䷙�;М��>9�WYD��t���#�;عv�l�$^f-���n�O�Mn�/][n�ח��5����g���.ۮ��-l�r�,-�߸���g�9��q�Pi^}��	4tE��
@�a8��)�������8�|D�D�re��Nh���-n>���Ź˯��e�d#~�`��?ڵ��M؅&PS�;{sXLe��ް3���'��YO|}�f�B7�;����7p��*AW�f��Nu[WSˏ�I�9�����ZZ?!��R��hC=��G5�'��p�zwgsey~�}�hٷ��hf"�V"����4�����ё��E�_���W����im��4ck�������drlM�(�dA��$��/	��m��Փ�c�2�X��z
b���ameȌWX}���c8,EZ�rs��K�Qo3��D�HQ	�O��
��A�3����z��O��mU`�氻 �x�Ո��$<�z&�r5Y���蘮3v{�I'�+��\��C2=�]t�2��]�mel��`�B�>��`�Z��.Z3�/-��z��<���A�Vŭ{A�gfΠʃFGf+������ɫ��R���O��:�k�+6QQ���jKi)\+��U7�:p��	fP)�U4�3��u�Ln�a�f'?x�ֽW���xw߬�=�j��@�k^p�rYY(�OD��Ag�����>�>H����*ү����gD���[Lv�tu������Qs 71[�a��5�Y�ϡ�{r}ş�!cYb%gu�C��^�J��8<hw��-�?����̂�8�iG[��"N��5Pxxz��+srv���7���_�'t\�ٔ�%;�T��*4�h�҇�t�UϠ�T����I�- ��Q@���RydH$I�����r�J8׼���ievZr֩��
�F�q^ʎ��◵Y�����c������{��۶��3M:�i,��ik�^�TybPc%��� E<�m6���k	������fʌ�ʍ�Cb�sԫ���(�$R�L����V��Z��K�sW��ǰn&��Ʃ�v�a�ѻx�:*��H�/��^�zzysrypF�H���i�Q�N��J�4'
k�!bH-�iS��X?���Y��'.JɊ����s���[��Xh͌��RL��R1�f�TTDX=����,~2�˰���ӕi����l��&���Dh!;bU���q��������XC������|��t|�M��5��O��L�|`!�����I]AV.���twvf� ���:�Vb�Bnb1�Z4�+|��"��x؜�}�����xg��x��������]��Xvp��,p+@s.[�L.��K�BC
�+����n*�B\��>s�;��V���d$�$�ݘ2�8�������R�Ã��-��nl�����A�㖑KS��Xy�f�;�Q���4�|����X��`�!r����si�pQ
0�YO�gOv,92ID�6%���7��� ������`��_�_�\�x������ɮS��2	�g�|F& �ݰOBc�LL,�v5 d8�,�Hj���6P7�*r� %��lҭ���զ+sЍ[7�y�v�J*�J#��UUh7�f�|�tDF��5?� -QG[�ý��A��(����X�Ed��ף�F�C4�1U�8"(8+V��΢%�����yBƘn��U����Lf2c�t�Xߤds[[�د-��}S����lf8��T�z����~.�����ԥ����pu#�L�
7�{l��s�"���$b=8<�"�8���4xB|vm��C��b�\�'�s�6�I�a�D��m�P�7�|�~1J^�8QQ�P,�jJ�4
�sd�B�'X@���l��:��#D� �x5�3e5�BnJ4A8�Ġl8-}G�/�<C�f�Y4͊��a�̪V�˃��H��\"�,�P�:�K:[^�o̓6o�hY�̩3��c�y�l���t�d_���t�ڽ�W�mm/�:pҒ߈uEZ���V�Wp��Oث'�~&W��X���lnXNe��z)���(��(h]B�A�o���w߾9yq��	5�'+�� �W�;6�O��A�w��Ў|��d�ߖ��Ta�qgF"7����<��j��YT�#xo��j46�S�7�$�	~|�c]�
>*����0WMf�!�{r�����������Is�|v�5{q�����?��I��{DF.��ZYY[wm� ��F�II�2�F&�l��7�H��J�z�وz�q$���1�e �VkVn�/���߽�f��<ݯ��{�g?�*3Ntd���K,������>=�d������h����f��mgw>�潊?A���Ep�q}#�o
�ŉ���z\gt�#幋��7d�k�a�]��&"
Z����{?~�����r6�k��@��p��;V00��h5�'<�����9�c!W/��Ɇv�l��^UP����奨��%�>��$F�VG?9K��V�#ex�T��p
�n�f $���o��/H�O)w��{�s�h�$#�0�;�f��m�6v�O�/_���HPR��������ٝ�����'xXey(�!�2e�Nk<NQ(]5B�ND��`ov��<��V��Q:�y�}���yzv�f��P2�n�{x�{�<n��pm�\��b"�4k�+�l�0�_}��O�F�')�A�+.PX�@���|�1�ި�!�El�؞`�Y�L�_;tM	F)����9��Ï���E����֛�+���=��"��d�yo!�QèOX�w�Z�U6[�����{_'B�e�r5���'o���m竛����Ip(<H'8� �!cn4�B�	�r���SbrЩ ,Kqd�L1��X���J��3E�X�v��½��?x���`��\CI3~M��b ������������͋�/?;}y���7�c��|.ē,X�)8e���}+�j�m�݄D�H<?<*�!aCpȃ�DKX*��@azX߭�����rԽ��(�t��w���8���y4]�m���}��Q�כ#�\w)&����|���f-x���M��w����_=��a.��Ӹ�������"0��
C����?z��ÏVyYƣ�B^J\ ����6�⟟�z*���հ'Q5��y{��%u���E3Z
�+�_��Y�k{    IDAT1F�h\�DO!�0,���i�FP@�Nѣr����]B��
8��i����A��}�N�7[�c���7�)��tH|m��὇w�}�/��q�g�$�m���o�k�@$�a��q׫L𬐙�?'�;*�' \΅����W��4�-/L�ݼ$�,���f��������Ǜ;��dl��9#e�@a�IRqaL �c�������W_\}��ӫ�ޜaq��F�A��%�����M�q���S�L<rPۉxI\�pu-3�i�R��d��UD`���PW&�R���ў�Y�8�ڲ���W�����`� �ѹw������m��)+�ɚ�Zn֥�p���(d*b��>/�ǝ�?��FatT��-O\��-��7��G�ɼ�I���7��Z?���;���+�S��K�ߒj�RӨ&vDq1p��W�7o&�ߍ�^����J䇹A�id�,茹�׷d�ǉ)�
�����x�{�<�����"�P������P\]�F�:�����Z��m����v�t^�ƿK�s#�p��{�����]���Y��,����XTb��pd�0D��D UB/Ġ��`�s�\��@�8\�o��ni�O�kP�k�p�ኣl�\��z�Sź(A��j�Vy�^U>�qy���{C��E�Ѳ������ך�ң#(Z��m5(@��F}=~t_���b����9���i5���c=2���M���G�]���v�+iŌI
{�d
[�,r�H����+ޤF!ٌ���1ɔ�y_~��[4\^7�O,���y
�yRl{�m�ӦٳgϸӘ�M�Dp��o��#�Q�O��o6��[�~0�X�+���2i��G7J��9�)p��կ~�+��8����?��GON��x��Bi]nȬ���DG6'�E�з(o�':_N�3��Nt�ğrf����ty�|�E�Z>�)�qH�j\m4(����7ȇ7���ۼ����� ��2_ �i�O�tW�|�=n ��)��E/�rS�.��W������~�@}�E���]�h��B��Bܢ����Zo��P���G����3 �;ax�-r<��c���X��hvU��]�ݩC��ӽ�H{Ƈ}c'	nM JO�4o�08X�~$K��,[d���&�S�H��!���K���gu���_�=�˭WO+o�����§�ܫ¿w�R�HvUL0_��k��6�n6ח�^����ѣvgG���\-@3m��tl�`��f�56
͇Ym\q���u�6���3��i
�B2#>W�y��gg��a��?mc�^���D6�� |d1�����?����/�;'�r����ۯV���IlH�Z�����b�|��׾��lL� � r�S���y���O&�wW�Ӊ͚�n�`��śC�3�by���W��뤼���.�����[N`c��yQq�m�s�8ҟn�B�!5s���{��j@�u��sx.EV�	�U�CJ��!-Ռ���gi�6�`6Y�}cзY$���_S�L�N	�+dB}�����Q���ȅy�`��.{�]B���bA۝���ҧ0������i���2�L������	�cmkw����WC�3��$șH+
.�;���u��yl�~����~n{�B�%�� \����4)%ar����\p�;w�[h�[���}��v�4&���٪�:���ɽ����+I��$�g˞h�py���D7�l������Ո�z{"tSZ=���3�3�6���O"�7���J~�Xګ��x�Դa��G�#��{US.��xd���5�HЀŀo�su\�M۪����fl��*8Úd��٣C0AL�7�E�G���O'�mWdZM��օ=;<�J����A`2pM�D�U��%�H~hY.(�*��u�AP�[�AF:�wŲEhn�4���V��6<�5��T���N���Gӌ��> �]�z�c�˱��m/q��]�:sX��D���DӤ_܇��E3��
{'�9�r����A�W�������b��0WO���:��a`rX �aMo�;6�X�+����۲6���RA��6�>�QGi!������o���i�o�{����w'�օT���BJe:�O8ND�$��s^^t�w1;�цۮ�6N�I���dt�fp�S��6���������]���P��y��o��q$!�kH��!&�0�����U���gg!�D��X�b�L� lg������v��滭q�:�!v�I�BW-uF5�o�Ď0�Œ�O4��aY%�<�/W591���QC�Z̈́�r$�UީKD��|���G�Z��l{���H9�Y�e��<\/�f��G��K��
�G�� �����<:�.���߁yI[J���)�]����Vx�)�@mר)`�dC�;�{���ZOf�6�PS�7�ׇ)�)���y���]/z��2��iw�bF������yD/�	 ��Y���Z��	�wi\"�o
?�n{������6ٽ�}p �#���4�}}�z���Is���V�l*:So�o>4'LJߪ���׿����n�O>|��ϖ�����n�N��W�o)� J�а�7��Z
� �l"��m��u)�q��ʣ�+B{����̑�����߻{��'<��9L����c]MLO��D���}_����Ȫ?{��+����E�D��ƪ��hP�Ċ|3�TVD�4�1o�"��mk���y�tG`�)X�.��mZ��x\�
&'Pc��N����������j�����%O@. �Y�_�s"�3mη''[��Z��c��esH�C�!�U������{�����,r0�E��.�'h�p�y9#ny7��Sn(�6*/<x��u���G;����Æ��m)�TЬ`�e�Ӿ�/޽:})�qF����ƃA�5�	B�������'1}^��t���-���IY�"�l5�nQ�vR}�#�qP�Ry��*L$�s���w���v��T�OCL3�+�f�q�9�J�)��zu�����̖��bw�і��M[�
O4�U����������IZ�K�&��)�
�%��Fm\Y{Y<⺔�@#,�����>�{��\�!0�L�B��,����1�S�,^�����JU����|6aY�)d�[\��ڛBƊ���PD��כ���V��8^�p'"�$��"D���3����ڰuʎ���U*���m5·�nzRlEj�<��bf�Æ�x�5{����f�����|��՗}%FV���0�,v�*Ce\$�*���Լ�m���85
4�m`��@� T��F��Syߦ�=ܵ�y~��O���ˮ�Z7T����
���$�e"�8��.O�^��|g��iVDqx3��Ǜ��ߚ�E)�f�� �p]�ؤ12��rKd��TL�fo�m�ǢE*��8-�N,����l�0���J�k��t�WEۣ�@;ҎTґ��'ѳ�Ѯ>?~t����1��s�.�ђ>�E<KЁa@�-�A(Č �PX�"�.�jy�wN\/錷y\?�ߏќ/���ӟ���q��֭�]2h*�ۈ���H��ҍ��|�\�~g[���5���&�·�4GZ����a1�����Q�>��#s����0�["��5��,�_�7iC7�BT�}N��_9/kl⹀��{�����IqHX�Ί(V�p��`j�� [vǪ76;{�omo<|���ov����Uv�n4��ǧ�R�-�S�<���`R@l]ެ���PV�!C/V]��·�ol?q���Ͽ�Q��c�@�)���A!#�ͦ��>�|�̞�Į�Wv3��_�;���P�R�����$�8�ʚ�MJeԢ�+y+p��Hx��_@Z��v�!uM�-mh`�I�6�,�u��]J�����e���gGLU&vR��b�!@����C�L�\ͽJ��O�w�3����p	�o��'�-�[���m'u��� ,kc.��@���1�9�T^���޴�b2�
a�aN�\�ɤ�t<���t�1��X��|���ýM�L�Ҙ�B�Ss#��3�S��D!+��W���՛������6`5�E��j��gf7�M�w�C��K<�_DiBs�G�fFʟ�¬Eiu���䡚� 6niʦB�PL�`4��Qg~��Z�4���E�L� MН��:�G����7o֝y�����ns� ����}���
����n��MU��[t���k&#FՠJa�,�0�Mqdƌ�s�Zb�9*d1W:~�u�夓��^������S��Zg�0�/�.4#CpS��*QM��ӗ_��~u���fg�r��wY?8�J�r�D��@��=qx $�B�~������!ͅ���X�d�$t���S@H���j�k]^�!ۻ3�!w.D����2��O]�mv���6������o�t�.�bQ��Gت[�%��!��n~w%������?�Wڔ�K�i7�b��F�D�����P,���N�������R$_�,��Ѕ���
�?H>�w5���6Ԛ�_��	 1[v<����)oJ�o��ܩ�L1%b�_�䱃@���
%iķ;m��H#�S�8�O�&�k�u��2�A1������������kU�X��:k%"��)�󦆌�iۨ>|�z�����E����B4��Z��������.�0��8�CK�u����C���f��Q�	ֆ��اy�~��û�e�{*�M�o�Ij���J�$f<%zfF�;������������&�F�GE�M��-5l�r�.㹵�{'�$4S!����%sE��5��
c ��}]����x�"��1���zM�p}|����IMr��Zz���̰���
я�r���_"%6�;'�����F�qmj����L��~A�X�,��_૨�$�+Ԛ�\
:�_�^���s�c^H���x�B�"�O�����'��{?����ǂ�GWgt+�x���<bfb����-ڨ�8}5|�v��o�6����X�U\mu�pr2�Xvx@�)����  g�/�� 4��y�Lm#�GM�J�G0E�w�2uj��{w͓�+�AM�8V�D9qN���}��h�yurv���U���p��jo�a�8dR4�VQ�%<�$���D?���2��D� ǹC3o��%�:��Ew�x��SK���u��V������~E�pPW������+���{�/o�u��"�D��	L�,�70�Vz�t�����Ug��W_��so/�]����/^\��Pq>����~�)"��9�NB�����Fg��
z�|g8�Zp��!���s>ޖҬ���տjih����.r�����U/^��)�ފn�zj�)cDU��]~P�v����̫J� @�]���F<���?��ϼ�����M�Ө�������{�;m�=q���zΕ���)߉71�Y����qX�������(����U^��r�xЭ �t8/wb���8P6��.��w1G3 @� ~�^�f�����Ӕ�ƥ����뜣�ɓ'�n��\��K����6��m��["��X�N8d��������_�%��?��)�Q�_|�?3�{��z�s}�ҹ�:�s�������b0��A3ŒD��@�(�@�D+r���P�����U�QVV�h�4B�`��L�T�n14�.��>�}�DqXM�A<1'��A�zcl�+�y�Σ���qK�����َ����޻�������f���j{s�M��-����`���{s@I��Tw�N������}0��n�.�s3I�Fh�ާү��;�v���@az ��)�V
���"�'��_@ٲ�D�9ש�ސ�é�����+
�r2��b:��F�fuxy][l|�Ï��_�ѓ�)�@D�J5���{qm�G�ݴM�E�ֈ��-1Ub�/t�E�J<h�յ���� ��5t�
����i���p9��E'ȋ���;<�q�	��~��G:��_�T4O��D3�w�#e?������-O �l������f����������ڃ�hC��Jǘ�
.�5?bb\b������;���N�����eb�eb�+�b�R�:�����ΣcV�RX�D�����	6�nm�t6+�潱�kU�m@���Ѷ�J/�������|[i�H;��`xќ�&����B��V#j��R2e%�FBd�����{x��B��r&���Byi# V¿��r�%�1}|?n!�ڻ(��ǈ�鬋���Nu�%�G���v���{����i����@Xi���11�D�*g_��d֟�g����?���<��t�m�?���nNu�� � �@����|9IC]�t��XtS[�Ek���fʬ��z��2o
���2L���Ge���p:q���N���d�+:��K�����h�	 ���e�qy�y���G��W/ή�I�/��;6��Y�&��K�L¥,�V�-�~���EH�p"W :W��d���Ey�D�����ns�U����2fbi��H�P�b g�1�b�|�v��_ΆtRʒ�E��ڦ��O|�c��pqS.	��_�a2!�D�����Q�,y����`2~���d86XB*�������_��2�f\B�H�l(�YÁz���a�Iq�N��5�RA?$#�8ÁE���k���ޭ5����?�ս��u��*mj�$ࠂO��c��=BP�A����L�e!6�\"���)�?*����r"�o�Z'����G�����ϟ<>� �'ScJ������Y���٬����we��yo�0�63d5�BSJ� +�ޡ��f���ߎ��N�a��+&u�Fl���x�����$���z6g���b"�A ���L�˳�C�t�ӆر�<.ƍ�Ɍ��NFW�=���踱����0}g��U�>jH�ΛB�R��O�;��`b��i6�(U:�*��W�1(Y�iAR�B	|��])	���̃���G?��ݬ��W��9"5$C풑�faQ��-wm��^�˯�^^-/�We܃v�^%Qd��Q��X� <_M��ՄHo�a���,�D��7&u�J=Y��K*�-KMR2)Wy�&��m��dT�l>�r�lx�v����Vu�9m�6<�{Z=���7U)�9�2�KP�����/?��?���}�K1:S�TD=���AY)P�9���<��<)��;@��G\�6��R�s�X�����t��Y��)ŏ���	�@��k����Y1��T+�2yw���L�幝�h�{���5����3ME�j���۩Q�cAF
�ĎY(a�v(���w�O��u{-o��DPP��XM��4�:ol_�y�h�`KGf/�#���'��X���JKm<ٿ��ݗ�3^�]ŲX3T�`Zi���D�,� ��d�Iy�y�V-�!�m}�e�sK��{(H��`2�+��ǟ~xb�a�8�r#���:>�J��Y��'�f�U���S[���c��F�c�$�c`ƽ7�=�QAk��]*p�*Pt��|��P���pKM����l]�&H����vaW2�� �=<����Z������Vv����V��h[0P�w��!���@�e��(ܹ�����G?�?6�CW%����~⡩5� �F2�X�a�3�? �F�3����@M�+�S]��-־'-R�n�����?z��U�P��/��ly1�B:��Uұ��N.g���<�ϯDvU�w�F��Db ���K�XlV�Y��f{;�����4�4�^8�
�G彬��]��Zb��8�?`���i����NO;j���vn��~S�g#}��bݠlŰϞX���q}�����Vլ�hO0��A_hf�W������a~W�5¹n
2Ԕ֊�Q�'4
�������|3�l�y���x��ѝ�G��0�ȚT�)�62"�Eʍ4$��)k>��G�����|4S[�AM�a��F���Ͳ���t8�5#E���+����'��ء
%EU�
�����uX���'�F�#P���Vhm���wmEXyF�Ӧd�fc��j%%%�$P.�}�rB��3�n��z��޽7g;WyjR�Do�v-�1�,H\��P��2Z��`h0/k��ΉfY�a�l��	Y%o�q<t� dt�����w����G���P�l���C�;Q3�����z    IDAT�Lf˯ߌ�fv�&F��ƾj�ͩ� ��`2-����J�$�8������pT�����"N�� �-	��~��`E��rEP��w�e[����P]W�7FG�+C�R�lk`�b�5��e�[ǋ�7�N�vd�\@}�����ĺ��j�Ga���t� �$4Af0�J�bȓ��)����?��6m�]�eƺ��<�?�nlĩI|�P��Y�vsP!#��F�1>Ex�cp��xy6o\UY"^���N03�E�C��Y��@�C]�5,����J�7�BrL��R0�����o8^�|s�zJ<��X)���"lNF����������B�ƨ%�����z��厊b=�/�*��+��[���W�Nk�ד���b�w;ީnT��&�}�s��� X���v��cSf�����	�fK�[��	h����|)�C��_M�c4�Fņ��es�����V�g�`%��Ǎ���t|ʣ����Ӷ�V;gpu����/����SW+
��snW�^(?`����4�p3O��f��OM�k�U�(��=*01/p9	�#�C�;g	EN���H�{�t�����Y�ޝ��Ym���r�����{#���f������x��?�Tqzڛ�<-bYQ
)���Ff��#rF�*f�2��u����[R�S��%g��MAO(�A~+�V��O{Wg[[ݛ���g�&���VF���1b+#6'���җ�׳�ị_����{Br,���)m͠��N�(n�.A6I��ȃvoi�R"Q��4n�D�$���0TN���5]��i�c�L�D5e��w.g�g/;]����UZ�"ӓҊjeM�.jj�N�`/�n�`�����F���zC�����\�����m4(��"�����9LQ�[�/$��H�ț]l1�aм}�����ꛍwW�i��M�H!�@F MAM���_����+Q�;�A[� �ӻ�Cզ��]���>�e�yI���gM\ͺ�V�v'U�7o���R�.���\l�/��>EL��w�5������E}��VD,N�\�N�q�<B��x8�6l?\;x�����^��J� ���G�5H|��F�J($�k�.���p�?��~�3�8﷔����73���A%|h���O���ǩ�3ʒ,b2���c�Sl��� ��ԕr&秗�u5*&2�z@�-F�FR� ����lx��.E�,f���UJR<"�cI�𵱱����0k�nʂ�k��P��՗�s�t�V�����@�4kAĚ6=)aQ�ҙ�U�%�9A�~���'��ˋwWo��]@�x/��I�j�	��5���oR\9�HL��P��z�%`�k�if���:���DH 0^{���t���=x��C����l>�i
�,�Lh0%�5lL�jȱ��o_���򫷗��x��#� C6�|	E ���Ӷw[M>-E��2Py��3ڠ�:�V9<�'��T�^�*,��/�(hi���`�{	�T}���a`���D�E*�s���{�׽����?8k\�Uۋ�j����{B�|��O4����DWq�gI��=
��`��|��wL6@)DDOi�OG�L\/��Sν�-Wʗ��f�y�P�㮏��؟|�`�=�],{��z֟��vM�MhT̞D�ƸO�_�SLy��u���߫�����/�<-�s;{TU�,ꝣn��Q��۷o-��uS����|�
)��m/Y�^�z����F�b�.tm�Й�O���5���f�}fO�l�	�50d�]��=���Ç���|1(�λ�18k���>�Z�(�h��tˡW%�|�+��T�)}���R��3��;nw?����#�׶�ޒ�4��lg������F��n�]1�ğ̵O�UΔ�����š�+�jS6+���p��'�lh~�g-���p���r��@<���h�
��?AɃ���6һf�cUzU�HyL�o �h�O*�]v�E�J�6���ʴy����־�o�Ϳ�L.����rV���K����� >N����y��d.�wj��`�������<�,_��P?��6M�(v��C.���ݮ�}k���z,>F�h#�%E�}�B(G��E@s�m���A�$��� g�oaa��nmwxN.���ޡ��!	��}Py���������բ7>�Z���[}�Baw��R!����Q�ٺ7�/��^m],챞�:�����S�x������\�L�H U:��P ĉ�L�-�2�~5vˉ�49L��E�O耂��#�T{��j����*��U�]���y�������o��d�A�����b���>�s���0T�!��0��f�
-&��DmFwM��Zx�_��Ԥ"��P{��=���?UG�X��ٜC,̡��c^[^�B��5��4�k_^�Ѳ�G<��Yw�[.B3���[ε.��Ox��2��UN<���G���-� N~��O��6�F���kh���$���2����O4�׿x;�vh�H�P$9C�1��6��F@ϗqi�a�� Ԭ���x�N���jg/�nvt��	�,=��i���S˝����	��G��C�ʗ�F��*/m���m�����E��'fw�c����`s�����֮�f#c�%��e��$1d"
&��t �s����������>WJ�p�-��eI�vd*����w�s��oA�V�h|QPV��������� ɣr�`�r�S>�w��V��������'�E2۫'�p0��X���)O�I�&���+EK�M�͎n7�"�9��qr<�1>���2q���E���T���mE�lo�mwf��������,��Y��}�Y�B_W:j�Zۋ�N�q�Yow�5!aʘ�ׂ�@x�0T�N�I^�3���
%�5bb��:|&��/(G,2�{$׆���H���{��ho1}�E���y
"��0�eE3�f��T�sE5&�'ܝ`'�T�(�|-��,Cv"�3�������l+��+�\��R���W@��8?��gbogI"����Y���Ԯ��]۲��S�F h�}<�Nb/��6'�EGf-wV�B�$+�کՒ�������پ�{����W_�~ym���ņ��ꐂ�c�"��G�?�.(��_�$ ��x�s�j�[AЂ�8��}�Kc��ӏ����O=}���˹]�Z�-.ź qGvq#-縠���~�<�x����=������x��Z�� �q�Y5*i	�7�4��,�SOV�u#w��IEd�=N%F��t�c<u�6��_��0v5�_^�m�ɪR�H8DH��[J���RSd��p#�E ��b7�/wN޿���dT_a#JSȈ���X�s־Џ�In����I΅ɴ;02N�k!�0C3#b�Ke*��Pad~�������x9�9:�:�5���_=���Wɚ<}9�^$�����ͤ�g3d�x��@g�LL�>�w|���~;�^�I0�0����Cр��r��:$P��Lg�(�J�m��,?�Rܨ���Mwonk�]3��E�2�'�)*0EWh=�!�������7��_]N�n�v)�ݒ,*��Jt="szz�U�
S>�KKr�u�' 䊵�Y���D�S�7.p���O�*�t���:A�Cz�߱ ��3"�2�8왭X����ͦ���a
��}��0R�䧡��⥸��Y�Eer�J��4��-e�`B�+Œ�P�P-+�`>���ʓ>Bх�l�#�{1{w�Yow��Ч�Z25(ؕH
����g8�&���{�8����J�=1!�N��*Q^V˪�s8��� O ș�����R4.�������2��s�kdU�Ń'�=�ݪLm���.6��" v���B��	Ԝ���i�zu1��`E�| ۔��M:$�#�|�H�p}K�S|�mX���DV悻�ND�l�����5Im���G����������u��F���r��yg�Ug]4�8'h�H�crAi��$ģ�Ut}'$��?�]|y�S~xA�u���a�#c5K�J	��\[���>]����b"\$�8�� mP�°MT"K3�D�gO��9hm��V�!
�f_^��cXG1��U	q,�o^K�~}5����r&�����Wv�����,��TW#,SpnX��ʆ�����]�g;�o4Iʍ-�<b��qy��l�mX�0s~��T��ེꜳ�ק{�ݝ�n�1tC
c�Z��k��T��x�/)sk�ٓO~�����'{�.����'�]G���(���*�
�܎�lĭ����xɯ1�@�TQH�!��a���Ȉ[^-N��ӧ�K�i6H�)	��GV&4)_ �P��C�����_�` ���o���O�Ց�S�ٜZxk&�Aؠ�� p:�S�-4/�^5�K�Ļ2���=�&Jk������g�(2��R�����4�s����q�b�Z5q���]l�-��<.p(

xw$�j��{�p�yi��qj�
�I���� �ެ'��N�c�(R�1���zZ�u�SQ!����BY�C�0����§R/B�~��O�;������ޖx��Q�jRc��c�I��5��xu�ŻI��q*a�(0���%n����`6c�-A����8��w��o'�]욜�l���2^m��$J���Ck9�t.a7��eotq�zp�Y�}��k�?Y-�=l�MR![�5�[`�����'?��|��WK��=ȽW6�R��
�oH�5r3OE����
̮<���x��yxM�{�;j-�Z��r1!L 
�tv�t�'��1%AaDx˞|L�B�4;Rz�<�^C�������ߜ�z,M^�@��!mc�~%���	p��ѨM�͆�v!����r:�b�=�wpH���~�gY�BuC&e���xM5�jl�*P;����b�%r�i���ʉLe�U:\U�x������_o�۟)�]lu�����X��R���&x�2S���ld-<��<_���&<O��n��y��Pp( ۳�?+����N���y�?��'�GN4�h�6լ"1ylGn\ͧ�q��l�W��w}a3A�\�G���U���b8.K��9�?J��������A�߳�dKpQb!b�.w��9)�7�#��*jg����s�Fc7�|ŊI�Uߝ���w����e�-y?���L�`��EJ.U��d�ѣn���X�z�z=Tl�9g	i1�*�K1��$C0J"a�e���%/f��9 � ���.�AaB�#b}�}Ŋ����'�Z7��d�U��"��z��;j�� "��3�xy�իKDJ�%�NV �D�Oo�(9HADmq	H�����7n_HbK���C"�py���L�>�@ �H&ډ��x!;#��$N���9?����4PR���'�K�7Rv���E��+���n?y��ߌnN�/�Z�$�8�"<뛧������8J��'ni����w��å�.�9 4�B�A�I$x����ޟ��Ի��Uu��&������A��L2$	f�g�����7���r,��v�$Img����n���+e��H���8�:%
n����h�[(�tk�V�	^�c:�A��s��V�o�{�E��@��U��&N��틫���;��d<Wg)!���6�p�l����t"!��<����ӻ��*\��ʞ��1�" ;�h	��Ԇ�����s�^Bz�M]���X�S��(jآ��ـh��?��-�f6"  ��:J����+rfb��ʀC�Io��ݬǄ7������ѭ��L+Ku)����5n^�y���h^�R���D#��F��q��&� 4�`�^�l56�[�z+r�͑&ק�&M��(%���̖M�H���v-��#8c����ם?����/��Q������H*83��_�l�@&�g�&@.$�H)$щ���R���S�X�����,0[;�`V�������ѳ����A�L�,;X!Ԡ��,�����E4'W�������w�%�c��aTuiK�,�D�'�0�� �����!3^�z�ZQ-�%��r!eC�eG3���ّ�O�`)��_]�G�������a�T%���*�ȌKu�F(V�ƕ�����������<?��w���lq�����p��o���@K� �iK�6���_��C��N��]������K�ʋ��:�ҭ�Aov�T�ӹ_u�Q§�U�I�	�E�~�Z^q�L���O[D�J��e�a=[TL�b�S����N[b��n��fm\߾���7��ZC���E�R������l>�����*ȉ�V����߽|��_t�_�E|����+�,#"+by����z�u�e2p����!�8�dM,�ܚ����n1Q����E���2>�и��8)�5�h+;������-�`������m�r�u��{�bC���B���bÙ�xӄ vb�#5�0W����}c����_��^�+F����ž�:ZΚ?5�G�;w˹_G����x]��;��������'�0��F :��,�����J��W�={�9m��
d\�g�}ԧ���?����=��>���s��kj���u�Wh Q԰�m/����`��c��k5�>U;�%;A�#�,Qg��B�g��)��x-�|Һ��^_S?-/f�M�;A��[�OLY�)|a��>��4��0C)E��L+�?�f4�)C�gR������s�F6m[xV\����������~���o7o�%�rJ=:��Wj�`��!��Νc�o��˳��h��=�4��ε�{b��i�8(�R8���O� ���m,8��)t �έA$��P�8a@���#�h�Oꫂb���ݶ��������J��9��O��?�?�T�s ��o�痃�W�!RѨ��r����6��3Ӂ�\��uz�=�I�)uG�cG��밵��XL���p8 �3ʿ8�MV�����!3�r�x�+\)��9�p���\c�rݧ����u� A���uW�[y^~�|Ї�������s�f(]|=+�
�;L��Z
9�$�k%���$�'ܦ� ��h!w|�38�"���u��lj�%$<β�w��\{��d1�������nl��٦����!�
L� Gu��7��8<:�I$bܝ�x��`>%�z���"��ֳ������q{�s���~����(�ocn-'f�8X���;'��_���l���VSZ+%`�	 |7NJ�j��f��&�s��ֿY�QE�e7כkySA�i{�|Op��r4,x�(=�C��� ���;띞����F8q����n����9��&�߶:T��m�B0��+6)t��Bu���_yL8"�n��i�ی&�-C���aGe_���ƪ��l4��M��ZwL�gsݩHV�TKnV�1&���UC52��-(�jt;w�
C'm��>�k��F�M���A�訁�&�/���B��-�].
��"�.�&���?�[��mw�?�+�<I	f"K��C{);G�9N�'�ո'�m4\L�R&�^^���m�eS�)�o��hQ�g�@��Vw���L�Z��cl�C�o�/�:�@to���Mx�ͯ�R:�6�l�E��;]r1��k?exX͆W[�����u۪����'D&�d���F�����Zϫ�Hn@�DVv��;��dz40�7�Զ����aF�����ނ�(3J�Ŗ��]C�����3AD�F���G}�O�u;�X���ど!h�ł	���w��`�%�)�iI��H}���)+��1��7�n�(��.��ڬ��1+p�i�D�|�ZeZY�ꐱq|b�M�ʈ�`u��	�}b����M�bPS���p��6�W�{�eA����w;��事b���'/!˒I���U�ͽ������O�������n���=[�[�����h*�Ig�f	���0�i�l�Oܿ��#�\���nƈ�	q�>�%�BX\15�9�
�DQ1�L"K�^wW�Y��fK*���&L�de���y��[���_�Tdv�zSj���b�[�z�[��]%�|����nw���4���WC�v%����M��l�@غG�GΘ��� �d�q���-P3K>��ʦWFR�39��]\�҉�E����/���L��AP���u��l�Nc�&>�l���ՠF�N2S��چ��W� ��    IDATGvl� 0�l��`�#]�� j��[�c�.:���+O�?��!��%4�J)�p�
'1�0xB���4	r8�Qbc �PK^��?�d�Z�\�#���Z!Gp�iD��!�8�i�X�A�P�����I�Ȧ;;��µ�۰L��N��������G��B���)�(w�*V"g�V�!�����Ǐ�v�@��rcڢ�l)�&'Q\����	��u��r�����R��m�k�=pD�P[I��Z{����?<�Y+�ô�R�LjFY=�"��0ɀ��F�itx�����D�9ĽQ<��i��<o�(ȗ����'TW�l��Άf�D�U�V6۶�n5�̼L��D��z.h���o��#�ߌ�Z1������&b^��~��4oo��+����9zY�9��r��\H��M�b�=z���_Vo^N5�o"g	�#8	ۯ�5�YjC$4� ��s�a<��`��`��Ȉ_ʭ?]��c@I1a�Qe{3rpؽ�hFY�uӕ1�#X ��� X� S�R�����}v�+6.������>\��3�Y<��Jm��M��������Hb D�V�R\\��!d�J��!"g� �f�"���[bQƓ!w�`4ޟ*���Z��#��Q�.��?�H%!�7���rgow���F����C��L&R0S�V�K��b'2�N�vC��2Cj���o�M��#N�f�+���CrR=Vx�0�;�{������zC!��b��8��A@Q����ͺ�Y0�]�c��� ҃M2j6&s��ړ"�q{�Nk0�c1o6�[�L-|�/�W��P����in����޾���J�xgAϥz�1�QX{wvg�)��F�BM�ڨ�%��#��(�$�F�Ak�Ew�f��ĸٲ�|�M0�I���~K�t�bA�C:J�f�]RJEމ��7������.�s\������"��Pv���z갩 ���R�@@r���/�'����t^p-�T��6�,���e��e5�-����q��D�UhYn1ƎM[#��<!�)���wN`�����tP"�q��#�^��c��|i&|��9H&r`H�E�/&f��+���l����Sٹ��B�R�(�,]�OZ*}��mh``Q�֯V'L3<��dS���!��wc�a��lTt<����<xx���T���2��5n��"�f�[�(&�}y���xsu���oT�%�X�h:��y�v���]������v�.C�h�H| ��Xt*���Z�
	�3X�5n��րUL��9��^����<9:���d6��W�/,�:@ƶ�`,5�8PQ�"E#�hUs�=k5WUu�d����x<�'61�%I��r��[���.z{A�]��FD��S�u�+E��R��E Q�ޝ_�~w6��4���k>��~�b"J�%@y�j��<����b�dC��o^��{��� ���k�ڸh5<�@��������N�<�E�	A(Ut�H�t�A&���XN�}��Ƴ�5K:�'@go�IwIrD�Xt�?J�A�� �NI>����[Y� ��r ��]]oA7�<���iou5��'>�-GO���\ffKO"���Ra��SՍ�ޢ	 >b��N%�%��y�+��L�J�V����������>}���w�\! )V����E���S�/��/ģ��n'���o�����ƌ�K�G�5�7�-^Y(�	J�,g�"�T"����e6�4B,��X�bc�_�Sv�:A�`�P�$��Ӛ�d'Ic�CE� |��?ct�X�����;��dC���|��3��nww�?y��B�H(�>v�H��0�>iq��:/(�7�W])/��&�49�C�
_��
3چ<h��B�0�Ȕx�����'�s�9Q����IZ�)'���@�L�I������b�Mlj�(��
;�.����'1Y\��m����aEHb;_�ў�	��du�}#J9H!؜l���F&%�	2���MpM�m��Sm����B��AJUrKv���胟���ÿ���/&��{3j���:E:@3E�]!˅~`�ѩc�P�2����C���fDO4�ۮ�^ 9'JD,���.��1D��~������Bj$K�ZO��Bܨ>X�yxҦ��h���j�+i�PA�C���mu�*D>�/�"1,��y��dR�βBU�w�V�p`$�5��e�"0!�l3hHD7((�Ս�����]�{�W{U�����i߼�n�t�DDi �i��n�}�����X��H}NK\ �%c��N� ���4iH��i��ZV74 {�nReԕL�l�`Q���a��d�����i�ݼ8��M8*�^���#
��$֑������>��0%�@Δ�ɦ �/�DȱѨo޿s�����x�4����0�����i �|}{�6����wyR3.�a�%Fc��k�y�f�Ǧ�=H� ��/���9aCp�`�720v��{���KU����[�xVHRX�! bX"0ЁZ������~w�|��'�{�	0:/�zܡ�_Ϻ�ĭ���y&�8<�_-]/�'�'<^��	'ne��]q߽&x	��'�O��� ��)�7��1�Xn7���zG�ݥI���ߨoԟ��^TF1Ɛn�7���)�����=��{�><��$���z�������������G�S�2�-=T?ֈL:�h ��q���٦����a�3�W�^i��,5܄���IK^�d�-c/M�>�G�+�_�v����U��9��������6o�N�Ғƃ��V��I��#��w; E��OV��dݐ�	d��*�+�t��'K�zn��>׽��t�� 3Rv��rN��x˙uˉ�%@�k��%@���S.z�?�˝x�fny��W7
 �������,�C4�!pp�1�{��:/_ �vrr�Y�YӪ=��b' ����ϩ:�g�gO�>-_���׺��:mM������u�p�~��	����ųg�t��̟��]׭rTZ:\,�(��7;�E�`iɏ�
]ȝ��$����Υm�[�Ґ:1?�%�Zo+q��0Q������,�� �Ќ��[� �n$�(�[HO�z�_����T�Ɲ�������ثTX�����ԇ�׃���7�켓G�~�F\���Jw�ٻ�_x��u�����7�٠v�j�v���<�,ub���&������ �g&�L	`ʹy��40�z��]vEc�,�728���s��f�9���Cy$�Js�ֹ{�il٣�렵�������?���h�A���7�W/��W�{v�0*�\@T�Pf�D,�3#B�2�u#l�R	+FT�=������c���I��fW㉜��W���/j����K�(�5XG�U\t�.�(�	�l�����-�u����Y���]t��ρ�f� �����N�wj�p�,�O����c�r��S��'������.Fa4Dn�P
�vC�Ne{aGh\�GeCK�K��r)`1L���Cݭi*�,%�R��L?ySJ�uS�p��!�ӮĲcŊ(d":L��N
���5�PQ��gH����ƈ�ۃ�� 3�|�����=�$�k���a����H6����H�T���fb�)�Id�u�`��w�[��Q����xG|� v3��{����Ï�mF��m̴��>�}�3`oZ�	��y���M�jf�&�v"�:X	P�+I-g.VH�/<�g�V�5
X6Z��m˂�6�͝w�D��)�t (R�6M��IC�T�����nw�ngk=���ג1F�~*��*�ݻ��=�J�C��3zRk�;b���>1�������u�h_6'����;�O��ݺ�ɨ�����q�3LD���Oo��*�U��:^�~E}
j���J�E��Z6�aje�lt��?8<�n,Ʊ�����|(-@�A9~b�aH��T�Keh��U����W$Kl�#ͤ�#�1�e[�: ø0XǦ���^W��v��J��N�����n�ø;9'�ֆ�� �ͽ��EHh���?��^��UI�:U��B}z�{�6�1�i%oо1ȍ����&�u�/��X�ʴ;�������N���V#��	���$���j�[X��(��X�߀	(T&��C�-����ɘ�\����������uZဝjz%�!��d���$�;Xax��HJ��ҪL��z<�\�R󒩻�V�M2��E�g�F��6�b��)*Y�6٪�Pee�©�L������RZ�G��y�<$�����w��J;R�T,�-�I�ao��0E�C�=C��!	C�ba8d�AI��t�ew]�%^��x�����ۯ�*7o���Ѡu8i��G.mL��#ǚ���m5Z[�+�Ӛ�[L���)0;N���|	m�\q��	�Σ��w�fL�P�[wX�]%�ؑc��,+g�k��c1��P�@V�u!��f��k�����m��'/߾]ɡX���4�-�H9=ۛ|	�-G�vQ]����zF�g�:���M34��tJh1�f����<�K�>�h5)0�d����[��l�ƥ��(���瓭�|oY��ݯ��n���Z�M�#��hҔ�$���&�� �@�(0�`���P��Al��[���?Q_������?���a�>�T:X�5V����#�.�C؃�"푾���C��]�T4�'l�@V+=�۞d��C,ܣ����{�0�;�\�"&�؋��|��E�|�{Ifl��b��6K��=U�x#9_T�`t5(ѡ�j�O!�zA�L3�F�.[V�����6ܞ�u��fRu*6�r�T�B،+���`_���K0�a)���ν�#)��+�RFW�4�"d�kyx|���LC���|S�Tk�͖O� ɮ��e���7�B��K�B;���m�$B����oߝb(���dj�v��2f�JOL$�E�۔C�:����jӁl�\���=����Ƣ�$k5�Ϝ	�]�}p�R�W�2l�U����m^V�P)���� �W�A�n��vU�Σ��������q��K!f�����mD۟���LXx��x�����p�K��
����?��Cϟ�������Vs�I`���|�G��������T��p��{�����b����X= l�bणF���&U`=amh+'�\!)��nw�ǻ��SD��oL�k�_a����u�����(X��9)_@�Q��d��tv�9k���֊O(����1Ӳ�,��aυ���%qyЬ�g��d���S�`
w�p� P ���mJ���b�yw2��V@�`pI������@� v��ޝ����9=���
����"za�� \�P�m���լ7]�l�gWݹ}/נ8����O�u�|! @�.!�^,Hj6�bF�?`�"�M�Q֏�O������nlv�
��\�_����s��1��~T�V5t�W}Stn0\�Idv̗	'S�������kql�dYV)��ѕ/�`V�D�h�Q�JfW�AFQ��L����6���8/�u���C[L�+V+�
�t*X��������]�GS����Z���k;�e�W����~}:��f'�,��)���P-j=��7$#J��H��y�Ma̽s�l�Agj҉���3�"��A.~[H�����I�^C,��/�@�04��φ�����o���#]O;���)�!�"u�4
ʻ���ԟ�(�㽓���Ż�K5-�B�,,q��I+�� �"?  ��)p�{��`Ia��K�E��G��ng�nյg�z��kE��<��w���-��`�o9��DFYT^�I�����()���Żw�$�Mf6[ZD����h�?�T��D5!1c3h�G٘
]�b�L(�:��R�4d�"���A�j�҈��V�PBZ�(Y�d�8P� ���?}�Js��ح<~�Ȋ�{"��Pf}.��bHV�r/�j�}�|v��7W ��@��j^^��:�O`Ѓ����a����",5R��J̪o�v�w�!�h��#�!�]�IjgIFc3�١���佣�;ۂ>��kq�׈fAó�wQ��);_�`:ܜ)��2�"�!s1.�n��>�U) ����fk���@�A8�P�L�J�S�I�k�H���& KGڝ�z\��W��#�@���6.4�~�I��}�f$6V�П2�� 1��eA?����n�󪕦b�{u5i�Cg��uL��K#[u�X����v��%����:�?�s�B��(�����x�sC����X�{���ΓG��tH�N$��߇��$0��|�"&U�_-2_��:1B�C�����M&ʰ�4�����Ҟ,aDс�li���!���(	��#���LbMY`dc��	!A�;�mf.��O�������ި-5�N��:��nt[�_>��w�E��$�&Ї]G'K`��;@ �:�*��[`i �iY;��\DI�Rl��*�s4����Zm���~��.�׫EP�N��9P\O�w3����O�Z���ɫ�=2B"���|^�%���X��+�"���T&'#3(~V9Y_W�I��
�3h(j�����S��R��@��/!��d���s;���YR���ҼF-��/�. ���L����~�9�Zq*g�Z&�Ԥ�\��C�Pa�,�%�:x~�d���\/�ŧ���(�8	NYlWٗx�n*?�ɇݽ-�
ă��&!�YJl�zTÔ�����|kW���۳Q��@Dz�/�8����;�.��7�Lp@����A
�du�.���Y��p�ݡ�g*hL��R�H f٦]�9a��&\����r�4v��-� W�l����lށ]�}f��r>ە~~���ߞ��`��=�����R��P�`(+#7�%�q+����0���i��!~������)C�ɘ���Ӗ*�
��������H�C�&h��!Ez�OC�L�fQ���{q>����c鯌�19L�ԫ�	�,} �n4w����"���W��4�dA���4�qP{�K�cV/��@~�8�?�Ub�5�#�!o*�^����
�a���d�)&y��G���a����X��[��҂��G�����
Z��=��9°G�ß�sGyѯ���E�M�����]� �@0����x�G��ny�<�����B�Ԧ���`��P?�%��^[~�u��_���5F�ˏj��o�D�`z����DW�EbCz���]E�싎[���d��[�O��і*�k�$�J$#mv`��*�`�77���s���īr��}NM�|�0�^`����a&��E� ���?�\��̯_���w��so�B":�(��BJ���O��hP�?��&��ǳ�❌�h�o�@��!t��\y��~�Q�s��k���$b�7�eKa\U'�r�?�!Mh�/D�!��iJ�+����L�?�)'ԉ�2�s���FW5�ƹQk��w�k��*g֯�e���Kc�'e{����$?�����o޼�+W<��Yz=��L�*z�9@҇�uE��Я7��q˟>�i�Կ���Ј����T'tH�ү�<�����ʇ��o���kT5�}���+��@��bل�#�ҧ�Ʊ �ڞ'��AWR��zr��bu}��uS�B<.If��@�I�@�0B�L�>1_E�v��$ |�Of�Q*����_$���l1~�Hwstr��׫4�z���R{2h���?zs���]m�7��xf-$dcUߌ�7:G�?�	���4�P��O�%���t��6aC�.���z�Z�Ц�իWV��)����j[Z�}yq�}��t{�K8 ��QO���lڶu��Fpe��G���j�ָN�[��=��G����}��j��d�j�r���b6��!A_��Z�K����������|}+�E����+(��oyd&Q^sOWP�xa���/��}�,�&�bCrw���b��C��#y�u�U������t�X{����c꾚dˮ��gVVzSY��5}�7��� $�GCMļ�ARz�ЄB�`HA��b����6�߲�MUf�~�s��<@��<u��k���qҟJ����x\¾<v�a{�O�����D<�-���P++"_��J�d˕#t���Zv*�i�r�T"�W*h�(�b�"(
��ʼ    IDAT!1�Zl4I< �0^(v��'&��b��<З�y��C�ԭ�A���
���o��
[��-��I�IGjT�Z��Tü���V�����x�X�<�C5$TC�s���SX9���i�:ӱ6$g��[W���`7$������
,L7��U�'^X��{�1+�%<=Y�����r�|��{�vSl�"?� 20~���ފ����׿x������}�0���93�Az������k���\��Ke�bUR�7�F�楞�&�g���ק��b�o�J�h��C6>,�)�P��s�S��k�r�y��v�o�Y����Z��ܝ��f���7�4eKB]P@ 7e�A2���x� �f8:�jz�����O��8��O�$\*>�H��=zBىГ�V��>�r�恘4�� �YP���]ZQ̎�2%w�����t��L�j�d�[�
�5�K��c��ĳD�D(������G��P���R腭d$v�������o)B	�P߷ۺ���ƨ��R	C?>/������b[�쇺ӪUڽ�ʭ�sw�>Rn�~%�9�&u_��������}U���u�Te����r�R�1E�����c�?UZ�B"W"��p:��IE�#K��{�,��8ۓ���Pݕ��t���TU!�tEm�7w��ѫ���I�| SD�R�\�	A�ɏ�NK����s��%c�p���ec��pjr�td(�/��>��bDv�+�ڛ���Z�`_�MQcc9�j@���K�V�K� \R41�1kc���������L*I�n5,O�5��׷s��P�gԎb�';/���>C�w�[n�O�lv��g,�g7�'me�����ޯv9�L��wj�+��[���p��	���h�YBVg��#�kri��١������_��G�ڭh�hz��Ő������=3:�o�X%�X��1�Z�����jCV�(rz`�f�(Nd�������Z���)���#���߶^`]��W&��(��~X��;�������z=^�ݫ���=i_*���t@��T�mF�N(b�M�0gK}�]LFj=�zÏώw��Hβ�!h��
��[a�J����]���k��k
� bb��H�-��Δ��W�=�t���;�ȫu�S
�4=��)�Q�s��������^�����T����H2�`�b@�Fc�a挢��l����#�;���P���2L\b��������;xv<oQ{V3�>OC�ݡ(0�Ļ��J�˃L �z$��H��q��<��=r����m�''��n^�V�y��$���Kd#z�������BgJ�,�����
��`����ֻYWA�����ˏ�<��3�o{$R�`���c����Hed���7W��]eI�j�t|���6���e�Bkg�*�9@DmH�2{G�9���h�	5��7�D(��o���d[OwTQ��ovy�R�fKO�Lo߼~}�뜜u5%����F�!�L�/׃U��@����~����o�V��ەL[�b?�BLᨏ�дy�L���
�`�*1٨m�3(�8_"���������W��ڟ����gj�)����0J�;�k�O��`�|��v#\�����q���|��FV�:}4�sۀ�y��͊A����i�F��+�Xa����x�M�='�sP;BA�·YڂOnSp&��~,�!a�?�;�~��ZfÀ<�^{2_��:�i6�g8[�3�x�,���6u#P="3�f��������R��T�7r���f����eK����b������R�@E��e�!0�!�h��X��{8�ȁ�[$�g_~~8��#���\U0��&͊�G �i9��m��������_�aC��D��(^�`G�m�Y!{���L��I�1(*�R���kXV7�/E��O�V
#s�?M�0��欬X�eQ*R"�-�Vu���* ���v�.��5v�6��B	ۇ�l�ܜ�9�����/ꛯo����Ր����+�(�tA:�t���|��O u��Iח'3����˼� H�}�h`�˿�Y�[2�E���Ӽ!���ZN��*��g�n������(���r`
��ml�@�Q̚��J/V/#8[S���A���sJ��'L����M�nwDY��X�"*
��Q��bD����勫Z�䤵;�ր8un~I�N��<�[!T�-����<<�������b7�U���Z��*�x6��yʣ��,�	� {yx$B�����c����Ӌ�#���E��o޼����h"���'�?:�k5��R�z��"ӊt}�T�Ƥo����W��\]kѐ ��;P'e2U�?3���K�PD(�U����T=Ǜ��J��bΑT;Y.��&uD����5NU��S��f���-x�a���o�gg�����5�Z5M�A#�x̬t=�5���St�{��<�8�m'��R {����f6:�K#�h2?n
��
^=����[mjŰ��K��p!���L�qK�b!�,�{��ߌgsS6�O�����m�@�/j���BO_I�����R/����lKQ��#r�Zb#���	ߩz�1�}`�T�,������4ګ��A?����Z�z�޺1�Q�ă����`�H���hI�L�����>����C���Ez}�������X\���5.(����f��\����ް�<�ůV����M^�j�!sk%9Lj�J|U\ �9|)i���Ϗ�}/�
g,��.�$&.3
�q(*����~���g_|*.4������h��\]CN�&�����0����񷯮]3���2�$��e�����+!��i�w�|+^�a�hΤ�n6�n_�+�aaWyPRI��T����4�� g9�!�4�M{܇8o��a;�u'�-�������"�d�;�i����=:{zU��no۸�>l���F&ݰ�(^�+���O�4���.(�z�@vt|{ �W�h">ɻ0]���ї�����'_����}:�1�{8L%�Y%8����ņ���^q�k�OT愭04e<�,�%����F�b�^W'G��*R�XD�yS$q.3%��u:����b����������� �Q@vD�Di�n{z��R��?�s�`<83�W���["h�b��<?�/^�$4���UAa"f�Ƃzx\`X�.��Q"kN��7��΀' ���P�¨���Ԍsr�/y�ÏOi��TB���\ƪH���JЖ�ѳ�_]���~�А�{��P���L� ��#)RC��9�V2��{�!�(��CH�޲�Y�y
��D��U�*Ԩ]S;P�+�x���J��3��noׇ�gG0�N��S��VѠl($;�,�aw�tOO?�v��n�����%h����T!�{���pTgx%�
�3?�Å^�_��m�BVAPc'�-	��"4w�ș�?~�쓟}lF7��"颰#S�5�,I�A_C�@�Bk��/x/���c�\��"y3-BĨ:p>vdG�
aM��#���o�uk���gB�Q%�T+�����D�\�=G;VȀj�j�;�O�v$�͚�^�ڏb��2����j���)J���E�*���?���w��.e�Q>��M�^cT�,�	д�(A,�ٗR,�X?L��\�'�;ʅ��G���8�U�r�&��#^z����1YD��_����'��N�t�5�8ﱾ;��3��R'�{V�<�0j�*v�X;�wj��*�Y=����z�u%���t�=yz*Q�����d[1�z������b3}����Y�|��~���|��;�7c �����7���&�����w�I�wY9�����3�2��9&�j����Lа�����>=�������Fj�:�����8��w�}Ǳg���\O�b��?I����C�6lT���4f��d6�[V3U�P9����4&���Q8:���O��d�hCs��`�X>�%v���HA$�,�vrތ|��q�黦\e'���|����2�̽�Î*�����zg�Õθ����|��>N���KOvM�q/}-~IO�7���0º�y�=�˱rq��՜=�;�CFa p�:���vSr�?��,g&�܊/D�l���T��Y����8U�j�5��������c��[Q�@髊�U��w���
��}�ʘn��.�|���h�mTJ�].� T�݄�Z�y�n=�v�?W?�VO�'��v�|t���Ż����e�z\����N�����Ҋ�͗��XfM�)���t)�NQ��Φ?/X�؏Y	f���k2�b�Jl����DH�������Z!�����j==O]����:�۳����pws������֮���D�'�/?��_����ŗ��GH� 9��oW��Lo��.I��^"$�(��u
�z[DbJG�SF��^ѝ�e�"�ݙ�Y-�6�c����Wo�\Gq��q�}�]�K��쨒z�>���~T ᆟp�y�����%���DH_\�/n���k~z���lHkk�^�b$Ɠ]�p��#FH���|�'���#6�Y����"2-��0�u�9Ћc�3C�ڕ�	Z���t/"�q\���]mɦâd�����hb��&&��}*�S3�L�,�'��H]��RXL��X��7-F�T���d;]]�Be��vB�z�)E78�����M��u�V�|/ Ac��Y2��=Za"���N�^�/�Y/��"��.���'�	,ww	y?-�宅��{:�E/%ơ�,U+����O��2�@.v��#-V�'�S���2Q8 ��ր�Dp�e��[�
m��]�l�� ZV��Q��9Y�tA��{����N���Me���H�(q�Ѫ���h��Z�l	;�j����`+a��_����w9n.�ʝ�;8?$�׵�$C1����&�ў�O���I�2ov�����I'5it 3)҉z��韕�����^ �8T4�Y��W���EAo��[��/��(4|�E�8)� ���& )?=�&�Te�~�����>|��k��@ ��eoN��zqHzR�/F+�XR��f,�L(Ĺ>��c�l����OD%� F��D	`�J
��@�񛑊�Mq�2F��K}��mm1�_��[ndv�&��Z���4b���O��v���gN����m�MR}O!?/d��i��C����;��<�[p�2�����Ƚ/>��/��'�5��U!� S]�����ߢ�".5^�>��,:ۺh��SC����L��w�����O^��~xK�y�a�z��({>Z2Χ�Ȧ'|�~?[A�D\:�r�fr=ݪ��c�֗@!�
��R�Z�F�����!�w��o�&p۠�>�!x8���0
�-wc�SV+���E�Mأ��*:���bб���y�!M6�TQR�U��^�����h
�9Դ��n�i��nE�܍߿�ި:�<���0��z虍�t���P�-�'C��ח��ۊ���HKJ�&���}�b\�F���XPq���G���x�F�NXk�R�ن�YS�E�R6�a�O��q�;�aʤ۬f��X�{K(�ެPW��i�^��[<=v]�n	"NM�y����O�j��.�L&ϟ��y�+�Ҡ��k&�7wB�d�{��-R繫yİz�`���aza@Ɠ�-��$�9L>� �i�x`�z�>..�zlB�YXz�� =p{t(��D_�b�Z���4<ޑk�*���%�/9��%��'�7��������&��[&�"
NH�����?�r��`�+�C�SD�Zi$��t2�#�{�5f���� ��$��Y�"&������!;�qΦ��{ݳ���==y2|{�J���uC���_�J��]kvxD����"�|�h��O�˖�A���ǆ[j
v�l$����l�cB�rԵ��٣�//��֌oJ�Zn���%�i����b�-$� 0�*p��Okj����M|f���Q
"fL�f�p��]�x��QoX��̨�w��F�>Nl�=(&*��d<o!OFoW��ŕtd�$X�dG�([��д���$Pdغ��=�l�LҮ4�z#��{��J7�W�j�\������x6�5&�M�Դy;�}�%��f�:��F���߾�3^��4�_��5,d*�i�.�*�Y8�t�(jdq��U���t�=����`k�	�ْ���%����;�&@g))I-0���A�Bb$
�d��4�������TćN[h�G�ǝ�z�� �/H�}�Z��H����ؓ�7z�՟n.�o_,V�9�9�H�A+��nr}D�����ٗ��o�a���ɪ�i�N���_���2$�
�ڬ��T�R>�<5�,k7O��s}5"CQuɨhW��w7�����O��ɇk3u#��Ĕ�c�	)$���ʴ�?���Wx7Q͌[��+4O�X�x��,������"�Z;��%<��,�%��p�#�Z�1�"+���_~���X2�q?�+J ��Pl���[AΟȶ��+ѽD��NjL�G�D:��'���(U��H����IV�{�vH���[

3�@O�P��gө����0	E���vP7��X��F�D|���̽j��]�]���@�xC
!�*f�bo��������p�m\�Ğ㎸�~H���V�[$�'4���RE*�x�q=b��e�a5�<24��wF;M��Z�a����-x2C[M*z�iq��w�"���;���g.�Nd��'������z"HS%%⺅�A�T�y��;���2/���0�9��vr4��6J`<��`���J��
�׻Ӛ��ˡU�Nv|�$���ŵ�����Ǽ_��ouN?����zgW��f��CךT�#4Ŗ`0LY���ɯ�?����\OF�1�{�S���S���ܖ�^��3%1�`��C��OZ!e؃�	M(C�K�U�],_��o��?�Wi�������>hw*}���1���[�()���ma�]BB���M�*^���j�!"a
�TF�Ppt"���0iqw��>��tH��T�F���^H<����p�;,���`ꛙ�����4R܉�����X�%Z���p:��1m7�|ZD/[bA;Qa a57��f��I�j��>{t|��ź~	D�~���q����į����Y-�ee0��Ф����L��금Zv'���+	�rW/߽}��?~󟾚O8�O����ɩ�����øW���+�.����?�j*���lf��)�\�p�η�#���1l7O����e���5��C�e��>;��(|��_}|~zu)�����t��~�g.8�z�������������/�>=�?ņF0p�l�����@k�b&�.:��������n:A��õ���Ǉ�`" QJ����!�!��#�\��ź�?}����ms�?`QI�E˷?89;:��1����E�M���8�����L���Gx��������\�@:����Fm�x���n��K�BMIɫ��y;78g����6�n�	4� ���!Q]�qL����Xi%r��Պ�Z4��k�c+�{��˫�3]G��yyM�� ��(W�1l1��36�z��'����ǯ{?� /Ăxcմ��@z؄�0����d	C_<�D�9�E ��Y���F�S�W �
�z���'Cu�AAXkB�,��0+]�á�w�fkt����͛[jP���z�1F*%��
� �aK��ɞ������3#�oE��s�B"5���?��_�����4[�Ә�լCh�� JD��fD�4�h(�=�j��[ay�ŵ=ȃz-���_FEX}�H�Z�aP�������7�&�يe�i��r,dL	!��yp"��΀	�>K|qG�]�^�#��c��ġ�^O9�_��?��qb"SL���&��ްY����FH�.����$��SYL��;_mb	h@�Hzz|~$u�/������k�S�(�/����$�/�a	R:]��(j��/8�'/Ͳ?Yp�ʤ*�:ӳ~�6*���&� d���*�"�*`�8�qu����Ѥ�~b�[58I�&	�ΰW�����^��4񅆀0�e	�tx�[8|�����E~�F�Q���'(P�    IDATO>}68�zL��k�����#�i�I#8�Az�����w�+\6Ƈ�����Ìp�af�B��P���39���<������h���D���:��e����H��=��Έ�-5��P�1���{�A2��5�O�����I�uD\M��X��	�����#f�s������%�u�՘�r]k�o�jI�N��!��w.�pF���O���	Ɯ��;9j���SId
l�`��u���_2�=�y�8\�.W:���ΐ��u�|�����^팧��[\錟���ATTHt��l��%R�ڇ��p��$]u���kGXsL�+)�h���?=���Ǘ�?��]�+��������l+�qE6�>xrpЕ!���f�1T�ݒ��H3��Ʒ���x%�����GlƬn<2h̀���뫋Ke�'2 lQ"�_���駟�;��e��i*����lD�����Qͫ�K<K�:Ʒ�+�R��N���y�4՝c�i�e��1IS褪%��R	��F��7��(R�jd�U�
���ܚ��<�&�O�bv�R.My�<﻿����9�q�/�I�~z�wYe�=��Kds�f�����@���&n�ݓ��,�[bN�t�[x�]V��a�e��kw��C�p���NMspXK�����N|�<��V�����r��Ŗ�(-�?���Ax��3Օ�3��K9a�믱2��e/wK����Xh�	ϧB�������zy)�������-��"����,���Pӽ�	9��I��"6�	��"�&�Ϣ�ci�b8��Ͷ?Q'c3���N8ftc��x���'������×�/�˫�K�X�\Y�,pdj?
��-n��q�;l��p���#Ll�I瘋k?:;�?��1N)���neC����^* ut��,�����w�sʪZH��DP��v�@K�e*K���DM���x�����O�V�o�{�������}�O�r�|�^o��Kv�F-��+�NW�	������l#Q�/�Y$����������i����@�p�8�r�!cY*�%PPR����_\K� ��r;t�u�L.��n���Pz@�!h���VC)�8�͕>3�b7���O��te��|�'������� 1XaP�ď�lw�'�/^��|)O���0_�T���`�L���FV�����A�`9sd����VK�M��nʖ�]὜<���(��� ��iL�l�T#K�VOMt�bv7Ma�ّF�������;�w[�̍�%%A���A�J���&1,4<4@��(�"���-��㉦�eq�i#�e��L@W�[+,	u&	�A��`:@) ��]H咕�*���t�*�R.����.`�����{�/_�ɽIg���XB��'��$J �Lg���E��� JuS��_�	r	�����������d8;�P�Qi2}�ȋ�j��Ә~T���n���Ƚ�bt�5���t8h�_�Q�{ǩ�n�ɀ�	wb|ٲ��S�m��*\II��:��-m �k��3��a>�8$�N�;>�z��^�?"y���P��H��qkӮ	I�w�,�Mp�e���xN%�/2z%��O&��0UBka�@i���me�J�����Z�~~����~<�F�`Ze��H{܉����)J7O�,�M���\v��*�sq�շ7rz-:-3z9�V`d]VK�]E��#����i�l=h�^\N�Vw��Q���t���t�F���&*����,�n�Ͷ�EfT?j�^3)i�)�t��� �Y�/J��^�z��ʛj�f�
��l�]�'�ֶ>�VU�+ f!H���	hR�4�������d`Q�J�ir���f�}Yh@�H����v|a	H#�D�]��!��@~���D�v�I��W�F�d/�D�y�Z��V4uXr*�L�;P���U��ӫi�7�I�`ǩ2}�tXW|�V͗����(pΰ�J������Fc��u����b�/�8������n:\P��ԔtoC��`D�$'� \��&��k�f�ǎ8L���ْ4!D#Bt)��%8U==}�������G^w ������g;������8���bvg��m<h$K�U��X88
�I��Qaswsq���ܶ
���"�a��\�V�/�}Ҫ��~��@6Jۖ���$B9�!�8$������r@#��#yf�X��?�z��E�m���Q�w=Suʧ�$}�.NCY�vs��G��E+V���GĄ|�T	�4-K�����z�r��ǫW�ԯps��0D�Pd�	���H|�a�0)���!&?�|w  �{]y�_�&��G��N���Z���ϑo�Rz��-!��&`�i���dq����Z-S����F�I�2qB08���'����hæ�d!�.|6|�M��P�΄���h	�?<�;�����Y�1�t�fċ��[��)w.��J
a�V�论�oL��G~)|��E�d]��Oh
RN��w�����i4��v;���&bk+��\�Q�N�d�p��HV�R|i&R�Sg�+Y�����E�tYL�R�lN�V���>8>hLٗ�3�5��%���� �(\�H��aU�O��E)
HT���태]�7MDJs�E���r�6۔.�Yݤ�3Y0I�0E�1�ᑪ��8�NFl"��QWj����F5��:%��z��c�>��d��N���x�}d蚋M?��ɺS�Z��V��v'�ex���o_^�ذ^�ma�<lh��S�6�	`�d0, ������Ѣ�����3AO���J+iՀq����i�Q���y�L�vI�(7���Las�6QE��o�p�}}{�,+K͸�m`f���_�����v#e��D�"�#`N�z��[����s&2MQg/t��w|���@!D0�$c���v;\���� �5@��#�%���m�X��j힉`̈́��V#& � ��UU�������Q�u�*����G慑���ہ�|�K����$����;�:�} �_�C	��H�I�g���<9}��_K#�5.lb� �8!,l�?���&����*~Yw&����1��FU�_��-F���S`C�\��U�lt�4fP�\[{ݸfY������/����e��e=��a��Kե9����.���F]޳N��ѽF�_�%�.b'�E��'i�w9����ē�o�g@���j�{J4 0t��O_L	$��/%����%�]�A��Sd��<5��@�����죏�=��*4���S�U��g1.Eh�4 �o��� I�}��Rw��~��S#��y�PnFE�=@"eF��<�<E}o�
�p �S J�~HC��T��ˉK������K�_����I���ʠX&�c�$�}���+9%j���b�b�MY�*zT�4$�1
xw���9���C��	A�\L����7����B���n�Z}-��wR�56k�������o_|�����O�T�Jن5��5��No̫�2�[��|5�X���["D��y�{wuQӻ�"�ƄS� ���A��s8c�̓�V�Q�S�\�*��/0�&*�.ݿ"��)�p��a@�E�"
�����Q lu��h߁�~s1�MF��v|�䒨e^�]�Lf��L F��0��nw�>l��_�t���"����+~ ΅fd]ib�\�z�a:��*F�[��=��JQ�@S�������~��o{�����`:y����t�>"��������?%(FH%�@�{������B�?@�v4��>����5�GMdh�Y4��B�i�	l���:yK���t�+@���s��t$�_�F*��V3A{e��;D^���?h�1��xz��J�]lj��M�ɘ����Lpun��[���?�WG�s"�����r��h S�۱U$�)��� ����gI��y�${�\��w'��@�;Q^8����7�봞r*mRwަ��<�R��c5fN����4��~���W��3��[��}�"I>�:�3{���H��,)������x�j#q�{������ c�Y!8�ILNee	�J�IN񄙘c�p
*#=��^��L�@��)Z �c�����u�ي؃>�{� �%˭��k=t�+�k"�G舆��m������΃m�c@�����9>B�G�E
�	d5��V�w}��������0��8Z���B���Hy1G�E��9x�,вk�
�|�2��i�A��\��ۊ��6���Ἅ�v��Y�AL�[S�s4~�-�����32�V�-R�&��:���:�� �eCXo.��5fOBN�%�_�Q<���$(�(����|�賓G_��n�F��b����n/��P�#��d�U�� �&��a��>M�f[	��~�iL��Ϝ"{���5}$��0�3��Yo��vV�xFW��b��w�\��T�VAa��-VۉG��%U��G�;>H�L��M��a�R$��RԦ,2�@�v��t�P�Btu���SP������� O���f�
-�p
B�VɽA`�o�l��&����g�[�C|rr^��GX�J��
�$�%���UU����cL�9 u@uhO!�8S�j�0z��_m��&������d���-�!�y��7�� \H�!�+�S��t�yt3�.wy��r���U0W����G�S�p�ԥ�h|�����l�f������V]�}J�r$�����c�����Y����Pe9��.��:E!��Y�����sʹ�Yh�T��즃㋻n*Y��\�F�k�u�m7����W��ɖ���1۬����I6�.<F�	o�<~��g\\ߟ�����.�K���V�\,gʻ�t��>˓Y�m�H��W�Y�)��ݍY�_�1̥�k�[1��FW��s���ź�}T�a�٠P���P{��5u��Z�;��]M��q��������������ͨ�3qvJ7ɛy����}��Ϟ��sS�ަ����7m����}�@)����	;����B��_~�����,S�_��d62>����_��<}��_X�tH2��o~�;S���|��x�R#�=����'��&�MF(p;�5;�W���F��Q���5�駇���}	6w�1eɩ�U�ܚ�Dӫԯ���lI�1f�8�5�1����I?�%��
?��/�Q�ɕ~�q��a)=��Kb�ro�d׻��ʕ7��>�'8�Q��7��!F ,��@�	dlw;�}���`[�3љ�n������y��45O0���&���V
��%W�~��˾��+߭��NW��zja���\�?��>�Zx������2�AS���q�����u]��i�:��?�� ��g�F�U��@��Zg|�7�}D����;l��
!q����c�CB�^��RP���
W�� �� @�e��L�'�@�;CuP����Ǖ��ۏz�g/���������	���<����z��1�ǈ�,1=oŠ*e�z��)��O�<��9ad�D`�]��HU�j��&��ѭ�R�r�HM&dV��� �1��ٳ�n��ٳc$y~[;X�k{O��|X?{6���O:����^#�=�V{����߳��"��3�K� �e��i"k����ˀ_�ʖh9�@p�%��n��A�GK�({�u�]VQ u�W4������9K>�{R�y��a!�%2�g���8���i�8���	s|)7����wg2��FX������W�b�O��R�t�OO(o)7�Du��N:HN_|������w4�?"e��ZF�hW��{G���� ��(�P,f��(y�d���P�$"Q��tO�H<\��nXt$$�r#�=:���S� 1ЌE�V�D���G*��T�d,��蠠�P�]S�)B
�wԣlU��,,�ӳS����
�A�R���Yb�y�v��*j����. �
0����k	y�u�*O�	�V�d\�:� �������/���֦�5ا�:B,z[��N��X^Pt/&W�\���݃'G���e��#��Ʉ%&���הh��eB�f����RDKB���t{��J-8��r�����٩"���@�mjk��H�dD�E�S&"
QV(�����ā�*��x(��Ԏ����/>}���t��*ъc�$�,U��|�L��"7v��ʒ$I鿺�ؾ�'K��_�#( lȖc�tJ��K�5��+�����5�ZX)�H���,ŝЩ���������8$L����gSٕ�B��ةd߶<Ql�J`"����M,7�a`0R_����e>O�N��+��8��;�~��c�y5^�%��@��+��ON��B�ĸC���*����w/�bb۫�.+��)��CS����2��}�_]	ҋ��!Z
o�2�!-9�3�~E��V!T�kY߭w�z�Q��R�jр#$�Y���3���b�b�,̵����~��&�y	��E�����.e�x�*�=Ͷ3KB����8�K���C�H^���0�*���+v"�CF����z�u����{��@�[�yb�c�k7�W�w�fB~�R?H�{-��`PO�����.'ж��l���q�jէy�̈́�(�X*�fD��t��Ry�+�(���B�1o�!��ZtXţT�P��D��4���Z Y3-�&�g'H2�d'��R�:�!��?�)�3�	�)��\���D�X�>��༷��F���q��CEb\�6�#W�6�����2%e��:��j��?qGS,g�g	�,zqɎ�]:��L��)��!�^���a�H�	�N�'�����۳�>����t,�������R�O����.4
W���x��׍_<���R		<L�-�Ah[�~�f܎�W������_�~�F�ԣ+��E($4��3@J ���`_��#,�4o)(�k�g�>�BG��] �����t;�S��U#�uu�[sH��\����F�[��b�&z�D�,hZ��{2�^g0<�D��̘�{�C$�cثo�nW<��}U�%����w|���᫗���Z�B��O�6� R�C�T�p\&��(��c)�=��I)��an�%L9S�7+�ǅT��殷��6{�0�&�.g�@B7ƜW�D'���HA$����	��,�+<ft�ś�#r�yU�R[�d�|x>���0�,9�"����:W-�#���^��:��//rC���PR��QXr
	H��iJ��H�NJ���u�)r�l(r ��Ć��U[�e<z>�o������"��:�Ns��ZS�W��cII��!����#��f( �b`�c&Q����S �7!G~Ւ/QiX���[��b#툡-b�����h4*Kl28�d��R�q�Dg���B��bgER�8���]��G*��xP�+�i�O,���-��D��66n�Jc�u�t���f:��Jc�G�7	�%v�E��f�N�|�M�S�u�"��ؓ� ��[�Q�b�=Y��� t�l��Wo��l����i��V�z{5A�UM�n��z�6��b4c��u(~tF��n���W����?ۻ�:��o���'�k�4.9�2�2���Flke(��4~W/t!�C�!���Ɩ�O�����?�P���]g��d4���[�'Ḁ6:����`r�R�A�NuͩiV�B
w���^r�'#0�
u�u��G�}(���x:*��Ы��&��B��2��u!��Զ�ѻF_ �%�U#�� �m��i�ai��J؃�������T�S3�W$�`HV0�[�=��ٱ�8|lz�� o�gD�<$�)Ȃk���� ��W:Y^Y�4鱼��ã��-�������������7=���A(N�SQ$7�+�	jƽz���Q��[��� ��%a�mv^�R�+������j1E�yV�Tߩv��L�*��9�fr!u���z�o���?x )��_��"&���WW��AN��W����n-��;=��s��0f���4����6k�Z`(��o���-���ƽ0�z�����`+V�n&H��Ǘb3P ���{�[������W�;K��e�2�뷯U��|�g_�4��J��.GK�X��$�5�m�^�v8h�8ͽ��F�Z�_�ĸĕ!�[�k��ȋ����������7��I8�WY�kb�[f-2lE\��Ս�ɔ�'�X�^���z;b�����z    IDAT��$��t|��W�}/��)�K�)7�A"Q��3�4D҆d7>�R����㽃o*���w�7�ڧ@j�U�)hip�X)���a����N�F��ǧ'Ϟ����w�>`�W[L=F�	��v3�'cA���/�ճs���J�oR���Uou���A��C��S������]��]���I�T'e�D?� ��@*9<�<5�H-&F�ǌ���4A@o$TM��]o�s��Zvu��\D�:I8!)%���Z$Q1*y�}��t�y}�VN�F6�X a �}$e+7R�:'xe��$���v8���n����&�MW�N�`i \0��!r�Q&���Ŷ�s�C���#`!Q*�����¥??��P��j@gJ���|񇑫�A�`8Dt�dbZ�zs��'�=]F�IWh��w�s8���b�I�G�I܏φ� ��|�nv{�[���Rz���O;�#E�Pj�c��є�B��z?�s�H1�k���R�zm���Ǆ<6��,Fx���?=};z���Vą.�wg+ǜ�S	s -@����l[#F$+up\nD1��X0Ä"f�&�`��@m���G~�I,���/@��ր��VZYvbKx�~+��	S~�*�kōs��ȝ�	�fJ&d�B��v�e�ծ�S�Q2.�UP�pb�)�e��Ѥ�:e�~V�k	�I�qJh��]vh|UHu,�T���U�6�)�C*�,I����(ITu;�@r��%͟7�0������`�b��X��T@?�%_Őb���$�C��Zh,��n���p������]�QdMЁX�<������w���+"fܕ��Ib���F%�~qu��T�.��B���x��A�8DS���bD�G���<�Ps�fb�*��O�N������߃ څ7����3,a�vE���q���&�q6Z��a"�
v�6}=�
;U�D��EqA8c<�J�cL�Ma��Ɔ���M����:3�~؁WE)6�N3��� �r)�>T-	���M�Uߝ��l���B������İ�������:��h�U�md+��!0�J�!��&�ח���^�dO�]W�P�u�ɝ\�JNP�R��AW�gԻI~]-X�mO�T?쳴S^�g������Mn�s��)hۃ*1��ж��"�k��j:� �M�����0�n(2�+ڮ"��g��dj3mWc����Xcb�9㬫4���@�G�
{a
N��Zz��N����	 i�BO@���u�߳0���5�W�������˓�ϟ>��O�;_>�s}y�w��LWa��]� ��� \�	��L�� W�X-�i��7(�-�47h4����͖�9���N�f�%������ݟ޾yg�\���e�\�_�J���q��~��d��[�f.w��k䡝���3%6��욮iuk$�1���eJ���_�R� �×v�����]�7 ��v<�������yI�r�]��y��ȃ���/~��/Ac>��zu���%eٿ����GHޠU?6>>n�|�􏺭a��WQ�V��\@� �C�<���k�&�ժYY�X�
���E��`���Zۧ��0*Gy��S�v�Y�������O��?����nt�D��2�1��z��_��?��L�t�W��]����->�`!G.�.�H'����<�q��������6���ƹO��z�ѻ�)��g7�p����x��<ȕ��᤟����ٖB�'60ѻ.��i���0�|6���61�?l��R!!�g�N�^�S����ǌB3�A�qd+���/���gAb�3FL�3z��Y�ٲ�QrE1$C�(��'����w�����;��RK��3R�/v�_����Щ.����U]N.��nv���vvu�݅*��'��Joa�'bv_���X��u��<Ԛ����0���/�7��fQe^׾bF�&֤@��r�VN�g���b���2b��Q�Ch
��џ��OϿ����O��S�ͼ+�������lzɯ�V�l��M���4%��D�:u1�'�i�X
��#7 e��B� ��A�X�h�A4��ڡ�*���������
�>X'�.�2J&`�v�%(q��ΔhS.��P�B1����%W��myMV�8�^\�r8�'��q�9<�5��������fS>ӽ�����]rXP�8DP�]��y���)S�ݥ[�bǋ���0Cp��sŏh���버,՝	���=� �-����ۊZ�y�_�e�bW�nA%E��X���z���3�B���F�'�°������ަ2�h�{u9.��ʳ�����b��h��xA����d��Dq�ꋗq�le脌�U�.1J��+��7���7 I���iE�G:���6BC\��jog�//^_)M�[+�/{��J,���}^���XX�B���F��Z_�ث�o���j�&�F	�h�8f	O�L�|�^>&�h,��P��(��$���J>����q��D* Cb2W<�E7�f2�ŽK������|�� �W������P�I4UR���=|n ��"BSC(2;�p�mV�U��+T��;����l�B+&o��x
,�*Rl�,8G�MTG�*Y0�'���q�aH�m�2&��Lҹ~���G(C7��T�T8�ͨ-�<z˽�#m6�=(�B/�r����s u�G��:��J�H��&˵Ap5�0u�J3��Wm���d��%��6U�G�'��C�����o��>�u`��.gʚ.gWK؈de�\�i�e	T��h'�[-(�Z�!�n�\�d� �=�����d�v����ҿTb���U&�DzG�
'/�eg� ��W�Ů� �Jg2��B+|gj5�d3~ů��[�EWr��K�?��`��.,N`U�@��h.&��L*�ZPO��:���{��$lOhw����2�Z���+m���.���&-�{gK��A@�Q�nRCL��L�բ��f-�'�������F�|�V��|����!Ё�3�$���Bqe��g�� b�CM�Ԡ��+����C&K��1�?���^�]���ҝ��dT��gh�/�� 5V�I���S(;��׉
S�ӟ���njm3�k�ǣ�i�m�D����F��Ս�X��|51M�������͖�7�U�����i(��NF�o//�ӢF�QWțux�vO:�����/�GV����LS�&b�H���X�
��2��\<p�s��^�~wt2�z�� �]Up�� K�=��&Ay�kn꽭X�h��-���+�^��
"�����b�+Pl��-��mP����Og܏�8_b�����`pL�Q�/���������7Y6w�H�y,�����q��w��� )��=em9�'��2��>�׷)�O�F��b56�Bg�ۈ�����Ӄ�R6O���>��n�7�k����l�j��F��~ЈsOi�͝Yr^A,�����4�X��*�)蝹���IL�|��Y��Eڽ��a�q�@T�A�e���+UV��p #"8A�a/��|�!�U�$-�G�P<|��FGJ�Q��z{|z�9��6�����HX�ռ�R�`YU��{uP3T<}W�*~,� �%�0P��R*��� VR;�[E�3�"K;޵�5��m��J����2��?:9b��#�E����H%x�)$j�b1�j tWi�4��Ȫ�"v3� &�:g}��p|%����y�:���:C���50�,�8�b���t��1/5Ҕ^�d����L�@��[�R\q�\Ea�*�H��Ǐ^���"ַ�j�t�U��ÀX>?�`c�m���ǝ�\����r�k{��N�J�e2M=����4j餮'T���L3��i@>!�U�"
@^\ou߽�)��W�<�E��1�D�4�V������<��dʝ�n��]��Xa���e ��i����T ����s/�u%�d�0qu�h�MW6m�VNaM^��̧7-��-�A�#���:]��EDI�!:EcR2�g���}R�7�d�� P�����8���j�Ȫ��*/�Ap����$B?4c��Ha�JJB�򐼎�H!�i'��ߝ?=����r�ΐ!�މC��w�N��ݓ'�Ȃ񓸟��Ѵ�6q{�@��@�G���w7��}@ R'�
9��ѩD;ӵ�L�]�`���_�滿��`9��K<+@4Z��q$��&]�^�d�uL.f�V��{{I�=' /�-�۲��M�����6U$2�� .L�)���,��ћϻ*Ս��BB����T�(�nl$��Fl�X����N�Z2��%&��j�!�g���k��v&�V5��N�-t��o��b�apD��~�F��X]�R����A�ߪ.���,SF݅�L �r�WҮ��öO??�`��ոq_Q�5;�		���LPp:bI�΀��  ������W�ԠƊx|�uw7�rm��\�ɶ�.R������4������v��r�\]4H-�
�K��  ��{Y֬���pX�j�-�پdƺ�Ã���)�w�S?K�WA$+�g	��Û��vK��^�	6���x.#�թ+CFr��`���J%H��.��LUoş�)����֑�Vc���qgة*��;'*,�얔G�А�`a:�r_�T��?><8�?�K�=|�������B�lt[8�f�#���^.n�ᶠ���هO�N��	!�&�0~p��D/����'\�|����N��3+K�n���.���n�%���A��KAT�B���P�P�
'��.�t�rt�'6𫙩7�#����*���éh$�A�'z�R�#���)�u�?�f!�o.�q�7N�����x���t�+��y�,�L���ӓ���ףo���ۭF�����t:�w�vp-��& �KP.J��#��Y���B@\�O
��<��y#֚�O`� S�QtF�!��(��t
}�&�?�^�d�vZ��(�gD=%�C��� ���N�����|��;����<��r��Wl�Hj���V�JKW<��$&ɑQ�peR��$�zC ��ah8"D�9h�lE챵�܊��{��ص��Ϟ|����#h�za��C%
=��~dy�����`�q�	�4I(yoP0�s��C
����V�:,<>;P�M����/4/�����]������f~]H��F�QE�'�Z��#;��Hb'Q���ި�*�L���Kpu6�G��B��1U�T���@�Lm���UB���g���'>�^<|G�TGMl.6oA�x���L<�zB�E]6)��B��ܶ�G����+��KL��`���� C��aq&�:aBE�%{��.p� ��t��P��Ь:A�D�\~�ѳ�Q�v�c,�Trw�/
��. �X���A�?�ΐܘ�8�u�5 �E(c�h�h�F�M,&��ѱ��:m_ "]M��������[����m����fʣ�����y�X���$�$:�B$�he���[ve�B�
�d�:H�����j�B
��V��������X쭹�1�jh1���%
jy+���Ƨ� \R��u�D��OvS.N�)�6�/P����H���ln�.T��MTW$��<�"Q�����wW"�(���EDi��M�q���lB������^�td����� n��$uǸ�.���QUe*4P����U�+j�M�D�6�F�(���Y���J~�,��t&�O���Ǐ�#����^㭬��$3�������~��rv�Z\�ڴN�%����1)[5��QAK_�����m	F�nF'�r:
�FxqMyqhAa�*/s}���K�@.v��=R>�<Y,�[�R�Q�'C*�	�>*�R~��yGy�/yDq����R���e.(L��"gWk�a��(I��e^k�iOT�N�����G�5A��NV�Ǆ/��	��S�?��_�b�S����~��_�V������;�������!+��M����Lk��E����H�W]��w��7
���)��\���S�����������Y�˫�@#��-d�'O��z��wҔ��7Av��������Ǣ%�ht����>F֊�S{��B���j��z��?�.R�nq��RK�ڹ��bu��BE�E
Z��Fs�Ua��:������U�����'g|�8��OG���w׸�<ぞ�J�.vҧe��O�ȟ����
��z�\�~�$  ������؆����n���3�
0�#Z������
�\��ŋ�<��c���W��<~{�TK. �{�����fe�)�RM[��W�0P����v���r���PJ��D}�� ��ſ5�:o+��Kay�,Ux�r5��y�.:�s��	Us�.Ʃ=�.��aD��i��䌉�/�A7��(\�@�i_H�Т*��!<���.�t֒Zz���*�;C<w����~>��/*�����_w������`x3�\��Sb�I��F]�;���n�ig�.^1��,��}���b��O�hA����o�N���C���a�=�`E���Ã��G���ڣO���!f����֒q���T�<Р�J�<��3M@�M�C�r_��N|�sE�Q�E����
�TIIS�G$�A:j-��ٝ��ɺ�*�����D�?u7v�S'��V�8th+�p��>^W�U��v��/�r}�Ŏr�3v1N��Oœ���lX�ێr@zw����۝�|[ ��0.p�c�hS�[��ޝL�Z�u�
Z��R��,59�;� �J�*��h�7<�j�O���I�1�2�$�B8��Y���I�����P�"�t:�[�N�����w�� %��m��.hY�!p�1U����w,�z�	{#˝�ޯ��'ZHlg:\-����D��bq�����m>n�J�G�M�30���1@.�>���䋝���eֹ/�Z��'Ã�F�e�U8�\�x����bYቲ�>�Q%o��Y�S�������3�)��u���y	�I"IS1���xO�QT��ʹ"q} ��(�L��.n&6Bw�67��ٷ�	��o����K�5Mǽ�\���NWq�'�'���xk�Ge�
��5F�e�G�h���If��f)S|�ˬJ|
���0\(j	}bK��R�
�D#\���Lېa@
'I�i��P�Jۄ�Y�E@�ʔ�����ھH��/o+��wfZTn� ��[�_���&�:��ݞpBa�. �g�%A7��L�q�%��� �6;�j3�@���},��S�1a�v������e��]�9M�ݬn�g�����r[��~!p��gT��������a��x��퓿��~}�P��Rm��yY�q�r�R=Ԡ-AH��e�%��{ݓޠҥ��5 ���v�� ����ލ��0o�0gE�7w?(`C}�l�x��p��[�z�Oo뫙�y�U@/�ʐ�$�<fK4�to�9h;�W��Z���:��\)V�F�hYH��n[�E9�EmF�� B
?��"Z-��٘X�������g�~?����s�59W��e*w�޿[�Va"��)v���0��}��{��2��s�k/C��/���ZG��R�=�Y3ƀ<��5!�Hs�;Ғ=J4�������`�24C��<�j ����k�T�����؃�M���V~��~�I#�1��/�J���bMG����n~EϦgw����[����UՔX��
 1�A����O�6j1vǼR�3N��>����&���j/���6.�g�bǝ���/_������Bv�Om�������E��u�K��nw��zy�y�O��;8�V*�/�>B���P8@B��\8����Ws��n� {B/��l<^1Hĩh��Uj0@ "a�8j	X�K���")ߑ&?���q8��v���u���W��œ=�0%P%3%<���˛9�@q��7�"��̓F$&�ٲ���n.?��F�I���]���i�^a�U0K�B�5~�x󖎾hT�:�Mb����TP,�"�(x���������S�r>��O���(?̉zI� �!A������7M{)to�wp�Ӱz6oԇ�h["N��S;���=��N��2��ǁ���i�@�(��|h5�    IDAT%��Ax�X����Z����4��4ڠ�@<����'O����`�x��:k�d�q�/�?��A%�����ʦ��*&���{��.��e����ziM�yk�����\S�n��ڭ&��*�T���[p���{dmC���uSA���]rd�f�[�4��w-;&P��^���x���α��\�`�l$^2�����VZ�ŗ���fD�~6l��p���t�I�\\�$|��Z��Y��U͛�=}�}�pG']���R������-��]]���o5���0����4!:zG���?p[�{�T�W���7����$���;��2A@���?h�a��|��z����Pm`��BYU�7�ل��V $����Y�V���K���a���2	��!�sM�H��$}��nX�$�G2��}���,x�c!/v���A��������8�]���Z����pr7�aб81�h��'��|��-4�'z;���/�`�Ai���{(E#k�p����o�fe~U�R��Vg�}i-U��N$7��$���E%��ͱi�1��! ֓Z��胦���XU���WI�:
Sf���8��Y3���[)
i��A5��@i3��<���+Q���3 �i���)���dgJL.?��F�6�u@j�l���?9�=�OZ�SVh(�j-/i�s�O�b�<^�|��G�DFJ cO`�@� �cQ0|��(�)A�J�{�W`��7C��G��7s��Г��7�#M��l�f���	Y��ٓ3�yy;B� y~�b<%�yZL��|���E�����<h\���+�����������k�K(n=�5��$5��׷Q��B!�.��XK4�񑋁�g�鼠�
r�����|i���\��㛇�T^)�C�D��F��]���P�.���zB��v<��YM|.�x���0���3�F��!7�
��9$�3�� ;������Z�l"�vFo��c,������X\þyĚ0�}�Ƣ����S��'�Aڤ��;�0120�hz]c�k���O�_]O�;UF�����X�0�,hhia���~��,=�}�y����:dNMY����2GQ"�*������<9b0���@�j*��ZᨳL�IRG������҂ ������	���]U�ᣃ�u���sI�+�{h-2RUVV�@����,��5~�} >�f�F��4r8m6�-эB��ԡ##3���;�8��(O���=�h��a����$�Q�]Sf�X)[�e���n]�'u�f�\`��:72IJ���]"?�uh��`��%�~���JP��V$�h�K�AI"1��(u��FB�[�!cNO��r����}���O�_V�����*�� ��C �`�>������B�Ό"�_׀p�B���� ������A��@�s&J�ZA�"�{a�F\~��~�O����[!�[�nh<-6�y��4�P���mR�.G�KW�N�O�?~���'$.���f�X,*;��\�*m��G���B�7FW;�df�����]�(;A�|�F�zM3�Q|��d�����DH���������h����F���F�Յ�,<�v��[_爳`������ qN�(2���U�t����CJ�7Ǉ��Ios��kK����"��(��Z&��f�X.>Ʉ��,\�|��ص�b0�®�S)��c��(��
���C�����r��tu_Q XO��nr��F��֨i����v�m$�Ŋzd�*��d�z@rqUTh��"��M�R-8H�P�L
W~ǆ�8W,�s��?���u��^�?dU([a�-�z��Ϝ�g ;���Ҿ[|����3=¹�@g1J��99H�������J�Ǉ��-N@e����!��".�6��+73�L/���PF�Bx��Tu����H57Ύ4F8�]^��y?��r�T��O�0z�1~���PS�q����i��+3$��V�[�qx"���A@%��X��#�|y��åBd(�EV'1^i-#��V]����i��_~��O��{�T�,S,(�/���u#�x�"#��3l��?��qv'?���"��H�a؄;�\b�W�_�����"c�܅ѻݽ�g,�=y�{r��D�ٴvgm���>V9�c���]B�ngsB2��&����(pm?H�Wx�h��7���P��P����=�ܒ�aSms�j3�r�g�%Y�xo�J��iz7R�@�!�T������{�:��_��OԔ��wƓ�W�)v�wo�5S~\��I������s��h[����i]c+a�?o.�9U�8^,�1��3�x9��鸃�8�ys���|�}�lӢ���'��Y���R����y���,/6Z�+�?��)�Okv\�.�,�354���'Ym�ް�WX��WG`K�Xo[���}��NéS5=�W�F��!�gq=���f�9@y鞋�k0`����77?�ׯ��$���߲��`&~P��4���Z}ӯ���@t��/�@�e0����Yt�{��Ͽ�����w�y�j �Ag�?�������~u2�������Z���NmyK�(�v!k���z7C��IMF�h/�H�@�o�}��b1�J�I�^UnF��O�y~˃..����?��������,�)�8��N�ה���N�>]�7>g?��K8���p�8�G�W�K�˅5NGR��Ϯ w�wy����c9�����/�h����_��o�ֹr���cd\�0�T�z�����8��?$���U�V*�뽛���O?����;�R~�g��� I���8�kEVޏ��h���J�P[[�_^��^�8p�y����X�ҘHK<D�#Ma�ކaL�b.�uV������Ŧ�9�0�
������_,Tx�h�xe^��T�]�?+F�O��������������ӿ�O۫���@̅N�J?�i�t�tiH�uM��f!��ZM�.Y
u`�:��ۤ��\�"$���{��t��3���gϿ���|��n��V;Ǻp[��[v��'�ԛKEM�����7H���/�=�����֭��%�Z�kl���h��L��	=��ZV,�F�T��W�x�0�6>�Mx?�tG�~v���܁ʱ��dXn~!�}��#��V�_��N9�:n������Y��PV,s�ו��C�i^�V�ٜu����o���J�s[y���+wz��U��� Nv6D�X]�Iq�Z��x|��Rk��[J2����M	�7D*�sj&��Pn���&ڂPz��겚 v�HP�Xwog�۫�B]bB��DA��{��V�������ՕL�t�ۓwl^���j:���A�z�p_�vrzv��ߑ{U��zd:�/�t�<�v�S�N�5����,�;�������J0�uЯ+���b4L�#��L�	H>c�=����$6Yc�N�"� �����Bj+4�A�D�:=c��^|��@gZͧ�%g0ȧ@D�K���3�c�!O�zu�I{6�|&�+������O
�� ��}�Bg'��e)l,Ts����w��*�a��*~�"	�nX%2_�������ݏ���#�@�)��TA��I�槫ʆ�۬�q���CQr5D(B�`[�hDh��R��P��X4��$�b>%�5)f�D��g��O��=�FGg���ˎ��$3��[$�:�Mprr�����)�4��� �%�_Y!�1���X����bI3�}��pD���m.��
�(�z��d�T��*�w}��_it预�O�C+�az,T��q]�]n�jM��E�fw�gG�{�O��wT<m?#�Ǥ#A Ѐ�mZ(#��o$9C�ƨ�Q����|P�[�#�@�r��`��@:ь�K�/�_�Ņ`P�,`�M_\6VI5�7����a '�Q�~���z�,����T	5,3ʜ���X���`/�d���J(�Z]e	ë�@��h����\h&;�fc0���W�������m�.R�6��S���B��`|`�<{��o��u�l�@\���d��Ǖ�а=�U��8v�$$���#/'5a�"\#��L�8dFd��˘i�?�N�
�z�[�vc,�`0Y�0� �	 ��L�@�J�5��+Jb���X�b�����V��m�?:��%�⌃�!�PYs}��� ���Y�k�������V��M��gZp`1n���ǕL���I�Ǹ_]��	x�۝ѩ���m��AYѲ���\N�̠ I�ؐ�5
���G�U�jT0B�ئCv��;�Ei�r:9aE8��9�$M:SҸ���FJ�iTr�	��	�EZ#kL��eH҆P�Ŷ#���y���FE�h�v�sA����~M�W��8dv�?^�R	�G�(��bez��|C gO����N/?��m��~d��Ӄ�R�|�D��v�o�y�qd����{���kL���f"]�V�4c�"%/�}��]��ō ��0�]mXWW7>��W��"[��b�yz���
�y:�a�gd偊@�`3���%�g%B;ͯ�x(Y;V ~6�o�Q'���#c�àp�0Jd�<G�W���	 �g�����\Y���9������z��̝��w��:��Vg4�"�r	 ���S�q��x�æ&~�����.�L- �uL�7��¼�́i��S�V��}`��Ղ,�sʵ�,^b��Y����7c�1[�v��p}՜��X��[~���%�X��1χ��9e�F��@Ћ$��7��po4�rv�$Zl��VS��@���Q�AЈa
l�Z&ر9�t�l�֮HL�����`n
|4�b%���yK)��x�o�w{��	�>Z��b-�1�!A[�����r*x1"/�$i>I��O0?�&Giz�Yˏ��Ƀ���Q$�R&��Ѩl��z�-1k�[}�(L�)3GQς�����~#C���|Se�o�"��FE�E��	�ٳO�=|!�XM��6l��/H�@k ܇�&�$mR��3!lF�"1&9�A_*X��v�ws�������vlօx����BˈI:!.��|�/:͏:��P�"4��Gb8�瓗d�����B�`�����wF�N�\��|���f�)b�� 柟r��?s�^����=�փNW���>�wx*y��p1�����pG����X
�g��zfZ�	�#��`_]`(�&�����`�	)��ȉ�Bg�o�c��ơ���VL�L@.�k	�K�����$ȥ/$]V*�@�^7ڀ�-���7+m��&�~���ݳ��ڝ�*iUdf��`>(���C�����+�"��(`	�rq)�/qG��D}��;E�M� @俢��{�(CP5�9�^��cZ���j��d"J���p$���]-q~x3�$1M��OZk�v�_��-Ԃ������~Ae���]�d�Pq���GĘ�[g�|"#,��\K+�[�\yv ܯ,���8����dŤ�\F�C�J�$	�ӫ��eb6��YI��8��5��<9��z��|bԄ(q�.n?%1	�@y��Ǆ*�����J��v�����t��<}�b���s�!�8/�2D�0������K�\��S�l߾�}�
a\��ZC�����C�4�(l���#3�w ��ۘ~��Gg���ͻy�nB%��$)����V^r:����t���A�5��><P���bK�y�����;<�����D��V
ڞ��Q
N[H:�OxD�9�O
��J@�di市%��:��	�M�s$ؐ��2�ur���Q�C���Do�L��M}�~g#J�v9Շ��Z��#��c��V��m���́����,j>���S����T���[zn���6D�`W6��qZ��1�����-2��zw���?7���Zm��h�YJ��A�_�
j��GA�b:J�%�.�?� _���t$8
�I��ګ�G��D��?cK�d�X�TH�a5�H��
��,�ηû�bi��
�Q�lؓr�1&$��^}��0e�a��BM:)��aq��.�A��^$��~H��@i%dĲ ��gւԤJ�����8�������	
�Y��4�ȐL�,t��0����a��k<v
�Fݳā���)��	$*a�o/§�)��`JସI8�Ҕ�ڴ9gQ�㜬��˂KS�k�_<�
���`���<��5=�]��M#"��H9㐥�XIۍD��k��gj�Q�j�wC�M2�z��#�֙rbs!
+13�y�SfK��JM[D�)���r�����CA����Ţ+�+�3M�N�@J-�
|���E�"9?�L�K��Eo������'/����{�t��Z;I? �Q1Zj�1�����{���|K�v�}p��Ҙ��|y�-D6��q�a�$ɚ��|��6?�p��%���$�2?��H��G����@M)�ć�a�%��6Qem᝭�����6;Q�X'>h��@��L������Pd��G���M��e�f�LO��P��
%/���k����)s�핻����HY� �Y�b �H
qB��:�_����mE���ÓA����f'�m�`<����Ьb�pP�d�d4Ex�_�Ņ;z~^��2����y0������J��oD!��`�WH�tl�,ė@z��8y�t�c���*��	�<��>�����u
����j�J��%�^HbI�1̉���J��7�%����?�����ˋg�ڲJ�Y�Ӗ�<rQ� ��%'�2p���3�.�H��#��n�U���2��b�n��]��	08z8xyx��Ԍ�_#�����dxF�L,R*8%� ��d:e*��;?OL1���2�g�?��?���,��n����˗Z���[���O�S�,����Y����t�G�����d�:�	�W�T�{>8�N�	A�Ow�Y��k/����~��9��/^|�����>]��i�͸��x�?�/�W��n/OO;u|v��կ����ϼP�P���ûQ��F)N^ �������LU�C�I����Q��3���RoN�������؂�����߷����{[4��yﮮ��H:�i�&�����ս���{���x�6ש4�0�;U��p���b��-���ŝ콦=�8P�|XB/3�(��2c��˅	�%&D�.���d����w���9�S��t�5���G���b7:�-���p��|~�9N��vpaOs�Ҿ�����r/�$=�G��-G�.~��
�d�r8��@��捎�5`�q7�����T#wz�}l� ^�x��J�Y��W���~�N�ܟ�G��88�3�e��;=���d+���5�h�ϕ>Lv?�/f
1�����0ĺ����7	���w�+��ڭ�V_�ٚ�P���ܣ��W
X!�E�rl��9���^�i�vŀ�P0%,=������K�/��q�V��.�3l�5�$���Ț�
k�J�?�y>}�;>=9�R���XN�ϳ7����k���9B�Ř`޾0�b�х��Ղ�J:�P$����;�t!��������͓�jw�����4o.��?2mܮ�?�q}E��ԴՌ�-KO.&1��Gf�{?=Oİ`y���!F�&B�xRb�+\J��z��N:"V. ̧tei�So����7�����^�q��)��d!��>���8��b\��)Q����8�_�r��CO�@����E�/v��l��l?�w���#q�㎔���imvJ$/_�O���2*�ê�%�U��@<���W'����w��?�8��*`����M�o���LI6'+=V&G}ݧ�;�UNN�iZ����3e(d9�#H^�/(/���2��{mE6a�+R���=V.g��:j�r�<h<�#M�K�Ȁ�Joc�<�Vf�!�T���xG1��]m��;5^M:��C.F=ph�;��g	#)��_=����oC�}~ސ�G/-|�G;��88Ѭi�_EY��Sp#vaV{��T��B��f�b�;��a��%���w�c��&Q5��r��̋q�V}��"G����d���	���B�]i��ap���Vp�����o&��m�_�    IDAT����>q�b��뎶U��7��������~������ԝ�cz#�Ki`#� \)�BH]��j]�|���� @�؋KA��iQ�P�X�l���2����29�Q� ����u�-��[\����\�A{|t�j2��.�9¢Y�� /��R��gg�T����t�P�'�L�"gLZ)Q/�]B/�i�\�����9�tL;7�s�RV�5���7�=�>]<�)!�C1 �j���T+�ZnfI\O2D590�y�1�ً<l���.�|Y�7�fn/�VBqO�`�G�K)�����!�r+3L"Q_Z`1`ѱ��-@�:�%v}'u�	El�n�	��F��Qa�	 |� "^�K����L&Ig 6h���V���|�=��ęJM�~�n5�Ȟ�����]�T���`�a�<U���R#�U��9=<��CQ�h 9@'�O�T��̰oGyN��8�K��65�7Y������byu�8=;������|9�O����4��Lݾ��L:X��G��_}q����(Jiw�h@P]�g
e�ȨP��T�0�+t)��ޢ-H�j-�DA8�M �H�Dv7 zа�Gd�:��E�偈��"���r,E(#�T� !󆯆��,*�Dl�����{^��6����L��,��=�p��$� e1A��*s�ҀS⣖���ވ�݊)����v9W/����f$Pi�����"?�.����?�ȿy3������R����h��g'��>z����}��W�����u���䛬o�����N91,���d��lk�T�B._K�+	�'�,-�`�D	
��AIM�H[vJ ��1Mw9yr�a=����~C b���SFc#��g���\�D��F�]��w�A�q֯\�L���BY��!FhKnB%b� ��X"��xۦrp0͗+�����W{j$�89����9����\E���?���-��Z��U��<�-�9��2J�j�4D�'�g��ӹ�[?6�00IMdn���-j�R𽧃��h[����cjt�^-LrTRhA �g�RP	OL�F1M(lg�H4ZAv���a E�r�䎗���4tPI�d9�u��樤Jv���t�t�|T����&���sٟ<�M)Z��G.19�K��p)Q���jO��s*J�B����4�r<NF��n��ET��Z�ws®����~�i����w���w7�\���_��z.��S�m�����r"4ZEI�s�-��h��*�;���w3E�t���$E��7*+�9�ɾ�ȦX���-�Õ�Q�	Яͤ�5&�`��LY���?;xѸ�9t<��(/'���"��׶��QY��֊bS��)b㏣����</\��]c�N;A0
K���X����(�6�4������e�R�p�W���x�8z���ť��H�2�����o ��Z�7򣗳g#�#��z�N�]��Ѱ�yab6�"��N/ź ;y$��K�#/��,Cz.���4���;c�p9�V�s������-�`�������s1M����"�`��6���@�hhu*j��Q�D���:��O��p.c��k��8A�F�zω$4L��et���5E��F��&�|�O4˓ñ��1������v�Rj�az]����H�"?T����{P#	�$eVj<9³���y�fU�?]�R��n��h����9;�����|��A����9�_k"�P(��m��W:�~�T�=`����'����t��*�b����h�a�
'L�Ay<�3,�Y��� Ҷ� �F�;�{��Aŭ���$�)،�PcdB]C�r|�n�{�Y�:;n�_��v������Z�\Cn
�(\>���9.�h̴r��{�O�g�*`G���`R"�XY���+�QJ�rn47�&�<yU���Ah!k!�����l�=�P�]���܌���A��|E� 4���@�xXǄƼ�Qia!�&4�͚B���m�`�v=��I?hn6���SV�>���$0��'U�N��>OR
�[�v�N�3{��=�=Gn�%촏ڣvKaA,�2"nķ������Q�4[��`��y�3)ID�0�N�8~�es"6���(D+5�K\M�50=]���������?ߠ��!��;9> �S ��e0��5�}t�?�i=	B�+���s�5p4��b9�fo�h�(�A�ȫ�L��pj��!^aN��2�y�*��Y��t�J0��2�\�!n6K[S���>�I�h�/9����l�I=;9&Xz�㻋~'A�m=܄�4�smW�	�J�8�"��4�����qɔ],�y�!�AܜL����w��� @�!��Bu�0����c�VE9� iL�҆���n����}k9�<t�ű���|l!�!胯<1ב|rA�qe�[\�>�������Wg����7�*6����[��cEEY��i��ʬ
*��%�[Y�vrB�$,���MY2h{��*��?�hGC�<�U�$���L�-�q;m57)35��*�U�ta&�Y�pm8oH�Z$��	�@��_�������ǫo��aE�B��O�S�H̦?sI�M4�^o8:=��n�W���6�	Qڕr��\\6;%�
����B�2�O�-04WC4Fm�����*��Z�j��h��/�췹���P�*��H��<&�[��̉e�NN8�
���)w̙*U��q[�%8�FF,���<�}5:� te�~R"o=��b�Q�i4M������'<4�Y�z[����A�|>ej��Ҹ��x�46��	��Țӳ@H3�
�6H
U(�����v{���m�����}�b�/T$�� ��ݘ߂� �gq���k"�9^«��+�p�=��I8lA���/�{5����P�Hbt�La/X--̋��8�ry�����
[j�nV;`�%G&�-��v����r���y9-ↁ">&����I����o~�����۟.e���
��5�\H�V��1ޔj"t��Qk[]	�)⢀���أ~*G����tve��}@�"�<p:�$�J�=iO�_^���a()�F��vb�q  6�l>֫ML	g/��J�\c6���_� l�ânp{؝<�>С �gӦ"�o^i��:���zbw؝ޯ��zȠ�n4�H�	g��YO�:n���VC�p��,�ŝA��;	:�/�9��+J����Ke!���ƳW'������v:쵏���)�!�Ǫ0rVӄL�����ޘ��B۶�����zqQ����we�jI���NP�bWS�oO-����]��D�b���JO!�0���X ="����?->gqzs�#6��uAy��m�����<R��	a����29�!v<����v�d{bgl/����u���~y���7�� �e%���|�k\��r=Z�&;OU�Ȫ�F���ܩ]!r��쌆�	�Q�ҟ�'>|
A��7���z�l�N'Ϟ_�������������C:ҕ�{��ս�%U]�n4�%[����DR��5Hh��IFv<�B�:�9�G,W!��*���( �\����L*� �۟����1i!��;� �%C�ǃ����3��Ú�G8�^=3c:�ؗ��]��͜\B�@2��ɋ@[����yA�"`�g�ˉ���w�<�J3n�fHκ�\����-9�2��?˳nq��v<�Ľrr4��w�,jNMH� �j{��ݛ7o���r`�����{/�����\�4���,�.+1��'���Nn�����|�Z�_��2����?�>��_�}�h|���3t�������[�?�'�Ţ"��@�R�R�%����ӏ��Ma���n�W:���jO�^T�B�6��������>�H�న�����D�T�eS�ppFD%�F�D��FUvw��%���Զv)Jl~�a�=���fv�.�o�������n�l���j������YU�������-��]��h_`��c��a�òȪ5�<B�j�^e0�������a���)� �L�~�N���j���yEG��F`^�&�`�_�*&�⫥Y)3(�^�%٢B��8�)He��MQ	f���E3�x�,��eUؔ7��-�����vV{�~�a6'�>���ݖ̕|�8��wAZK�٥XE�����X%�-_m^˳&�-P(3-䭈���
�k��?w��ӀBD4v�G�ׯS���es}��b��,WZ0ioa+V=�:
%K�=�a��u���^�=�IZ
�"oWV�j�O��Я��O�ִf���|��$e�t�ȊJ*���Բ�l�s���a$���#Q.�����P�~ܝp�p�a/23|��լ��5+Mi
�'�*;��^���~�wEx+���U�˨���kZ�)���H��GJE=�E�qX��@�� �G�9�9"�ғA>��	
��R�+IZ�yԝmG�=�!E��E�;����P,�ŭ	.N|������2�l,��Dŷj�gB<8jT&	�Yh�o�i|V�\7����E@J����������w����B���s2�@BɈ �m��v��S���'j�r�<<��*m߬L ��:�]ȋ�B� ��W_�jn�Ԗ���|��Q�N$��F(M�4�!B�>��r�3����@�,�%f�PN8,G��!�.��A���H�?�j����]\�[)r߼{����_��X���"Κx8�%jkw��{����{��0�-���nn���%�>5S�Y"l�G�s�׈Ԋb�4I�4'ҝ�Ƌ+uk+_�>|��^~���?�x��L@ЏF��^��n}kM&6K�R�A��G�̱YE�98{����w��iu}c�ኅ��[�p>_OI��q�j���B�xΙ��H� ���d�1�4�6G�� }�>6�;j�%������������ה����Ҫ�p=��YPf9��,���z$ؓ�$����o�w�� �9�(:KƬ�cFsf�A��0Ne@�U��3�'',� '#f+��4���K��v/_�	�0u�����/.S`�m�������-u����*%������v��u,���u?�<_4jw��O��_��8�4�/o��;4@P�g�K(C4��|��L��L��Zg�����g��U�WbBHR��ʹ" ���9!�@M��X@�yr)� $�O��h�o�Ĕ�S 7���oV 3����p�Ǥ������]����kφ�*&�_�S&���t�-�t��p��L˔aɸT�hs���j�0I��Ϳ�ȷ���p �d��)y�9��=�T��խO�Q�w�~{P�J�臇<Hē$O�U(E����~q�]��f:������IG��8��t+��DY(ݡ41����#t�;���v󑧡��	��҅���_b����,�}�e t�����LvC�K������o����?��ɩ��y�7���t��6�	Hc�o�d�Ȭ��y��xI��S^�W]m*�È������>���z7$tͪ~� Z�>��b4�����o��ZLotC��J�u���걠M������a�r������L')V&`�F��r�Ѵ������t��Av+���^>xn4؂zP,��2fßa��y���YY�P�4��M �,�M$]q�
������y���vߩJm��
�s>_��R���҈�������&?S�s,W}	OI�N�ܨd��l[���b%Sm�dV`���w��,O�w�G��h�Q2q?<������|��A�=�ɻ��p���q<^}z�,�n�M����IB���!q�Ȱ�Ĥ��Cop���n?��;�!��[ON	�Ft�Ε.a�q]���4�Do���,��_W:�m����1��&���-.���:�g��G����M���p�{��W�@��aw�J����VV����r�ZpBΟ��MzU�ѫ�le.�"���G�Mz���O�����=<5�ܫ���=z�m�ŏ0%H|U�ɽ�Y����2�+\��i<�+{&JY�����F�A�
SS�a�atrݥ�2130@@�9�t\�@%G �����K;�(�� ��B���
]\r��~]f�� ��l�:[>�|�������G
�� ~8��Y/��B���!6��Wr�"��5��*u������")R��Nh��YG��s�	�Y�J�����T���D���q�W���5I$k�G��|5���p��e�`�������D���8����~���tEHW&��;�����Ļ	o�d)��u"'|f�
h�}p��V�}����/^�p� e0/���{�s���#i�A�f�Zy��k�	h�S��<V���0ƈ̾�L+sP���'�X=��M�WH��F���S��6Yf���~*��t���.�������INr���!Mw�w���7T�P�A���dO +���ʢD�����G
�"Q����E���k��-onC=СD t6�_|����S��?k���R��(I�pM	y@�C��[��Qf�YR`/�
۔0��/R�nsH�\4F"�:$�r����@V[�^��i��u�[��ꬨ��H��w�?�+��&jPJ� �!�S@���x.'[@�P��p�v�_��Q7�ոz���"������Z6,�!B����v��(�YiP4�jX�����6[��Ɂ�]-/��!L��F�/�y��E��杈f�S`:�'4���!=`����r��`q�<��B�bi�g�G�Fw� �?q�7+C��i�-������a.*!L�{CQc6u�J ώOl���v��bKF�H�����+	���,�9�X�D�p��i
��XSi��f��_q&F����a�t�r�$*k_�w�&�K+U-������8�MkJP�E���z_Ɓ��w-�SfV�9.��Nʥ%� ��h�����	��vY�_n�ش�7�T&y�����wb�׌�aq��RD�D���&ʋ_�	�Lv�I�p��3�q��q3n�H�}��G5����y|������@i���C�$`���,Y�	�n�����=*2������lfU��A_�6�J�
' ;E*:�*�S�ӂ�Q&�wC3�Y5�ay�/��=����*������H��t��EWS�2��+P��6�C4�a��5�mne��q��3����zML��n4<|~0y[i跒��R؂ WIv�
-� ><xH�.�H;! HM�f��]N�RK^8X*=�t.��]|��W�|�\lS�Br@&<)D#�[bC�Q��Ȍ��^xGw�%&~��Ř���$H�PL��ٷ��U8o��St�B�X�XM���q��h��Y�Uкl7�����|qu1}��v�l�64�^�>MI;	u?�¢d2�0����?����a�9���F�6��[�b����"�a[�F�9Æa�$�
D,�D�e�\ ��|9..1���)�Q�+`,Je�$Jds0:����Cv��ɏe��S��ag���ʓ����/><^�j4Nc�����"���O�:�%pC�"��н���`�u���v�޾���*�]�&}c7L��t��~|{�[�O��pY١Y�Р�	76����J=}k,SZ��[]��bQ�+R�⚀���A$db�y&S�5K>#ļ뭫�ԝ��^%����8]�"�����g��/�J����"�*��!�D�]Y>=�_�`��<ٴ"��Z�G�+,~B5Zد�:t�3@#�Z��Y��r49Vnor����V���6v�����<zP�q?#x�&����p�X$���;8�j�J��h�8>:io�O������2�]1��C��pm�p��t���d ����f�O����	�͑�&_\rR���c��S7/(�Z7�t��El(Ȃe
]��A[�X��>:c�3��m@� 6�#�@�[����'e���,��2g�����ӎ�]Y��Ny�|r9�r$����9~��9��B!����7� 3��~"	7B��*X��z��Dr����f4hM��YM��������/��HJ����z���孊?쩉�|Tha��߾�Gۢ�w��y�vrz���_��������o���͵�TD˒!$�B��.,��    IDAT��yk ����`2ַ��S�J,��b��V����4���'N��X�q���ճ��D��ڱ�шT|�LNj��� <5=g�K��l���V�>t +�# �pϔ����R�T�F ���Ͼ�1/�\/�lN����7��)'�A���)�q���%z\yM9k���c�����.��f֍~����"����4����k[�q�v�x^]���DYt�׹�ݽ<8��ԇ<Щ��g��r�>��&5(�Ip����C����7�y��m	��/�%gL�YQM�y3��S�Wˍnw�{�*�V�*�p�܅���)Nb�ȷ/^"f?^�3��T��l�&�{yw=�u��}��+��X��Kbl-FZ��}rc�O�
2n�����(ya�TNFga�\��-��V����T'T"^����^��=qv�n����Hѓ���V�LF��W�����$r�V��і�|�X��to�5���Ct�HWU=M5�P��*4�4�,ÆM����i�5��E)+�&iP�{�����a�Xz��G[�`t�mU}�=��7N>Ȗ�;i��U��h�2U�Or��[��m�>�o�ۏW�Ww�y�#�'y=&��4�;��t�"�$�>x�c��'f�V.���C�^b�#�tK�9��b��t����u�)��}�ˊ�Ȭ���i��sϻ�fu��<-#x�+�NBҤp���+�oY�5ڐ��	`��g���a����&P#�Z�eW�/u?H�(���m�
:� H�"�QkT��9�\]^pV+\E:'���:��4鞼�E�W��#Ug~=Ì�eu�?��e굥h�,��ޭ����^�z�4�o�� {������x�4�Y{:��JI=4#��  �T�����ӟ� ���m�mĪ8^���4D�5L�RgZ�V�O�(Vm˒j�Ws��xF�TSt{暌Z��8��~o�����Te�%̟M�G����$���O�Z�a� ���4�a%TP�
WR�3WSeRp���fJ�LN4l7��t����"z�f=m�X)�Q�fP�T�$�,�ꢷ���[x�J�0831;m�/�_���:՛C$=�2%"���-�;DA���UQ����`�֖�_�`� O]�bae���M�ϳ�0����]u�h�l���W?��d��2�/�I�`;!�H!e�>������'�
)q2��@g�4��1����邶���6V�8Y��)��8��LW��f�O�+�?H���N��X.;�6�h���nM&!�"����%uS���ǂ��/�/�꼷�\��XV]�ons=�X��Zp�9cYsdΩ���IZO�1D��J�		�A(�<X��f��i�j�؄����;���2>}�~}�`X���d���n�
O�1%�S�&2]{lލ%!c�&�Z��V|�*�H��NPn`���j��0���f|�7z�_ڱ�N�E�̨==0�F_��+�f�� ���d���~��&nC�u�/�:��'A��,�&������ZvNL��������o�y���:�uD�&	�Vc�Bz���R0�*���L�a3[�n�g��}
C�~V�j-��T�KՏ���\��n��~�5|���2i�jWg+��T}�0?����nys�['�5��>
�+%1֬��^��_��'�>����_M���k�|��aV7Ɉ���ڣ��2;��,(K�����K����c*AdX�ӎ��������٣8E��k�n�RV
��E8�>?y٫��u}��Dj��o6�ӜA����x��_���F�O�g�y�hQp�^�]��#Z����U�^
V��vM�g�(�0���:4�4D� �>,�{�#��-@,�/�M��ArT�0�����5���u�5,�2N���#G9����2IM*�}U˯z�����[�<}�J*SJ�Q����R���;i�H��{�U�c5j��a�L�p����,ȶD���j+ �<���{298>W��*xw{�Ȉ\�Ç.�Y��U���w�)ǅo�g��Y�.7]%.]�Eh��ņXK���2�lC�G6� �m���n��l��z�H�w��`	Ki�y<�kl9�b���,E;rE;�DY�T�0���d�:������
үϷ��U��)��[W^�%[㶞//��D����eL6��{?�݊��=��u�Nyށ�Mp�1�U[�!͓�9�Ez�`r��H�
�R���T_Kٶ>Z\r�� ^J��-yP����f�ntCnݕ�_���z�enחIj�>���Ο���.��E�3&�K�7�b�IbAQ���U0��t�T����HAE/�!�(���Ci�%%U;Vd=�}d戝�V���MD��y���D����'Ȥ�b}+[g�ا�*ن����nnz|�Z��;-��_��� M*�<�DSg�ZS���$ �B��P$T�۝b\��mg`�<�B����<4�+�D�����`�/#P������2(h\�3����v]/.un�)F9�CF]��g}U���e�M`1Ơ�ҭ;�6v���s	ҝuL/=�R��JSr ���Z�iLH1af	z8��W���w��ЊH0�$��?�a5�r+I�"�������d��܆.e���tWbڱ[!N��%vE�0u�K���w�YI�>O҂;�y��n�n�ktF�,d�dO���A���)�܈�S�]X�ӵ.bt�4ݑ���)��7$�1f��R,e^���Sk���k��uyBG������c��(n.�+ݘ�}gk D���S	��F�X�nw����'�$�v�y��R�v�e��J���*7C��'�>��w�Y����jvH��P��o\�f����)KEY�#���rd����a}{H_i�T�)%?�Y!��ջ�}��yq]�KG�b�Zފr-Q{>(�+�d=��oإ��r�;�d�ӮWA���2¸���́*���?�͞�|h2Ɣ[�T�K:99R�FQ՚!b����W�D!� p�QS1�yЭMN�������ɦ�*� -!s��"���Z�D���qb�<D�VD<�#@+`M�I�x������K����F.ئ&/EC���֊M� wW>��	ڤ����N�i͒马\��5�"�f��mĵ��*e}t<��I���u�����M��v��z�ڰ��{^�n�m�7���n��]a㵢W�V ��'ʮ2����F�:50w�*9�oT��ãzw<���W�!��ª�bUn�+1px-�-�����h�`��d��q������3A��6�i	����H�p�Fs��Yȑ��Ĵ"���F��Y��F�	ᡝ��Ge����Rf�@���D�����$q����z1��[{�.$*r��e��h�[Ov���̩=9:R�����Km�j�6X���?0�5T���R��ĵ�:��J�5���$�aP��h�"k�Ɠ�#�a
{��h�\����=j��[��6�{|�S��	�QO��{)L�LDO{H��!�),�m'V��
8cC�mИ��([Җ���fCޝ����hN�v\��b;|J;9����iyf�4�M�����f�����iC��X 28z�i�"獡i�K!�8YU�PLM.&;���u�t���,��Na@񵭕���3<��[�%	;Um��ɱ�af�����5�m�)F�2�8v{����N�r����G�c��Gu@��Q�CH�R�L3�'��<$������V�N�O��UA,�Y�����b����dEAX �|�S$�L	+I��\��28�뇌��w����_�:<:`b��L��B�cx����)�`V����\L+�ÑC��A0!f)�i���GL�i�j� B�1q� �g!��<�c<�	o�2b���΂�T%�^�S�noS�Gfa������[	]�QS��B�M�W߼�q�U�����j�H�����r�>�L����P��dU��a0NE,�
���T�@�a���S.|�ļu!��V�*̪���=+�'����-p��}u�`�� �� ԍ97���=���ŻݷU=������Ԛ���Jk�"�V=Lo�V����O�U�ҧy�l~�U����<E1�ږT����������������p�� ��z�#F��]�P(fŋ�S��|Z��C\���S�����p`k�ྉz���vc,�a>;"S�ݐ�^0���4�(�60W`��6�=���F��lA9���S��n�m$���ɋ3�%�ٗ�O�Zl�n�@6���}��n��q�e� �=����r�F$��pB����F���^���3�z�Q=�������W� w�}��換��y���"`�ͧ����|6X(��ΰ9*�d����H2刴�\�#Uu>:�t��=��b�YԪ}�Q�!bVB;��r��u��r�S#A𸱩%ږ�� S�B;�G�A˳�"T/�+��Q��Tyt�� ˹ز���rYy�oL�#��}=��ܑLV�)�)$��F���O�|G\�#^����縋I���o�P�-�e��)�F۲tBa� jh�H�� �݌y�I���cm���;}ʍ��5Bٺ�Y�����^K�ۍ��O7�0�\֯/��O��>�1�2��>6���
��g������X����t҇��9���=i�J~�W�O_�JNዟ����W\l�Q�Q�jƬ��>�i��r���X�׆��jܭ�G����h_�j$%�SS����.t�*�H����䤮�p&���<G�c�5����A�,�s9_��/������%�S��r��Ys���]ls��+w��;[.y�����|H�hT<��_���?PU\oS�����e^K���q�tU:?>>�Xwq�:(�+J�L�}�???����'OK�H�T�=i�������;~�_8���;�]�cń�w���W��^c(:�5<�%���:�J7��o	�r4���r�.+ټ��9 ��1���Ie8�@�Ľ��~�a���:}��`�]�N}W���\P4��@�H���LQ�Վ��(&�0�Df�xQ�� ʈU��<��2CU�Y4�OΧ ��V�Y4(�.uFķO��"�zq�W��2�F��}bI%�q�`�Гr<��?����n��[�F�+[�ڥ.���Nn�T"�кZM��4�o��4�����=��j'B�2RA�'��
FB�ȕ�Â�����E!�X����a�~�R��ӽ&f,�?}��py]K�J���[N��Ɠ�y�!@S,�4�6�u����:bߑϋR����rǯ�|�V��D��>_`%��)p��=�N9��������[�{&����e�d\�b�D@\I�H�4p�-��C`�a�k6���w��� tʇ�Ѹ��� @�	(�+�m��}Ex��
��x>�t���˗�ό� ��͇�J_�ր�EFc1
�r��#�|�fM:��~��$Z��?���_<�n��+E��S���
�!)7�,E��}�}�:�H�xb�
���!�*'��y	4��q=0����TnL��p8�D���Z�����қ�����Y�UT���e�,�'ŚO�5��>1 ���6�@Z�ɛ�o	#��sn��Oɾ(WO�R)a�Qeݎ��R����ˣ�NG� n����V�շ����Ё��i�q���N���ܺ#�f��rЊ"����N���$vh�H��V���qmp�@0%�Hc���	翕�H5����sL�mp:C��� �<�yj����ia����p�eB��]T�>�7/��̅\�L'�C�̦2�����lp�_^/O�nIV�Bs����l$�<��ٙL�]�����5�Qk��q����)̬��7����a�W21d��RK�|�G�v�#KF-���z{{��mF���q�����BOb�G�};˶�cfMU���WL�F���������kR�����tD�")�B@���QX��]�s9�=j�ѓ|�2 �RAtJ���R�#��)�# �T�H�)4�0�RS
r�dbH�~��˟>�]�}y��ʏ�K<)���;��0F�7��?�ܚdk@���N(����_��5�;͸SY�|	�	+�شr���f��k��۟�r4�BxvxLpW#e��R5���$٩N2���W	!ȼ{<�_I�?�����Y�c���}��γ0�ȞV���SG���GX����z�C.#F�D�!O	M��� z��CM����[O�wm����N�x8���諼���u��@]����'�b�cs\4�\t�Kp�]`������V�G�D�`�)��a�g43&�O$���W�����+�ʃ^�b�x��Β�-�U�b/O_Q ��:2��NT  �FT�B.\#�l��/���씗~��__�4����3>�iQ#��_M�GF62~��4�wS�U(9P�%��O¥�����c��D������uv�D2!�ᡡ����T)�i�(�HXt�	�.�.����j׺���X���d��w�S��}G�iߝ$i7��͏��_/E2d���m&q�HMg��	���譣����>���ۏ�馢��Z��B=V4�#�&��DC���A_��D��a#�S�V�!=h���Ood=	ϋŕ@�N}�tq��.?ݩ��h+j=��oeP���Ś|`�����P�48�&���7<�А�V�B.�rO�=p�JImX"Ԕ� _z���T�'�<���n�tϻ�V�1ֿd����[��fؤݲv�_pN��Kך����ׇY<�l]�}7)y��q�Q�I�6����Sx~��7,t����C�ČKQitk݁�k�j����g�N��pNA^��$����v~�&�}+��{�ϥ���!�Pb
xj��*r@��J�U���DmX�ɢ����1Q�<���_��E�a}��c8J�3+��rt6x���R��,����Z⢷���!:�(��Lxj_hɂo)�EQl��x ߟpؾ�b�[��"G�3�|7�{{qU[/���~H������ԙC�n�5��G���?��tѻ�q1zb(v>�!����'����u�� 5� eW�N�\�n}r���N��̮��c�Ѣh>c��|�zV|Am���7��(O�2�AY�* 2J�o�����e���v~�4[q ��W4$��A2��vh(Ќ��k^:|�����G��/Q=6D�9�B`�q���^�WE���l���H?;�� �����~�ތ���I��%t#���Q_�"i
�.�P��dt����]c��?.�GC��v
��`��+��i�E��WuǼE���z�hسXno�I}{����G�*B�W7w���ӡV <8=�����b�����~�2�빺���XMO�s{;X�^���4wHX$�J8QdA*ic��Y�h��,�G���/w�ЎS��9 o�5`ka)Q:�]lYF�L</�)���x�ף��%��)MI7v>*���1�B�-`�m�T���x�:_��4�R�<o!;E$BR�V�.y�gz�����ao���E&�_���f%�B&��v, R��*.��m�&�(z5��ah���(��!�X�ggG�燛�E�Q�W�u�cɇ�����+"�t�����fzæn7�7p�L�Ɋ|P���Q�E� @&�����BO	�6&9$����嘜\��_^�`D�x\R��(<*:RD�]#�(�0]�&>r ��8<�2���<��1"���H8�85=܋Ѭ��Io<�Vh��NMc͎wJ��Qf0WQ6��
~�P�|�g�}�LT�c�
dn_�4��S�%�ћ�&�in4L;o�-Fa�����r7�>>�����;Y��%r�"k�h����*Q�r�K�o498==��
)C�ڠ\�����အٰiq��0�Y�!�>sZ
?Fh�1������c���c�'ޤ �rE��稑�	A�6�޸���teLa��Nɮ���=%�]Mn�D��$���ͮ����Bf��5�@ؖ'k�f+�$�J)yU��6 ����i�� ���@8r>?ݧ�R��9͐0�U�o����ǻ��"!��v�����8�`_ڵ��O��B.ę�#Z�U�ĭ���H�e��Y��g��h����-������g��$��z�'��    IDATdؑ`����0�g��~A���e���(ک�́8�"�g԰ 2�ѝ�J����K��4�8k�f�A4��F�%��dE�XQt�
y6)�������5�[�"Ã>o� ݇D��Ԣ�H�\�$��;U6xD���,�E�_D1�ݧ����T-s�ͺX}X���`�"t�[�.���
��Y�D�ɩ��&���	�(����MG�W��l������Qk0D\vʅ��^]��Z��o�?7�MB�b��b���I�hǊ �{����������Ο��}}�}{�(����k�vJ���<N�*O;�F�[��fq������i�?��):d�L���Uc�������~�+E��#�kt�B�
��Eb�����G��G�@	u��h�����\��'x�� `sQ��9�b� it����/��0������Wt�2��h 6�'��Ҟ��%��$�A���~zu7��݊U5w������At��T��:s|$��p�éo�]��/�D��$�����G��wz�D�	Ŋ�hoO;�(��Xs3�����v��HD c����WT;D��m%�\�BH�$¹��=�#/>g4
ˈG��OlF�{ �x�RXB��m��!sk1A��[?��l�֛���ޚ��9wQ�~5�9�Q1L&އW\�@2KD��y����{�L���ɐw��KT�%R
��̦ҮVS�Q_��悔3�xj�9�/������~$�i�-������T��{Un�8i�ʲ}�7�˛"ڸ5�j�hO�֪V���(���H�*��^�D�O��+����Gk�
��ByCHݤV~���B��B=��A�j�Sn�!_NMy��6כ,vlO���;�F��~qa~�>��s���e���<:�	���ݎ�F��O7�*�wy���
���f=�e��������B6��0�o+ipqc��k
7�7��ۇ;��n���(˟����z2�
��b��-���Y�pv>���q}����>����g~��o~|����t1��6��Z&&�&�G���C������b8~�bV� �Ԛ�O�OGJ���O�����a�]�q������/f��@�ku#�˦����yYN�k�m�6�Ӆ�k��ZA�����=!H	�R5(���V�Y�o3)`�#�G=�i�\c+�)/6;vʃ~�bi{���b�9�������A!³��r�y��Y�{�N��n��H�|���_��__^^r>��=����x��|���d$�o`F�^�]]]y�'��Y�|4��!t��/^��#uʰ���M�0�����q��~��_y�����z��%��|>@��+��q�oI�܋!2�A�BF����
tF�׈��v�����+����yO��SB�x�ٵc�Ì$a0� ���]X85vpp���"��e����D��)�Fl�R$l!ԡ��T���h�}�8Da�$��c�D����B�ċ?�HbE(�0V{����(�>��7V�B)l��i�E�c�U�4R���D�`����)�H��F/o��"{!*C�bU	'�M7�W���Å$
��I$�ą&��H��ⅪP�c��eȾ��_��y�����ݧ;m%�A
H'�K�H����AV��
��>�(18c+� �'�П����8[�^^\>�U���7�\�Y^`���Ǹ��7;И���)K3�wחw����e�ᔑXr^��:��Ƨ��a�^���삧��QME"����ծ7#[�ic�?>��ڳ
��j�] o�1���7������׵A�㸉'�Cu�t�����_���β �X�x��C�j�\ߕ�G�z��ϗ��;�Ƕ����������Hqm��=�4���t��*\�Y�s�J�4�Zn�30ao�L^��aZM���栧��v�0�C�]�80�>��������s��qr��]\\�����c$
t̛2���"����5���S��Lڍ^���^E5���=Y�X���Hyy_�y�t(*��6,�j���������e��<V���,:����^��Ak��ab�f���Э�`��8�	��E��&��E]E��C*I���V�����:�jb'�R�A��8G�,���x���T�)�3#5�d="���Ҕ�𧧕
@]�Mc��ds{CfCB�Mܫ��*�;u�߄l����*GF�A�_/�.�Kh�XQ���T�z<��O'�.�R9>�梣�V������h��#�[PS�&�k��&�9�S�005Q������l��Ǉ#DE]����~��وB���DSKR'��[w��ɁG�J����p2�j��&��c��w��5V�n��X֘�A.��BU!�#�G!�,/>�o>\��n���O�BHݧ$j������n��~|��Ծ�k6�&|,�s�d�������~f[��v?~��^Zn�^��Э���҉x�xK75	�ḵ�x��lr}}��T�#H�+T�����O�����E�5#	�ax~H6	3Se,Գ��1u_=�d�����ʲ�o3��1�jw�%�r���.A�U��n�%@
�,g8�}��|��������W��|�"OD�x�so�Kv'�WKײ/Z-�Ca昢�o31�ii��\�t����i�SX�ª���"SD�֛mV������������w��2��C6��� S$*�)@�it�X�X	�T�LB�&�q��穮��2�s�<K��$�S�4�*���l�x�p�XY�'L4X=�v��l���%+G�3�H�HL���;t��PE�C�S��Ulml�bf�@��\���͟��*��l�ǽ��Ӗx��������Y��S4������7�Xf���䘲��+���^���w�)9�ǲ�j"_�ӐB��tо0�t�c\C��W/?~��n�XJ%�H�Lp��$s������I�U5Wd�p�� c�S7���h��Mɧ�V�9�����݁E���c����d��I��{%�޼�k@�����~���Rn��3m�F����=�dG�_��Oݧ��&�$JNnX��������)����a)E4c��D�g�8R�D��F:�?������H���kڅ��枫��/.��$6�����<I�����D7n�zG�c.��׺#�N._=]���Y�ŝ�5������8�Y�?�}-��;�0�K�4$��L��k��a�g��`beZ���6����U(� ؽL��h�B��$4Y����r��x�� �X�,S!p(.����b;]�5����C:��8�}pO3f\���Q�{-��c���@]�$k�1i���[���T��ɘ�ʟ�h��R�����V[��λoo���XRӠyw��Y�O/D�"�Zo�MN&���e�O>���µ��t�B��R$�4�����o��09{�v␭]�?� M�o�2��r����=��d�G�����Rp�ZZ�),��ٟ�a%�tyk��V"x��Y�z|1��'����V��#�pG�盋cK�n1¢�V�9�"��v�����v�̬�;�G=��ʆ�F��쟄]]>?>Q�m8�Aaauedbl��[��{g�O����q겞�V�V׌n������Xe��ɸ}���G�����UC��wX�+|J��B�ds�`Ż��rL�L<pvd��)��4��T ;��rh�%�6`��+�r���`�|��&Ī���B�D�����t�M1�M�a>���|{'��کi9Pcz|��ǳ���%�z��tx�3G�V�:��Ǻ��HH�MVl})�B=7IE�ˋ���Z�]]ߋ�o���ZN�\F@��I�8����8DQѐhs�	P�7#�h��_L4WX4V���*��3(��
,�NlC�J ���S������>���c�T�Ig,\ YP7��e˱�e����y/D�6�d�mR3Zq�.�qM)<95Q"i|��7
�'����*�b������Dd���I&���H%��ÙO�r�t��3dz���}`���pSwg�z�N��n��_���7���H@���!i?�-�M�咫ԧ����iJG4'��I������7����b�!��G{�`]�Y�(��䭨�ẓ�	W����K�Y�+<�(	a�BFf��+0w�4 !����[��y
h#�(��`\L?q?<��r-��*����_0#	��c@vg��%���:��O׍��x��9}B���huL��� ��2\LF~xT���S�k�~)/fO�I����G*�I��=�SDT�乥���J��@Oz-;w�W®�^�.�?��p1m;���]�謥�H�,7�� 1��,�BL[8x$<!�Vm{8qJ%�L �'5�b���/p����g6ur��ft6�e @���1Y��.��ƶ �a��A��
 ���X�eCi,���9��x�6�!�YW�ZXGކ����Wg]��_�BYn�Yt(�l�δ�)WM&������w7W��slG�`w	����9C�Kp��y �$��Ž'�sc����CӖk�G}p�KVY_.|C�"�ʅ@�<j�>ę�m�' I�>;��
r��y;��M۰���\{�?��v��d`U���rIN��9ď�?�� |Q-��5B]E*`�&�[4~�=R���|y�n�z���ėioa��
�F?:���[xb���]����E�?� �J{``�X{a�<�]*�h
��#�wϮ��'�~��U�w��)/�FS� ��Z��	Z=����N�4���e�?�&FR�)�Y��Y�7���j�;�U�ݠ|1��CeôL�	<�k�	 �����\n\�J��qi��B�;І��+���9��Y���-q���$��b����ؘ����Y_����5�YB��'�Vx�X��ylW�(���G2��&ª��V��~�J��?�E�z��,�`,���R��l_�",����9������Z�I�$D�\��fO���08���bA�=!
&J��_�8��z�p�ߊ��v?~�z�x��\��	�Qpǭ�©-FD_�Г��G�Rj[��yz��e4%��Cf���H@w?���^zv�r���><����D��1꟞�"	G���Q����۝"�>��� ?���Sf����'����x<�p5�����ߛ$���(+������o��oO��<	+�+b&�H��(w�4*�i�j��Ht�#Kp����<��]�r���5�_
����c�*�)2���c���"a�{��o�I���g�P�_��3���򂓄�W�`�=��T��6�*������'���y:0��%z+Q���)��Ӑ�a?r-&v(ޔ�L;��<N��k/"+����Y|�\>�Ӹ5�J�I�o���y���5��2E90�PTS�D@`����0m��g��*IBu	���Ls+�RK�+�l�0��+�=�*�P��v������9�b�Z"�?qd�DV�
�� G��G�yIuul@u�v�W�}WKS��&.�n�ۜ3�B�8�>F:�S~D���KH�~��[�c������fn�� >~r7�����T�ɱ� +H�΋�Aj	��` ~Y�>�� �̪"k-�-H���0�+��?q�=���z]������8{��7�_?�U6�C�#Y]���û��r�E8<��T.f�����W�=��&_}u��r��� �&���k�������g����[��
��ul!
##lK��"qۉv-G#я�')ʱyl�eJ��hwl%KPB'Bh��W~ �w�C�I��x%}W0���
��o�F �F�`�o�.w[?Y�qg�q�&eHVǯ��ǁ���4_��m�I��@��'��7�|#��HWy���n���0�x�O>�ĒI�4��۷�4x�a|��W�����?���~��?��O.�q+�:���dM�%7�_��_�]_|�������Sr���?��}���xD9KM���?��t���ti��޽�b��t�ǃ+���9�f�د�9�ʕ�tNt0�%!��%y�T�F�{�X]��n���A������=)]�K�N�+�_�?;�����!����Z`�dy�������m�ܓ�$_sv�k�*�xF��XS�9L-#P��%�Sr+���mi#"���v�#�e\Rs7���#���4d3M�<-Vop���w�B�&���iR��vj?,R�0�� f	�0ĆyJh9���e_�HZ1��V�J���۰/���y���Dn��%��E���l3�(��n>ܰg�nW;}�~���	�q�{+��ƀ�P(w����� �U�0�,q��Lv��9�L𡠐�>���\���`���D��)�3Bo)��¼lي��bW����	X���K����[���%�vl��e"h ��zq�G�uZ/�����%�?�c�i�B����	ھ��II[Fy��w�;r�������.�����fH�F>Dȫ�[��"�@�}�����o���_?6��s��6�$C�vzzz�>N�ݫ�b|=�9�Ǿ�X�0�P�I�.Ȟ �'�W7��b ��=
9*�,ޝ�PA��7?�P��`+��tw �Ks� �!���#�%�{m7���yX�������Eh�yW�U��?��ڻ�V �P.�}�Zz|��L^#u�ܝ�7�=�$Sv��/!0�vI�j�_^>���9̖N�Q�Y�X������!�J}�sfj��Z��i�b�E.��j !�3�i.V�֨������~|��}�!zY��`�i%`[�0��Z���ٽ$����:���\�����������D	)BUt�l�(�� l-|,2�Y�����d�����8��	>�{[M6w@	m�4�v���ŧ�/{���������.U��g?b�
��_�x&���;3��%UY�i;�:���������3^��iW_/I��_�����/��v�~����û�[:U�K���ͬ�8E0��G�3J�~����1GeOH,����)�嶮���&P��~7�Y/:Zښ*A�O@�vP��Ƌ��1��<B��e	�`c<�Ia	�S
�#Y�	8���d0iO�N�s��Y�S��D��fu�I�=�L����Y�|ݧ�_��+� Z��<1(Tk۾�eR�,Kl�}2�"R�0Fz��
�M9��〲��]���S�O��f1��Ji��n�Rp�1o?�ܑ��Q)�׮gk���㓳O�I3�5_�_};��n��	w B؈{��N�
1� �S6�U�n9���Qh�w��I�{2~�	��H�B�w@��&����?��
zY��lr�r�E���s�PZ�$�I�"y���u�w���_�Sm��7���>����2hp������C���I��1Y���>}ٕ��֭a+C�m���&��.OT�/onoW�s��T�{�Y5����O��#�l�A�%�K� �99�I���󟟏���������=f����$�I�/������*ck��˙�;��|��2���xB[�M�p>�_����h剎�ಸ�Ba ~�jY�� �5-�wjg&߳Er�j�,��'���9}��?{q���]�ЗX��mz�I�$�7�!���n�;���ݡ~ǔH���I}@�m�n��}��s:�i}��yt~~<:??���C#���~1߬�C�љO�同|V��t2D@G��B��a�3�|9�����O��jA"��N�\�������]G�ۃH���ջ�f�*��q�l�D~�
&g�"�G�$���3}2�m$��H)E�S�I��i2�xx2�Y�Sp��L�.��)�V*c4$;�S�I�+��A�.��t���a!a�[��"��h�$�.@")�F�]�""sp���"r<�(�xkM$�
]��L�uݤ���8�}�}�8SU�$��������|��k��)��6���Q7��R�tV}�.pku�Ox�_|$���cH��CD�ϫ7��e��џY�B��r���J���o��l�"a��	l$nß6o��n<_7��BĂ��C�^�����ϣcXqԷO�>Ag�����CU!7i%�
�	�j�>P��Ad����Bl"?��]S=�)��^�ꫵ&	A    IDAT+���%�@?��g��P�Gh���-v��]H\ITY?��u������K�$$�5���9?}~�B�m1��jFf�$VLoDP��G�i�og�.Q�c��86�[:i�΁�%��,�L�
���0H�>��p�(�Dh`�� �6�P{���^�#'��J��p�2
��0a����a���vO&S�:YϦ31�,N2�S��Wǻ7Ld�
~,�ѵ�;���P�.�/^�u"ڋ�I��mu��s��LS�e
���9�&J�ٜ=B8º��
�\X�0��=��ƾx��/>�_���_�Moo�X�@��� �%	�}�L޷�i�$��J�����b|�������q�3)��4祗	�a"��}1%��G1�CD�"Tb( t:���%F�p��P8�Aj}s��k
�ח٩V��Otg��a��.�>�s�4�o��l�l�3퓑09�T�Ϟ�ON������Rp�iGJ.�J��}b �\	RZ��f��^��cJˍn�������پ]��)�g!�k�;��E�M1�j�-��|FxZUM'�g�F�J˪�N#�� ��Z�y0�ħ��jT+��yD�o'��H�ׇm�:�������Eo4d�7���z߅hCՠ�Uїa���Ψ6>�ٯ�������n!8G�y�I�if]։XӸ�������'��3XG��΋��޳�:�L4�>�٘�V��>�V�`�Ե����/T��z���!F��Cu��-����f��K!L������_�tO�?�&/$�*Um�6�M���8胰��
��6���/V�m�+��bs����/�-�!s�-j����c!�s"�E�6�x&�#�o_��0��+� �zI9bEM9�����0��?Lu\e1J�m����[X~�tYk웘:Zo�iZ|�:�j�U����UP���㇫[�f�h�p�V���0eK�d�d��A-���G�FZ�/�!���
� �a�)�<�DԦ�y<d�S"V'��{;�A�Re�"E7�z��kg������`��![!H�`⌵pP�P w\ �Rpz�G#u��tx��{@c���3���ōU}�0���Ƴ��ry�C0��<ܝV+�ւ�(�07%Xp��RN�[�j�*���M��P�}@FD�L�R���!�X���n5�0�u�PёUR�&,*=	!J"B�o�"^�I��fo�ѧ�Gr�?��q�{8�U�g����@��E��ܘ�"q��׭J��$	� ¥; �e4X�I�QEO�{�c�%\�a�"����t��kikn�#���DVd�G����T��җچIh�������WD��GF;$��T�n骾Nȡ]Y���k�v��WB��������s���'G]��D��ՊAE�}pp�v7&�VwW�,~�7���,l[����z5VQ�����k�nbaJ9��\ ��[\D`b9��17���+�'@����n��P��UsP��� s�oyJ��.E�b�*��
���H�d<֒�Z�V
L�Cfp����"b]����W�GK��$�����$о�ERW����`!]RkX�����O���~>y�5��|���͉P ׇ��KE8��܂�	�f2�QN���Ѧ�� fv���'Ң�����^}��}�����_�ٴ�-V`V;
23A�J)b�����IU��PL�(I�=`	l�����+zbE*�;i�*P����4���dd֖�!k�C����/f��g���Rϣ�g�(2Y�6����3�V^�ʱ,�Ln�����{����p}����j���['C7i�B��f����lJ��J$[b�7G�ztj�ǣ�L)�����qi<�Q��CD�JJ�l~���F�
8R����ttαr�b���M-S��as^ ���X�>�5�����R��d��V�_F�6���/��� ȎA؁o;�����Y�ܷ1T�nu��|&X>����ӟ��}[�2�X�������p�bF�֙��7���C�,߮u�a�`�q�z�j���YM�F7/�X�>��Twr=��X�T�H=�%,x����	h�@F.d��!�=	���^����]���G�?���p�o����5+Q��Í�~��0���K�bX��/߾�)ʵ[�m�C[������W����_�;
���.��/�G��AZ�d��<��k�
��I����wY��������"Hx�1 �f��2�xy+��Fl��٢���q��F����ժ��iWkd�;�%��Tw��tm�����]��;��
f��F�؁;�~l孬�ı�u�բ�	����12��}sR�*>�O��1���yFϭ~���6y�Hcn�����܅G�������yn������$�Ep7��ǤU�V�������z���/ܔC�U�$xh��[U�s`���g������U�6�	c�'��{Ϧ������X��|x�V>�"��}�;�s�=�-�zS�
�N:�f���ӭ�_��]O�!������`���.m��G>P��<��é��:���i���
2}xr�,�w�%L�3�5�AKac��6�@A0�b�D����v̞��7�@�dPەtH=&* ��1�����_6�2cuO���J~1É.��`��&ݛu�012���	�i{nn֦T���Z/*���Y YV��&?�0{���Tڿ��"��\޽�H�	[��,���T�m��շ��̯�ˬ�够��]��E5������9��{���1����[��%N�T�ʯ.�]�ߛ:S=�6sO�����?{qyy�i4F��%N���(���a��_I/'�ܨ�M<o��r�=���pc�Dp#L��
@�%w�Ș�7^"�NO�/N�I����d����÷�Mj҇�3��7���/^�p�#���uS�����V6��b�B>,_}���F�����v�"Kq+D��E��Nx=/n��B�-n&
n1��!&�%�b��PA�Z�T4�* >��{¶�@�i���p�Pb6�z�����c
�g?��l���4��dt�J!ZY��fo�J��a�}l���9���P	�LM��������uv��BҬ�6`ZH�/�.t8Ѹ��Xk?����Pz'[���@zu���!!�>�e�ő-��"�U(�8���xxU9?�7�|j;!q�$�ۆ�h�ݔ>$Ϻ�]H܆zz�����Qy\J�&��:*(U<(P�����s�Fh�Od����E�Y
�F��#�B{�pA<u�<�$p��Lc����G���y��
�3��B��ס��RɎ�&�B+�=
x|4Tv��tfM�O�Bp��E���ei�vz�6�6�6�*�'!��?��=��~c8�1U�̳ѵj��_�8ʼo�Q&�=-�@��������6��~�]�j-�L�i��^�g> ��������K�*��M��&�1c�rR
 b�12�Y�;~�E�t��E�"�s	X��H�Q���/�us���b���|ڒ�F�kD�Fپ���0�	�W�Q�?s��i�$l���c����`H�1k���PgRvZM������A㣕�jڤ�V��d|��SMt��z����_���z��8�Ed�8NT�^9�<��O��0j�%q�!|�Y��� ���6�����,v�p�r3doA�CU�_��	/ޮP <ؾW�N؎��^k���ꪬ.��m3�'�
�)�6"N��Y)�"�*��3!�G�?�������F{��1j[JR(�c=�$y�Ɇ��#��NO��y/��Qw��5���8���s�i��v"�o_�M�h��ޒ޺X��pc#2�%A�O�#�5�����
���X�9@o�[XɥY_<t���#<iY���n�b-���1C���}r��)xѝl�J�K}��p�
yw�>���Ň�p0V�T/����K[��9I�H�b�#�ZLT���6�R  �z)hCK�^ħ,Gd6�P��Lf>{0x�����G�,�Dj���d$"�C��OL �w`8�R�]���d!:��*��i�ƨ�.�������n�K�U$&Z�ˤP,�äb�>>�<�k�T_O.j6�����%PjPIy������}�O71kֻ��8}H�aoIk_[m���Q�zw�@I����zB�����o���(��̍ks�>r6BxK��OD�y/�<9Q �Y-�Gu��֔%��DR��+�V�h��j7[��Z;+�(j)��(e�����jJ��AT�t<��=Tݏ���F�JU�T�@+tSO��
I����������9�*�⠋?���w��7�&��>�x����퇩)w��NRX�,J���h�t�E��)�ߕx0a2���3e�9:y��sq�"�؉B�AR(��S	j�XvJ��6$���f1g ۄ���Ζ��p���Bs��P!}#v��Ё� �cQH����{:&��d��T�]�}�S��[[+ؑu'?'D(bjL��9"�J��j}��x݅*��H2N�b��"{sX-�aY��U�s��!V�$�f;;z1<]�4��}��YeH���0=5��l�"S-�����RA�Ƃ�7)s7 �F�P�DF�%wKW���5�(�@5z�K=�GX�dZ�M�\"�4�V�E	Uw'��A��:x�k�u8D���4����K���k'M̫]P�E���2�qreG�����7�����.�ddS��:wT+t�u����6fE��l���$6��D��"H!충�n�Yږn�8��#�_w�f�R�V�r����NߵCo� x{|9x��D��w_\O�k��A�f��Lo���Y�mC'���r��.�q��P��]�}2������֛9���<2�|j�D�f;�.$q�,�R<�>�X��U�ܜql�o?A6�p �V;_�tUu�\�lǖڞK���wo'��ѪvW ��ncr	W��2,�����H��N�_�Ɲ(�ܨ�+��?֛a4�LdK4��n�pW*�>z����X\q{��3�x݇'Q�p�gl*̓�Q-�gm����l��L�z���#G�7�u�R��$.?�Z���	YP�U%N�����=��r�x|H"���{�t���z�����C�F+"t#0YI/�ʢ���&b$�Ǵ�\
ۂ�uw��]f!+f&�0h0в��CE3��b��UA�q��,�G�3�Ay�ib��8�N��W�r���X�Vs.Z.�i�q�R!�*%�f��������KB�j�
9ȇ_J��%��4]�3Jl��i�ɩç�8&��C$�ۂI���A���=n|���+5�����K�ؘ�S&��V�rņ��O����(8�L���xb[�WE�O15����&�G����� �bׂ�9N��X��rV�܈f#�Va�'J�
��ޕ�A$>^s�(�@�e� @���6�.Fg'qq5�j����MJ�'�D��CGڈx��#n��2��NVl��4Z{k��~�����iCT���M$�DOQ�k�U��T�2+ӳ�0:鑴�����ڏd7�I��t���O��	����j�FúTy��A�Ǭ�QA%(�ӕL�w�����V��|Ny �#�p�O@�sA�Z�k:��L^��y&BC�o��|S+ϰ�pL�2x
�c�l��_�����5����o~6���M�u��)��^Sd!��E8�,�\�Az��.�B�L�6��\W��Qd|�W^\@ͼ�$��1��C5���n�+X
�Z����t�\I�NĢ�.Q�����W�|���X��?[qL��-nfNM\KU�����wL��5�_\6����k�.�܈��2�p���4`!<�J�S�6���D���BI%�:/��$�Q<n��B��wVw�K
��/yq1�5a��,��T�Z	�d����aF��h��T� l�C�Q� ��C�Fц|0)NJل���6���QW�Գhr�Ŋ�q��(��G(@�}SVYޏ�~4
��$�?�.�B(��z�N��ڤ�jS��1�r�A�ȿ5;{�� �6֊�5�a�icH:!���Ȣ3�AI�6" 	��$"'�` �� � ��W ��#&�ep�B��8��G�^'�
:L6�'��X8Y�<�'�6���C����OEP���i��¨CW;�[ugbɣv��qɠ[��$]��}��K��� ��������ptz1��� f�G1D��>d�Ճ�}��MW�خt����Dt��ئx��%��m������u���/&/�f߿�R�!��	`�f��N��|?}u��F���Cm�u*zC�\	'`Ԡ�
%� ��Fs�e!d³~T+�;Bx����5��k������궅�Y�Ɖ����ϤK�0�������u(��u��g�I��L�ך�����c^X��Js�2���f-��_w ũ������^�L:���-��V� �T� obA�C!9�͞�^�C�}O�T"�=�
?�Jar2���6Ad^I� �;��G4�bm��r�f��HBP}rg��1bw1�����������IKPA�1$:�ul���G��a~�:�}�j#�x/�a�=�t��Mܭ:�]-��~ U��=��V��4?�θ�a>������<��YUV��+�$}�vy!xb�Y.v$��=[��f�[Ζzc�@*@��'*�������rp�0���Y\\	ںӚ�������B#��iF�����q%u���������������ڵ/����9��8>>����La����ۯ���9_��2)��%�O�!��Di(-uu�Ӑ����Yu���y�g��H`�`���:��F�E��!D��DhЏ�3*��@s&�:��T��H�'g������_��3~��v�����J
���<'�w��R�Lr&�/%F~��7v���!�\k���gq��~5����7&�]�\��(��F��ۿ�[��ʫ9��t[7����/~�S��߶�����m���3�r���S}�4c��lw�'��{�����߀�_�����UM��� ��W���~�P�K<B�A:ŋ��^���Q���0s�
��]����g�����CM)�so���1��u�3��T#�1@���,l@ŸW�`^�LBK��YH�H��+����6��[mn���\eD�)뤲L륿�k��)�"��E�Ӓ7�4� O�ē@be�E���mZ��|���&W�)����B��r Lu���Ƙ3�(���*,�TMb*(H� �%��9����צ��`bb~��Vp�[�Mme����Dp�f���^m�/�-X���;�BO��쇬��8���^�T6����Pӭ�?N�[`U�c�`�L|g����Zwp�z�_����������+�]��� $������p����*�	�C��*w�����G`���Z:[��(������y<���k}�[�]�p�������X[.�񸬦V$�~#�� �XSW��-}8�Ld���q���g��lO9��iFݭcm	Z])���>KC���?�f�v1�,����p�7����������a�ၑA҃ i�e��2Q�<���^n|*�%�ɠ�LWUq��,� O��j���U��l*�$0E ��Df�/�J=:}�,�X��4�yC��}�܄
����G�N_��e)X`�M^���JABE�~�ޟ Ρ3�m��\gHJ�H�`��"a-��� Bl"��ݧ��.X�p�$��8�;f���.4�j!�W/ih�U%v��dƲ�Y&�i���git�jbH���<���Z��r~s{w�}+y��9�X�C���r������C���7�Q��oJ�ɑW������V�B�k*��-�������Z8 yKt�:L��6}\I1�����Cɠ�"1�fO	@�	I�E! QDCI��J�8ZGo!��4���OE��fc�6��Y~0���� �ݔ}C=���F룐��A�~5��/w1 ���}��~��W�F���~��MJ�Z��kf��G�^k?�x酹ʟ�W˻��ۄҶ)��\�ky�`8})���/��x�uBGb�� ;c��(َ]�4!*wRҭ��D�
��L�� A|{�:���5�$�߽����h}�01N�$�,E��bJ��DHA4�k
*�G��:(�ȵ���j�V�n�.�@�'����y�����    IDATj����˗�b��^�tz �?)w4L#4:dZ�Q��t��m���|���$U_+���]����:
w�ql�����������j���o��v��� ��Bv���M-@��i����yu	�QR�t7I�b��A�i�6�	��$�! �n1�U"([��5p�|��Y ���7�+3��Y"G�r� ��n�$����op�'5k�?��i�'=y,�N���]��򙒂7���E\y�e�y�R�q��v))���RrG�`I0%��'Gǻ�F���{4���P�?�k׳��m|��?�����`�OTfkz���h����c��ů���SK����=��E4��+Ί��N �Ɔ+�Էs��SUfF\�Z�E��$� ��&�,�A�)�78�<�
���̡����>>�3���FoS�ߦ� e��&5�ep�\葀'I#�p��ί�����/���������b߾;4�7�G�h�w�B���jb$�׾d�	1SqA�l�y�ak4�RAd:��]�Ҵ<บӰ��;�t`���� [;,�+��Z��Ĩ����}�8��X&����R�'�?�.�5�OK&Hn�o��X�}Ɇ��������(j��`,S �U`�x\��كJK�@3�j���i�_k�3���+�Y���`j�Vڵ1ڮ�3H�8t=���ےB!�Oysu�S��s㞞���X��j��aJN��/>�D�q<k�,�������b}ܪ~�G��ɥn3�'U�"�4rw�A��艶d9J�)/]�3�ێ'c�&��]�^�Q�8�"Ys���ѳK> P&�/A�J�����Bbn�p��>���W�֖w����E�>�]0a�!���P����i �e�ng490P*ZL!������)gP�GkH�������~�XM�>D�,��� Q�n\�I�Z Gtk[<�����R��Ȇ��-�@����hXB{�;[)z�R��+[xGCV�3����/����X�TV�&B����ׄ���=%Wk�����W�v��n�`l���d����^�����n��)��U� �M��P�$গ�Q���AvL�0[�����ppO��
`*���	�(�p�zn��B�c|�e�lF 
B�/�9�ĭҀN�J����p9��F�(*�0#v�.�+����r���C�;=Eũ2]-5-������;<��u�#����ӌWy�����뇻��xA�[<rR6���=�u|��[�f�Tf����J�%&��h�?��)�AxR����HR@�w��f��&�����r��~�hz`��ż�d���=<<@Nf� }�x:L3U��R�w��r��[� ��
���@���h|��(S�nsw�^Q_1�S%E��������6J�FW�m�t�����~�U�LuF9���cO{�%19�:�H�)o�`E|���ʐ&�0iC ���-<z)b�#�E!g�ԳM�X]'$H�E�bg�!aO��H�$H �$����BX�[�+2m s^��� `/�4�߫dG�ۃ��i@%�Vy֔�8�!�3����jǯ�d�>�O������DkN�V�U���Pr��(�����������Ƭof'��ݸ�N*xq\&������֒Y[�=9��f�N�1�3��+����������k��5�lؑ^I�����[*�+.l#%�ON��_�x������-���ض��O��#Lq����
`:�'�K���"�ɼ%�1%��ܶ�׻���멥���9�ߪR�5��g��L%bؐF�J��?<���!}��`(���I6d��VU,�DA��$���&�q*�U�/8�Sjg�-%&L\����nͭ��ƫR�	p� q�m��6������ ���^�8�:�P}4z.F��C�%��>>,��G�
�Q/��������/I��4�2��a׋7/����^�W��&���犠v�����tg�(���O&�\|�1 �5�7l��X3ğ�c	��$�2AQ	>p�� n�b�Rk^�Q�d�.rB�Z���C37 �#A���mE|
�s�}"0�sD-|�-&iQ)_:6crI\>�ffI��*�P,5�������������#'5���Qo��C�A���y���؉?ns�w���	�l�r֧�+S�t����w�Zݞ�����9�(� �VT��R5~���iU��Fgj�NUo����ؗJRڔ���`b��jxy��+,�"A�����ZP|�Pb\b��.?@#��n{�;�u�P3ɯ\hvob��gM�ޖ�-�6���������kgXÔ�"v�H��sjԇL��|z>��8��h�/��S���ĲeV�T���!�4&���Z��$��6c�n1�v�<�������/u�%`)��LQ�T����#8�� ��W3x6�S+c��]���~�=4�������s8�ϊE ����|Ⓖ���'$�!�#?�[��C=�
`�ѯ0�`i(9K~U�f���͇��o�F���m���lz���Z �#�Pv�r��U�[a{��������XaOO`��X���V˝t�̨A��+y!v��9J����c��E��%_~�V���~+L|=9?;'A�T�'^L�8lsr��t�,��hۮ?.Ĵi�7�>���[�������L"�i$p��[�ٞōHBmH�j����4��=K����-hS�:�*P,AF�nX�d�̝�\ebxχ*
��-r�im���JRJ$Be�d�H�p�O������/?��_=���g���xxV���Pjm�0%��3I�T&��a ��;�C		���x����'�#�ŕ|��Ja�����aKS�[� ֬���7�o�^��4Wۅ��,%(��>=>��_��ί��;Fژ�G�A�y�hHw\�Lh��P�8�&��M�n���lS���"�BH����@|���s:i��@��H�U�yu�0�_]�����T���O�k��L
�v'��n8v�O?ݭ:i���_�iWw��O��0յ���c?����g�F��5Pv��8uC/\]fIbj�M�}e���+��3ۋ�=�?�r���`�f� �|�P��frۣ�����H������l�U�B\"��&Y���K|v�H#����Y�h����C�NtZ��\X��9=�
����ySU8[��ZL�rRE���ȲWltc����5-NJd�K���ݓ���`�O�2M@j0�p|T w�����9F�����ꠂ�cü��ޭ`�?};���6kQ����͛$��GR�����%�8pޜ}��������-��o#���͞���{�YrC��䯉�ⷿ����7~�,����.sR��~�J^�˸�|�編�ǟ^�U�ݱr�V�3�2<3s\˷?+%�U��L�d�8����";m��0��J�B��ѩJXNG�R�P�N�*v��I�\䴜,S�M�ăܓ	�-��S:��6&@��0hyxu��R�q����[�@�Ԕ�bc�.I�I?xJM!�I��lDJ��S���35�0�C�ȡ�[����2��f�/	g�P��5�H����3vԄ,�'dBb���Y���f ��V���"�ż�P�+Bq�0�wJ�J�ؐY
�z����N\��*�_�G���^ث����������[yT��sY,ڿ�ԉy����8�M��'��jS��rW�˱�>�W�m|2����S�1�L�����?nU��@L�,/�ۺC�1ޣ�|��s!�?=�ܪa�%�؊�]jcT`6��� ʰǉЫ��D�t9���w�X,a�����0m[S]���-�2�A�Jf�h��ѾmXq
x��u�ѧ�9._�Ň����/^V���L"���g��T���
v�&���w_ys�a�N��?�=�	1t�e�,nǯ�띫����;� �,O���l� qMͼ�a,V��btJ?�1��	4~X��兺�[�(���lE�i��b$��V��_�*�`D�k���O>���_��~�@�l:�b-��	��' eBWx7�e�<+ۑ�w}}�}�}�]��|����6�i�1�V��m���*جQ�]�MlAg�|��x8x��Rl0����APy�Ш���=yu7k�����4�"�ں�?����8�|v$V`�rd��)ͥ�0@~�v�h�R�}L��sk��;�*�kD���Y�-~b��k���z�.V�sE[�C���b!!�x��w����D�Wn'�����%��>���0�l�R����\�P�r%J���QQ�X����.8'�+�LbS�k��j]c-x��wi��l�`��Bd���N8��g�Fqm���;�ź�g���x�UӢVj+��U�O�D���P�ӓ>�}�]�S�
�HZ"{2��5�^��GG^��Z�����v�x�:��^�W)��!Ҭ���� vz�3���s��o�%�����䒰�rE�,Zo�y�(�S��v+o�SRV�A�4�n*5GVfri��7���\\����.w'w��$JI'x 2��&����y��.�R�dRv�j2����QkI��Q��ॶ���O��D:�A�E��OV������w��*��O���`E�.�Ű��[����3lu++N��h(2g0:��Ә1�F�M�q���g�=�3yq��5jV�W��ۺ�kJ�Ϣ"��+�3��[��a��eO����O��]�����[o6�悡�/�� �"��5����� �?� :�9	�S|ssu��u�7�eƨ~�N����Ľ�%&�?��znُ�l�v)��Q!<��N3�������ό;����vo޼���1$uo�ۛͽ����#�w�8�[�^I�g;`پ�.��=�Mń���y����w⢲Lj�����~�v	*Q�(�z��R��}���>�d?+�r19�=�]V�er�-�&d:��ƒ�+���DHK�E���o�j���pP��%V=j�]��Y�t5��Qޭ&�5;'���6��~v�����y��۹��G�m�b!]{6)T�� �q�P�����H�e���\�Z����*��뚲��W�JԌ
�����E�L��N�[�T���b��tE��R��;Z-�ǯN���n�����qҴ by�̅z�0S��������z�11�>n����Ŧ`	��~8"Q�[rs�Al�� �8�)ŕ�[ܭlb�|��͔��1�ݼ���.ڗi<���WDXO.��PK��hjUe�갤>��p0�F�8h�IN-~T$m��۞� EcU���q9�k��0��`��*��NH��8nw�_ߋrB̮�^���\��=�B4HQ~�pp���h��I��]Y��W�IJBy~~&j�pS�7�F%CEE@0�V���0��%��q[��{i�E��Ё��c.L��袵����'�;��bT��*� �c\H��Ad���B!^���Rba�@��۲�0�����a)���&5�H-R4"�}�i)��BL}Ƴ��5y4�l�fw�O��;�z���kv-SsN��yǓṤ�vc1U�Q�JF�2zJ��!P_��z�a6�����*�ě¶���O��ɇ���O��Z���L��y;;|N�튣X�X���+���D//nN�g�07�+�n�e��!�g �} ݊bXk��vO^�~2�I~W'���&G�8<L��_�����E�p���c
+/i���jL�������A,�*.��l	�]���K	�bBI������\��c{Խ���~yF�U������ċ��o���]ǣ�ꉧxM/@KDooԘ��Fu �mj����$"���H���v=1bpٴ\y&xST�)�[^xYa����S˽5���VeC�� ��1Ư���� *�^N�?s��%|��P���&؂X.��o;Bm���/44���/�2*#�������O?��7�p+�I�����*�(("v&�d�e���˂�x�YD^�\I�M!)=ù����lO���'gLi�������(�&�G��Z	��Wu�w����+�Q2�O_�)0��T�9�L)�c��K$.f����V�0�֬!�m��D��=�%��7�Y���\�`��R�H�_�N�՛�� R�)��_���2�}*���PU�\^G��*���DÚk�aX��ZrD�_���0������6zz:��Ԏ�;��]E�*Bă�U}QYI�6u�dw�=!r�5=�[�� ��!��\!���y��i���Vz��k��JĒ,�2b�U����8͓�
�������Ջ_�k������DW�����j�ʑX��o!�^�}�0TL��zs*�T���� Y�6D�짆��OVvNH��@�B?����d��⦘����Ja�����pK1��(FkJa�+q=^ϰj��>���_"o�=� �i� %�T��0X,�j�ۺ#��(�p�nk��*b���L�L&b}��	2��%�+�qu{����p�;�X7��Ȅ�U����j����Gty�)��Ǩ���(n:�ϐS�{�H�%{��_�s�Ě��J_D���(YV��{�ܶu�ި�v�����x�|z��>��u���	��B��(��r�V���I�Od~�GqO��D!q����|�nt�t8;@�%P��E����06y��j��P�{^�x��U�u��6�
���r4n^��;��{��фW���K�픻�%(��\��q7x��Ê'hN��XQ5��g�K����B�S��K}(�>������֋[�����^ߤ�A�/�eB����c/��MhLL�ؾ\���k��VT�$�$�M��E���:������œ����IU[��GX��Ug�N�`W�t�!�"�\)��j.�:��v"�6,1�uO�|e�bhE[�}�|rqv:�Z]/��#��d�W����"�]߉p��ӛ!�Պd�t>���"� ��Z����L�"�t4<��b�L�հX^��+���Vߜ�&���xI�!S�C��1QV��a=��G�g3Q3H�P���N�����	�n���xS�Qn�ۛ�8i�~A��3)'X�CM�7�v�[�񔵎��e�R��5h��o��zg8��zt����ӣ	M�ʠ랴��Kt�<<_�]�������/o�#�b��&oK�}x�LXCfr���9"~$~����t!�zP�L�:3>��qg�]�h�'�
8a+/<tDP����d��ǘ�c����ɤ����pP�⇟
�˘r �������# ��gu	I���;��AD�B�5Ǟ�5����q����mC��0��Etxt��wP�F5�������ѩ���?;���n�O����廛�;!��O`�F�r�p� N�T]�����m;��x��W��V}��廩t�t�?Ć,΄\O�
��=jx����������_u��*1��	��	I���	3���\q�y}0�+{K*$�S���2��ς�Cz�3��FSD��D����W���j�~Z�����(zR5�:p��W?YY�Y�H��8c@��l@Ш&`p����܌�\7w�������T�8�O5Ɓ3eb�8]��!�q��Ӹuٞ`;A�r7�h������I<�[Fg+�:Ier$��ѭZ��䢮���B�6�K�G�1]�62�(���q��&����Q��F&$I��!��t{-o٘�[%h`����
7����'j���i�@"!�g���Hn��?�n_�-�\M�?��`ª�T�������@d�_+���j-�4Ɵ�Y+�����3��������ǟ�_plѫa.���rw6�/^`�Nz��a���r�j�n^���h@U�����+��� �2�"rP������_ ȷ���6��.���/�0޴[Ϟ=��ng*F�I|��~��y��w(��i�[�{�~�n��Y�"s����+���3կ.�J��@ir����.؂�a�Y�ܐ6A.*('������{�6��	�E��$o���awC�9�	���!i�6;���-7� �qhjb��P�ֱ�h�Z�"F��fe��*ጾ�E3��H*�M�b]���B�T����K�L�1tb
�>�`%�D�ke'bI�̻&�ٝ���%����J�G�Vĵ0B$+[��\�,1�U0 \
m�C�Xkg�IbxY;��B    IDATOF	�AL�.��	�v��0�v��"[W׷���凛ǯ�M�_ێ;���@gl҇�e҅��0p�N�g���v����ݙ
�+����~���}*$1�Au�GS!Xy`6���˫��T?Uh�!�3�{Dug���؊:���c�a0����2Q�vu�6Hn%��	���;��3QN��g�z��:��qOB���X���ER�*�,�	�a�_����z���w��T/l��}�jW)L�
�&s+t�,�ʬnﯙ����b"�nS�<&<Q?K��Y�ٛ	Ѷ�4\��$�	��\P���fB[�/����l�~w`�+�9��
���$4��\X�+`X#Fv=˷�wW��B)/�Qo���K���O%<\��ݦ�'>+�&�zh�c������c�ao���k^�e�U}Z[�M�]cFrc��$�۟
�3�~.��uRgG6cY�}�����Z���-�\��vw����F��$i�,��z��`p(�����'p�_2vL>f�X����������ŗ������/1nE�$��uU��7$��z�p�j6Zʹ��|𹡃+s�ȑ��̅�C�~'���b���G�� $#HS9��l��QO�=y���l�?�*� ��TR�l4��|Hdl]�o��ӫ����'/?��������$M���$�����>�Hk������kJ����a��P��dԏ֩�I�Z�Xc��a��\-�g��W�>�l�5$��e����ԓ�h?������ډZ-��_��Oy�B�j�h�,�T ��	+m=%��72�[t���ҩ�E��y�v|���C^�k/�g��$ɵ1��p���)-�-w��nSF��Z��N[��l}ߝ�o����Ƚ�j�BޅU/���u1����q��l��=�p0P,�97��v���9��rU0Ez�,	��O���-ќ�
1�o��3��B�~��h9�Y��Nl�2��u�`.�a�N�.�xض�n��ZO����g�ۛ���찤�e�L��"V�8a��cW���f�^w������r6J�6[�jY ,T�e�qʵ�h��iկY�B��� '�@���P�h�&J���������	)𖵨��e ��,P�g��vW77�����Ќx���m��2yT�Uc�O�L��:Y������Z�-,g$�G5yEy�����j��W�|d����Q���߲ٗdm�����C�;΃#�㢭�̈́�Y��h8��~��_a���|q���f��/�
�@6�#����;�F���_�t8�e<��Avw��n�ݵ�;�o( �#����������(�ʅ�H�!�	[����w�U���k.���/��v��Y�Pn���?~�����j�5/AC���I<T���!��b���X���첖< <WJ2T�@q4��QV��K��Q���YW[
�ԶR��ʳ�C��J;�w���	�Y����dHc|Cb��J�hԖ����%����G��
U2q��f�ݾ[�����#$v�V-�L�f�`�k����$�
�����LR�	OyLD�J��R����nf��Q�+�d(˜f�}B���B�NDd�"�d� �r�'�v�%%B_��o��o6}CI�V�/��*51v������ND�*��JI���>��I�{urМ�W��ug��;ػ��6;�B>�I�Tlm��ލO5�l*�$�&o������A]ġ�H��;��I�b�~�^�����݋R<��yP�g�o$�����R�\�Tq��N��bT����Ɂ(-.R���ILa���"�v��")',�a
Y�V�9�W2�<�#�@�?m%�WCk�������d���VO�g��	�T�N+V���գ�t��
zPs#�6V�F������q_����|+��#�&�~���Q�qZN=��Ҩz�tB��l�>�t���~����ߺty���?:��ÞXِ{!�$q�d�M��t��!�>.t��B{�U�C��8;V{�ݶ���s۹:Y��i[ �OT�-�k_:��Q��}sNS*�VҦ��=^D~3O�D|Y`{<����-�\��s���G�m��0��S0?aѵ����Ӌ�KkmQ
�}���x�>�^\o�f
�]YA��,����c�L�e$����s�M�QҲY�L������7벚�g����jff''MӮĨ�zOb�SO�_r����	��
�� �OU'܌qޱo�ꌓθ�=�%~Q�R
"���Q��Ԇ~���Lt��CFE�,��4@T{�V�A7����N��}��:Y'r�����}ټb^����"���RBb��u�C�˴$�{�v��+u�;�T�4�@83X6Ug��~ A'I�҃X��,��p�J�cRl�5����	���T.��W��ޅ�rbgbO��,�$`:���lU,,�A��7��� "I�z����&"4 �� ց.����j㗏?5�E�m#�d�d 壂�`kU�P!�-�.UaTC�Pn^*�iB8����%��]_���Y!��������(q�q�࣭��lg�S�G��A�5=g$_w�6�bM����bq�i���_^UDAD�dN�ig�A���"���=�գ�Z�P �������W������?�'E��W�8�i)���S$�^�"$d��M��^��JN6�K����f�8@���8�n�d/ �F�A*�@�,&,A|�EQ1E:K�z�&���O�<#���P��Ч�6#���h��G�L��D>�6�Eu{C�#[���!���>
���:�胭Fy_�}\)#�Q���D�w��;�~�����p!e�w��-�ب���* Ҳ�ç��@tKw�G�����-4`p�q�`���O*�$��Q_�>KB�-��  
�1Z�Jbd�Y��Pc�#`J2���l��(���@p_�_-�>�m�� D�	���0A������B�$�$����E�[�p�e�m/��kH�	�i*m%в�
(>�,���1o�QN��h�!%:4�f�Z�{�͔hk4/N��QO`��A��ݥ���$�)$��dXz�]RCHb�'����N*����BY�Cm��I�����i�jv@�Osx�N͂���<�B�r�Pc�	�&��h�1�����#8!
I�<�f���D=�1��,���I�$�BgY�Ya1��$I�8�t��y^,RG�4���Ewx�+J��F�[|RI�H��8A
�,+_r�S��*j�O�������L?��3��c% ݹρ̬Z*����
�bQ��h0ب��^D�kЦ��G���W����E�U3䗀_l��3��.O�lI%e9 �2V�pZ@rF���1=�G�{�����YߝD�pK� L g�_�iq���8���JV3!�ݯn>�t"�"�:I2�f������s1qo�ϖ�^x�c�ǃ��V�cd�%[!�k�;PNI����{4��V��B}�擁N޽�&�����mM������k,P��ݱ<ϞHA�z(o@r���fՓ#��$މ��Ǘ�W��uZ͒�IԚ`Y�����S$�p���OiE�T�{�7f�lpjb;~8���Ʊ
�yiޯձ�LP�dՐ�R��j��D�^��
���i���p���NV�8!���f��K*�К�wbjxX-uh)U�%Ȓd�Q^���QЭxc����H�IC�ō�Q�˻Ii\��ŗ߻���9�i��}����$���s�gLE*�!�՘��wh��PI.*վil�gg����˳Z}���  ywW+*}��HiL>�-�lQ��!E֥���LgA/��=5� 8v�V�\a/�tl�|������;�����зձ��r�㞎�d�K��:��xk��rށ���:�������NV��'w��맂y�O�B�������yW9�r� >���#q�4�,��{"�-A�m����l�#�D7e��G�ĭ�ecx
������ꆲ�!C��c�zH��r@��2K�a2�G��kMmXru1��B)��MpI�4�\�d3wDߥ_�bR�m�j�:5TV��L�3E"3�(�Ax�L��Q��m�
�g{�'A{^��a"g�2�M��5��L@��qu'M�d�}�#ދ7O�b���ʚ����� �lG�dZp���Z��}������Z2ӂf#��8��FWu9���y���^���U��������{�O��0,z�t�Ц�t���:��k
�ҿ�~u[����/u^�鷸���I٨�X�W�^����E�.�{�a�<⥮sC�siItR&]K��N����˗�%&��'8W��gn������z����Ao�KI��9}�?��-]JI��m��u}9�cb>�m^ψ����2v��'�?����������-���-�P�xm�\|>���R��`���L��h˟-��������:���M��?F�(���V�?)�MR����=�
�gAc�j��l��D��m�6��	Rڼ������#�O�MOH�6a�RpB�wI�7cO|$:���ɰ6db~y�L���!Ω��fq;��e�ٷt�m��C��T��[���m֛�cX��|5a�6��=��Z
��J�J�9V"y�x�vz{7��n,�~�Mp�<|*;�y����Q_��i�3����e3�8/�|���:�QF�+�T>�{Se_\)[���bL0�|���-W,�c]�X�]��G�g�W@i�M���\AE�
������̻�����D:�ʣI��V�'l�9?��m����Emu�a"��"WI
���W(o|�S�n{+k!�o�n�)�($�A�ޟmg�\X �$T�)+t_�x��^��I�/W��hB;�Pe����R��݌����ˋ��q>zx�݉�@�q��`�RQ
��⠄k���(�Ǌ"�-��a���u�h^95�e�SN@���њf�#?U�|��E�)��c���=K�'g?�Ǎڟo�ߒ%7�֋'H���pB���R�|ӝ�v�T�;�K����?]���O��W�1��FR�b���鰨��"�D��v�)f���X�t�:2�j��hB��0�_W>\�Q����3U�#�<����9�c���Mh"��I<���6Jd�,;O����������/)�7ۙX�B	�Nd�&sD�3���v&E��-+BxT��z�\�:�1aa��$D�ʔ�	�9�_��-�u1�y
^�K��r3+��n�����tt�i.*�i??�K�E�{�L�B�]��Jġ�v���w�g�c�/ܺY����l��0���fIr�G}�'&���6����M��J�u��)�2��l?�X5B�O�9Vz�z��}����8�h�1����#^_������'/ˡ�2[��k�s���ϸ��Ǎ;���Ra8�P!����W�7�[1�%1 @�պ��c�����c��aO�3��,'��] �w#1߼Z0*�DI�v�q69���Օ���L/�d���ζe���/"�
�UI7�L!x/IK߬h;(��H��r�zk�@�Ȇ�=K���R 
_�V��M��n�}�S��z���?�|r�^�V��vC��&>�R�d�`-�x�r�HÆ�����m�A������+{�f.���+��~�>�%"�^�g�"���ݽ���.6�O�Ng��oۅgMr��|ύ��$��8��S��$��dU�\���l�z��d�욞�Ȧj�Ӟ��b�k���a���'�{��߫�~����̥��BK��E��nL5;�
�v�g��: Lw����h9���|ػy��B�����q��=���Sќ����Ջ.�����rz�)��{^0՝����\V��G}�<=Â�B8�4��2V��=�`-���0��,�-6hV1��{���>�C8���b���Ԉ�n�,%��AY�K��@�D �#*�w�\�q#��w/�����qru���[/�"�ǡ�JB�b<&�V�c}7�=6:���έ9s$�"���&��3I�! U2� ���A�1`� �4>��QB���x*��W>�2%�f�
D3c��,Hz�b��N0�e	[�T�U�dF�����Q4*�O_܄�:�1�c>�.��(܈}+����TL�Mu�?�ǐV�����+�"�"�VՍ	o�B08����PV�J�����������@[L�]h{�g;�c�`��r}g7I�h�H�o���nn#�>��&�ذB�OY��^��XJ4M��X��)��Vq��ZΙ��_]��5�Kj�[H��ڡɝ�	qK֎�~���/r> ��[���M���eG�ԉ��f��)%%��:�t��Wu�.����/+�;^�9�w5� �=�?%����pG�� �q���Ȯ`��M��?�}��"|d�yF%�K�cx�����c���J�S�<~��`=�.��}�����D@��MTn��}���bJ�(��0s�����;���9�4{f�w�0�@�x�rY�)?|�9���V��5� ߊ��&��� S�0[�=�'N N��ve����@�L��fm�KĿ�MԉID�M�Zg�P(�0>G�ڝp�H �̑�"|�B�L��i���s�鸑�P|�v'pK�3z$�Au��b�����`���ƴX\�1�����$����#[I[��U�Z�ޏ���P{d�xE�/i��.1r�� 1��k[�wdR�mAll�J9�#�����V{L�g"�$|���c�������L��a~?�?�V[��7Ϟ�q~��ٯR�p��=�~[�2�#���7�{6��L�Lݒ߫¹��t��,��x
�>�k�5�H%�D�_;a�\���޸�}���$����"���פ;[��:�ŉ�P ��Zf�.�І ��y�L�C��*���	�Q�L�������ҺH�����@��>� MRjm0��T�qٍu�v��o6{�2hRo0lp\�~T��,r��c���
2�9��-Xp6Z�{�0l�:L͆Ȣ��|�3��y�fTjĉ?b�;���)�;���+bP�˧���M%��"V������R�cb@�8E��6,Ӊ\������)�і��
F}�=/a�"a���Q�� ��?��f�,���09XHR~���f��+L|š+
�'��bJ���䒱� [$�PL��R%��|��<cdv��Bߵ*3a����֓���I�]�G0tMv����ӛ�dKq2�
La?ǗG�g��}�K�S���g�X�l^���,���O�M�0�a"Õie�����qzX��z�]�U�Q���)	���-�K������tG�!oq쓃۴Δ @���Q ����[ɡl1vPr.�s"_�P[�!aalm	�)x�P~�Y����*���b>��͎]8|�Q�N�0Q�^�	̑�V�b��}���{� �fxqN���V��'���N�c����S�m1���c1�gP�qVS���󧏣�º�
9&+�>����,���o��B��I�ټ�(��1����Ϋ��Q���#�4l��h�Ϧ���-[%x%����pV$�c��D�pLiO��0�*ATw��ig�)H�_w5F���C�=DH��F,iU�ò�DW�Eh��Ic£��@�����o�g��@�3�H/+��a���s"��jv�GV�J������z�V�x0T1��Mė�,Hko��x6:=�Vq/1�C��갡�V\::�m�h�rB%��"���L���(�L�\�]�c�紊��`I�8{�eʳy��ɵ�30�a��F��>��C���v����x�BO �ā�H���_�D��Q�Ml�^
�U�����4�/�;S����4�
�[��i̞^�C%N���,a�u����_��6��qa߷�=�̘'	L�pH����}m/��y�s�r��$�Ö]<�i�G3n=�q�!��.�Y�\�����x$j/l�\%<֮���X~5&v.n�Twz��?;9*��=HUD�<�\�9hq����O���tXϧ��<�[xj�/#�h��t��� ��b5��p}Էd��Q�zS����͡�v�x���f�t�x��=l���8�@k4��o��X�H�(]�d���An֞*�Y��6�Fʮ4f�%t ������x�D��d,j�1�    IDAT7lydː�޺�7�4lf����v���5�E��*��>�}� d�\J�\��7�4Zq��g{5�5x�<4��^���0p4�i���̀�p�+ܪ��[��{<Y�M��q\���
.$?�/��*�,�3��K���t #��g�|���N�#� �W#/�T!�	O0�� 1��w����x�렕E�^����-��AD&����#7�D�����E����:�b��8v��p5��b�̔���P՞Ͳ(��C<�v'�Y��lh��l��v��K2O�l<.��'1��P=����������ŧ�lPf��%a�j�._�8%�)P�����F��xf����*�,���!���^o>���j���[N�*a^ 0��s�:|߲�Dlm���͟ec����u�l��N�;�8�q���L���]�X�㺷8wI޿џ�8=��ʧt��;)�u��©2�E�;�l��9�u��b#��)"��͢2�/wH�������0���6Ps�V�$,��t�
�k4�{�N'�s��Q�8����I����!$ 
N<��[R��CF�X����'���̣�����\C�>���֒�0��C6��ó��8N�b:����ȏ��	�%5�ƯC?�*]��V�O'z��bٕf�,o��'<�K���f;�ʈGr�+\侏��o�"���͋<�D�*?��Qc�K�O?�T'���}S���������'R>�Η_~����Ⱦ�~l9_|��W_}e�L�D�rL�A�k\d��2ϓĴg�42�dF�A�����i��P>\�<�-%,W��Y%��8�S\�u��
��2g�uhc�$H.SB��D���"E�j�j��}�-jMJ�J�|�>^�P�Zufx�I
!�-/laH;fO���-��+�gk�Rk~qm(0��6gv
��,P�vc����5̝�u�0d7�_��X�#5��¬d�Z#�q�$"����C �%�C͢�0��:1G���b��0#�X�;`ڽr3B,���B,U
B2O�Fd�O� �w�LY6w�ߍ�}s��a��q���&�,�fX^xVE�W�u���bH%�j�JyW��8�u��!��5=�o���q���uzvbx���ڸ�܉!�F�z�t[��|���xJ^�Omt�Y<�-	��,{�R�V[�>� ^��~��;e�@��/��넲{;������_��N�q7�3�����D��I0�6[ �(6�g�~���	��A(DX���*����Z��7~����d���w����g��=�'S�y��h>�v�����Zm;A.�\$�Y���J���d"��"���Ǻ�����>,sa���Ʃ�#[A���@ɧ�)ǣ!�N��%��7l��E9qn9��˔cv%�%�W���������FD��������)f���h-���:�?,^܋]�&���B��C�r!���Rzuڔ�τ�V�n߸��t�(�BJU衛��A���u������=Z�����;��\�)���J͘i�)|�|��%�SeB9���!�����G/>��b�Y��Օ�y1SI��!������D��#�]&̃qK��� h.%����#��,v���.�����ѴR��# 6t���q�.�t�^N�m�m��1��~���\}p�fR#u`m�����-¸>'�*���\~����_\�=ۈǢ�*b�x��{�G=`��C�����,�dAUL`����l��Xb_:�q;��Jq8�߬��:�������Rb��� ��ǒ0y�Ҹ��ٓ���k���������{E�0±���9�3Gcxq�&:�5���$���xY�D��@�?�t����CDe`�/b��=s�k��X�׶MD���D[@^�9���XQ�[$���Î��T�R���;&�"25�Mv��@!�EP�_.(�j+;T�hn-���Y�r䰕`���b���+��mS���վL�I�����d,|�jmE���K6Ʒٖ��R����R}n�>o Q�2M��:�DY�D���]y;��nS�� ��
��7c!�C�,<�4_lF�:��ȫ�rAe�t����l�3���8Y�kA��-@7�?z�P�Fd���.<t�qL��:��d���-�H}G�iVBӴ�
0��Ɖ`�+��կW�����C�����hQl��V�:[�ٷќ0�&�*g<�\=�lt"!S�+'ݪP����c��d���I2�=���-��g7ґ� �^�kK�}5���A��@E�I�n�h�ME�j�������;�{!Z���ëG,,�u�;<[�a9z��U;=$Y ���- �^ߞ�&��<C�uY𲮘���B7<�+%�u��o<�jtθ;�b�B��W�h� e��4r�1Q�05$���Ѿ�8������G��ï�k�(;�����z����aN�Ն�U2�
�40DXk ��£��//;�!�U=]�·]E��Ȍ�'҇�^�}���m�f����/��C�/_g�*�u�[&�o������b��1�T�)�b7����vN�R@�e�AA͌��(U�j���9@̡O�����*H�z��B}ap�C��C8��ŧwaZ�M�mZ��BÕ���Y<�UJ��N�XD�1��� 4d�3�CQ�IF%9�i{�X�T�l���MT���.�xEB��#Ya$(��Bk3Z+������/>�>�]��.S	��O�Ȉ���Jڟ��؎�	Ay� Z/����.��?��b�==R���i��6���l����d�$��[�P�LW"k����4 �+b#�{`���>$2d������l(I)SAl@vn�������8�n�2Ql��	��5�L�^�B��ّ��0~ho�ٱ�)f�����ӟ���[�;��k���}�֋'#S��S�	k��ڢ���"�F3>X����� ����n���%�]s.��<{��⫐Z��6R���FRtxgė��:�m�*���:W)�fV�뛧`���~���@��wl�\_��@WC^d]����>�Ok�-�\��q�v��d39���@�8TL�Yә��� E������[qc@5�0^
'"�Z`a�5b�]���B�BcmZ�2��FZ5�d7m�/�~й��_o8���c�T��@)Z�e��N�qS���� �����|<C�#�j�/��P*�-g�j����F[h����s#~�NL�B�L���1���ƂG��dn���e�c.>ք�w�y�<��+��(e}��%} 5�J� �D�V%f�J�Fc.�\�ѯ#B�Xr�ߒ��/�k"� E>�AC%��B�����~/���a=����-��	�������О`
,������V�W�/ܤ�q'Fy�[���NQ�}M�Y��D�I.����enGLHb,�l��I&v�#�$��g�8�K�.T��a��}b�8ɥ��\���q�_dz�G��V���趲[�4a��+�A+�:ӓuQ�̦ϰ� 8�
����06&
�5M%"�ע�ͮ�%�M�~��r�a�p	���A��5��ހ|��m6��T�,+� �e�C��&�~8v�7��'�����կ/&��hg������e��a���g5Fb��U6ߊt��xeq��ȦF��,K��vyU��\o[ݮ�ϻ��+�0,d���
��e��S�V-���r���:y���|����y~�6���R�ߍ��l�X�cKbl�e2g��q��i$�T9d�T=�P�d�:�.�Ӛ�tˈbw��)a�j1�cfabO�I&���c�Q�(?��9�
&z���o��!�e���$UJ�kmp�]��Wc��!��:�ۋ�A�م�L��1"�Um��U�W7C,j��eU,���Tm�7��BXV�m�P����/żƼF����J9�}���Q1R��%�sε�!@�>��@�k����j8Y��_��߲�]
����^8;\�
t����h��e��������	��(J�3Zy�o�@2x�G���
�-ZBq�V�k}ڮ�_xs���RP���2A�Q;,��0�͢���=myQS�*��`:f&��:@'p���_6/.D�&�(�Wmn� ����a��Sjg�n��j����D��q#���c��-7�|y5��x	�\� u���^Y|W|G�m��E;%�<�[���w���Y8�d@��?��S��\H�s������O�n���`��[����H\�'���c㌋��v�e�3hATz�'��\�N�WW�V�	��ԄgM�؊��Z������d�(^%�]�4F��KZrkF-V�:m��Wr�aN�L����ȅ��hȬ�V)p#���_2�)vo&�����~;�8p���	�j7���ap��΁���`yP�j*HQ�0d�<�qGA�B�����$�l���%�ؘ����f���n��������H���lUbv��S4L�t酀K����Ye�Z��Y����לlZ�3�T��*�1���c_"ϰ�����	��q�p����%��Ƴ?�'s�eք�q��D.�'��h���JrjHf�yr�z=\Mף�rє�XHe*�H����h���
����Im��{�p#�0�1���A/d�|�ɪ��FtȖ372���I`0 �j����Q��P�Bl��%�P�{:����qW��F��7o]�(·&WL6��+}�X�|��Ӻ䁇��2�@��o����5rVh�O$/��9o���p�zf�|6���S��_�������������o޼��<\����׹��=a?itk�K�����쪯�L���o�m±�lVV ��)����ɓ6�� $kU���wPĴ	�A2�(��~a�q���s_I^�������K4� �攠`��؝�U�Y�u^���P>�J���Jy�������]�S�{��i1��Wai�ay�������wͪ���W���-e��O��hV�Yv�u��\���k�MIl߿?D�{����?���Ş�R|�bSO>R�+N������B�@_"hl��f/b��!sw�Ň��B�Ǜ�sI��D�ϓ��w?x�iQ�pc2��
�EG��W�¾4֥B'f����E���K�d���-���ùfAЂkuJ֩o){pݨ<�e�^�e'�{=�N�6�rx�E��mt��tns/{����ă�)zʇx���]�����t���B�8&^�4gj���c�����k�e�HE���/���=����=��?����˿��cb-��k>��C�3���9L&O�'-������\q]��߀�?����&�?]כ[�]�ɯ?}���Չ+��bp�������Dn�O��38DBe�b��K����A~��|���W<�0-C��-��qrG3�h��z�eс�:&�D՛���,�801K���=2�K��vQ�:(�?���NnQe�Bޕo)Mz���;�e��:�)߈S!��gb���*?�/�� �eO��$���xg�A��$���v�0mX��:�@yT�8]�G�C^��vM^Zz\�?�B�;�Q)[�l��J�~��n4{7�{ڎH�MȰ�C��rB����ˋ�������uR�x��G�}?�e{-=���u�͜�Rvŝx�\	nA��}y�]�;�RWν�����N����kq�|u�=� 폇gJF�x��b�����I�(�w�����ݽ�U��Hy�翵:�{a%��t`�G
�g#��O�4�����YVa)����1:��Ui�.���ϯ|�:��eR}�l������t��D�w�r����UI���
�0}�O~�T������8.����?� Y�1M����N:~�}�M�R�.�$)������\A���
���(a����y9ݧo%�n�袩j������_�z'ԃ�竷�yoѺ6�y�"���-;?�=�~x��o�����\|�is�x�V�&��:'Q�P~���F�L�JO_E���ȶB�=]�[$&�;�6�7�FQw��d�%&[��}��Z�]�.%�\��}&x)O���Uc-��?��^��?���Ooz��+�a�|;�Y� �%�1��"�������zk_�iWݏG��=��
>���#z҇�ho/����Z��X2���+Hq�=����^�sɩ�N*�B���w�����]��XE�ɣ�/ }���u��A����m�.�l���N"�I��6-�\��"1Nfsz�'��Yfz�\�Ծa�� ��*H�P����CPA� ���4�v�M���¡;�������ꨆ.�D��h��_�Q�r�=�%���_�gI�y�0�+�h$�uZ�Y�
A�(+Ҿ��a`H����h��Pь�
g�x4}Ƚ��)�1
$��J�^����?��lβbJ��=YM_��O~�[I+�)X0qN��B��G���0�!������?�����O���:b��w�zE��q�a<�O��'q	?���������8k���������a6�uZ�]\����9[�|�z�/"k�v��q\��
 ��5t����\Q�Il�ɋ��D\����������
���'T��;:t�Jw������0�t��C�]��	�n�/�.�hR����u�ܟN��$\���o��5�!�����d���0�k��T�P��k��� ��m��_������a��о������ʏ8��QR�(6��v�2�q��CT]�ą�8ނ9����[�%�e�����U�/��J������al���+�A{gW���lKX�y���o����1������D�^7��j�֐��j1�VP��R��LĊs�^=�nk�x\q���A����ż�a+�S���S))�7;��;q���;̐.�3�6={�DnʡmK���H���1������,�<V�6ͳf�0��4���\���,�q�լ�	�[%�,�����.�s<Q�٣b�˓NZ3�G� �����r<ݮ�Mgzsyq=��qz�ΌY,8S���S�$Jr׫�:���L����<��<��i��\�r�¦��b/���&$l>��^&���+�����@fh��HRR"s�pA�`�qwq�&�Xsk�'	�@(�Z����F���`�V8z��4ՈP++��F+���������Bz�V��'�<;���nG��W�D���W��Bb��v(��Nw�V��*���/>���z�/~����닋+��UH������>�kbPTtS��F�r�08���D��ru*��ի�3����
���r��Z�4�Y)���/J�+v�D���Ҷ����Q��6TC��<L	� )��Yt�)�c�	���FR�߀KJ\��i��MW4�6H��(�m��Z*8X�RXxmu�&��̗wq��z�I��7�����u�F�[�|�K�V��8V��Ո40��@f=z(�y��0q5��VG����lʢgԶ��7�$�[2���ի3E7��l.,7ދw�1���p������ݚo��'�_��}=8篸.���8#�H�xX\	)��}��ټ����MB���ӄ�DH#S�����\F�Q���pe���K���P���� ��֮���Q����t�,�����(+���ʹ*u1�Xx1�bC�mo��s>���o;���T^��^IIX̘5����r�"9,��S{����G���T�_'���|._%��Ġ���,+Ӈ�y�kJ1H6 ��V �D�|����G�:9�-�x�pPc�fF�ޤ��g��oD��T@3�J��ӡC[���F˰�7{k��~���A��Ym<�(|K|,��񑏉�zr�d�>\�b|�2��Y?�����:M������t��g��o����*��:��*\�$IT�;�=����r�{eM5N����r�yj�X�B�!c�v�@O.�/a�@��f�����OnΥP�/q������?�+]���Pq�(�#?�ޓ
�n��8;ȇ�����2v�R�AB�%�����Es�_J���0�B���E�u�%KJ��s��):w^��4�q]�=b�����jٕB1�{t�fCD�10A �.dG4	���6��u1<2�ɖ��<�rv@*����O�g�>֗X��4OT��v�@�QW�&,XC���:�    IDAT��^����9JKӽ�ِ	1!)aP�T;��M�u������U�+���v5��E�AG���'_��RQr�c������!M�L[U&�9^��sNh�7fG-�:�ͫ �L��o�F �g�Xgu�f�������Y��SSb���&|�� oa-�2���F��u�U��Տ/�K�p2~�߮7$��mҜ�7�jf��Y�sT��v��7�X���a��=a�����Ϙ�Z>��ݾ���-���D�~q�d��U�-_^cR��4�'��0�T�Y���[�F�C�O��+�}�G&󨼩���8��l�7mY������o"���p?Al�
��%�$�8���%�T���(��Al�.CO��혇����S��Y��{a��,/]�jsG��J�߹���S�lQ��ؓM�l�WB��uօdݢ kj�C,�,��#'C3f1��e"�P�I�����閼lÒ���4���9s��Ns(�)����Es9����i�U��ۦ�ܭ�Xـ��0A�"��$�AK&|XN�w�)��4�"�c?.A�-�9ЁaOlWLC(R��i��j�Χ*�.�goDA
7��=w�۟P�/�~�lx֗�J�	�CZ(�)��l;�X��gґ.ex�PZC���KRaFY���]q �Γ�!�cˌ�����dL���j~���E/J��;�Ո�ȡUMJ��8≕�+�4!o�Z|N�_%Q��]� �VY�L@�^�k�4@q;	�5��)p��s�*@j/��,T��'E�t��X�`9HW���-ȉ >J	����C��a=A_�ݷo�O�z^�C���De݅c-�|�*H��������	��~"/�#'�@�a�ƴ�^����B:�
Ed�D��ͦ���z��b�I=u�>i���W�ȩ,3x�_ĜfB�V[m��~OҠho��G�˔�Qλ�٪r��Ә%*��(
0`DI�#���r`*6%LZ��oO�e)���5:���|8��w ,�5���"y1w�6`�<ʋ�hV��]�Fq��b Z'
�p��O~��%%��Q� ���u�<�Us��������aD ��`.�7�N&����~���`!�|Zk�~��p�%RZ'/�����TO�/�~P?o�;���4��6���A�ߌg�"��!,��������z����������WAL6QV�L��"�#�A������a�@���o*�dBT�e �
�#ˀ��J�X�e����9Ѧl��
I)��}4~�H0;%WY���=�玿�l1�\)Ot^��j��'/G�q'e��O��)o)O����7�S��AQ��8)��ܡ��F�X�+��(�'���Ƚ�I�n-Sa'��p���,�p�F��k:3뀖hY�pO�9�yosAw�����1�id��
^̢���x{^Q| ���&���	�6d7cE�[�`4&�p��Q�P${�Oҕ_��D��]����6 ��ޢe�B���.j�W���t�+\)g�Pu�A͐�5p��.��E҇X$�-��G�5�9k����-��Э�������/�T}ܟZ2��L0:�"wu���+���a^���̩+�48�'���d���,,:�[���¡�� ��4s�������Q��X���1y��ޣ�Ѹ^vX��S'�9��uG	(�x8|@x�b243i4��i�������%VK��Um�P�O�����^e�SE���D�alQE���ph��{�חc��,ĆL�1�xB�"�A�p��E�%r��u�?ɪ�H�wX5�.��
��ƨds��u�,�clH�T!�E�B�~&�V�R) ����.u`�^�'Z7��y5N�L2�������$�A��|��C+ӻ,N+k5�%>�1i�|��0Y�|sϷ��R|����|Pa�M�椘� �Xl�N3�2x?��04+o�':�޹G`yٛ_m`��<�~�q�p�n�-u��r`eWԦ|/d�@Ɯ���xf�6.����z��\?l�0�`��l��ukF$+�AK��4;��B�]��睍�O�����'�w�s���n?���ANiA�\D�B���w9V�U\̧��Y�!�G�F|%����]�[�~>W�*e�����EM���<덏nڃi����)�PT��� ��?^=�}�ٓfc$2��2�3�ȡ��ὖ�WSh.V��Fw�_'1�Rġ��z Y���3^�^
Kp�����}�"'�i}�4�'_xȅ��|�v*��ZS0�C���|�y!bO:�����y�J�\&3��ow&�=�Ǝ?���]4��Z�@3?m�vhr�c���:�V����舄��c���J��h멜�&��t徬rԻ�w	���M�\ޣ�`��z(�����V��w·m+v)��L����R�H*,��O�&���cU2�ē�/L
\7Nd�F�t��������CA���@,H�5Ћ�\hd�H�|�#zY!���z.�'3��ŉ_��5	���B� |���@��\6����R͕��?�D5�����{ݿ�G��_�^�]���ڪu��J,�c�Q�;���2����7:x1� ��ò�ɅB�J���5IQ%���B
�f����L�.|��~1#��lR��ē�������q����o"��&�x �X�.�<��(��)�����o��E���o�A8v�|PJ��(���l�`��$���`���V�J�btɤ���=}ڧY��};z�̂���VU���T�Y�G�sL�."���0@����l�.�7�>�������7��cw�KQ�DS���cԼj�t���Qn��I/�e�!��H���em��M�K�<V�G�A�}a���Ϧ���tQŒ w-$�K8Þ���?�ڋ˦1Z�L��泻��#��Ɓd��)���Q�Wٯᩗ��c�Iet���}��Nt#�j�mS���F逧�Q��?���2/��J(��[��ͱ ��U�X1��(苅���@NSX�	J�KH��w-�W��4���}o��ZF*�\���Y7ϟ_'^GAzSŻ��`�<���@0��Ja�_��O���x�S͔����0�3a �ذ�u�}��<�"��'1I�-�/烟�\VQ��#&��8J�sm�x���{�P��Ż�^�پ�L��^��y������lv�
B�WAP�N����U`r��Z]�2�jK��4��:(�G�o^?|�C�M�wS	'"��@+�	A��������?x�\l~����M�a�����x�z���k����FUu���E�05�v1d�E>�y��Jlr|��x�$��G��ö�FT��x*bd����ux�E�%y]U����������9<W{v�T�ڌ��ʕb7�o+xK�ct���v9S���e��,�2���9���9���S�4^�$���wX���SLV�#�?�=��h���>t0K��"G���0L��|��/[!��BgA+�bvu�畓Y�t��d=o7�8n���L��lH?x��%l�(�e�f{�0�F��������|Z����G�[/v�@���7-�µ�N��,}�I��jJ�G�$�ݜnm<�eZ�o���v/4�a�0���������%F?�mѿ�1~'��7�z��V�^�=j��G�-.�0�	�1I��jM1���x��(q��ӹ��Y����9��PU�i��U�#�F�N�@��)�XD��գ4���Ɏ�X��E�};�u�E��D�rhcN��/�#F�狤�#���*0%˸�0��(x��6,h�tP��aJє|�L��}w8 )�7.P\�8p����D����+*���d���'?�Hɰ�OX�1�?��'삍��1Z^l���'
W��	��,堡����
=t�ɲ����N`#TNS�ĭ�:����/�K6,	�&���:�� �r<O=��DK�廛��kr��t/�}�w�{�����������]����V������c
_�GXw�'[T�UE�Y�Ī�A�B��oiw{w� q���c7[k��p���j��m���^������%��L�La刱�֖~2F��B�*� �@N_�"*J΃��a�i�"J���!�6�/�;d�\�zp�����2w��/������6I^&ط�U`Z�Y�~��zrp�ߛ���t���5����6�'�Jy^�>���U��a�vC���{Sb#���D�U�D�!��)H�^d��z"&��Կ���U�e"A��F"�
2@�`�,�������i����*������)ɘ^0��P=@4g�(!QW,��[�&%�)㻆9(��,�{u%�V����)8�g���}�I`�4��> ��R���VHxq8�ڲ/�����E�CX'���/z)G8��1SU���y����7���N��J ���@�@Cj��:��!6��}s���)I�a��G�,`vg43���df�%޸&���]����>Ĉێ��n+E�l�<?/��R��<����Ĝ�����;���<9���� �A��+n:>܍���/u���w���<�%r�9�i���ٕ
��C�I�l��e��ڐ�u�O�o���� $ֺ��Dv�%w!���X%O*�=bؚ�Ӣ��q�O6g�����	�} ���M�j�����&�q����d�dM:�
A\�����H���}eJ*���&���k%�ЩūRTE�j0<��义�o��ٲ&E���G?��jxa�m7��#�6Qn.�p��!#��`uY��b}���C���'�	�p�a� �v�e%~�z��R����XA�}�W��`��Љ�ZKtl�d�����vz��a��Vrq/uO)�I�zpqګ�\6Z��Z4Ǝ �Hh�.��3Z˓e��Z��yp���TV���,����iUd@�6�r�I��&5�f���đ)����[g��b�V^g�Ɂ�DJ��Nd�:Q�����d�	�l�Jy>����d�Bձ~�c3	=����tf�92�ڀ�m�a��s��48͉�V�-����>���߾|�k^Cx�`	���@�=ե5%5XN=�I�6��ӧ�^�f/����;��B� /P���ķ0����p�1X��z���[��+�NГ6�B�걉b�x`�y};�/��7�qУ�����G"#_ę,�i������^�Ln}v�b9<HM�52���,Rw���*l����¬y��+�4,��`�R��L�&�(��6]���@�\��T�پDi���v��B["�tâ���cK]��=��&C5-h�u�T*\D_��8J3��mѾ>n*�M� �-.ӛ}�cOa+���j�e�(�1�-�%UO4qV #@ܿY�д�o�se���Ʒ�#��8�7��cRm�<����F�4�g���[���Li����d��޿��C��k�%\@Z<�T�n�?,�'�8��L��������D�.��[� ����y	g��)���i)����Pp�� )��uEZ�{է8A�w� 6P2*�rWC��:f �[+�F����j�pR�G�8%Qӵk�{G��.�����y��%a:��o_���������!a'6j����������gϞ<���tFgp����qI��-%�B���] 	�������r��jzo��9��cC���l��G�1A,�o_����3�ݦ�Cw\%��=L*�s
~9�,� �Y�k՟�i���6�4���\#Ak�ן�k�Q��RNSٛ?=U"���1�n�gG=�O��k�G���u��ƹ��-�~\4��qW�`$ okY�߹6zv�|Q��y_�FjS~�W;�Os����j�n��|׫,�_<�p��[T(���.Đ���v1Ӥ��j�7c�?��C�myf5�dȨ�2D�|]�"�w����#�b�ٳ���P�n��+�����yى��ӡ���n9w��}m��8ѬK���O��+th�K0����Љ[`R>�D�p�hh
���~���̓k�CA�;��̯��`E\g����ޗ2�0M�p_�b���[ܺ��5��������6
h���������m~��^�]��Ȑ�k��QT_Fo�|�����/���/_~��W�k�Xcb"�:#-t$׉�����N43b-�G��Y>^N��� �6�8
	�m�@+HC�_{`��65t�����`�u�]�	��1��U���^�p��,X����{��$��4$^� 2�!J$ƍ��� /�m��N �'������@���.����H����%���O)��r��"���2��pJkm��-�B��K$��`z2h��l�vIi6�	@�^��D�$Ud2�Y�y�AŇ�|���aŻh|b<r�8�擁�&�+���������������hl|�w����LMvyL}�m�������"s�w	�w�#@>Y��T�_}����e�)-���G�:�-=^R=:<�O_��>3�a\B+�,N��r�V`����?a/�����,h|�d(4E&�ꔑ�e�)G2�6(�:�gM�*�t?8t�|�d����b�GSb��Q�@�k�W�{���X�P��.yJ-��[g-������:�X!���D���r�.�#�<I5��������v�F��8�C��'����	���_������zSy��`�(��MI|�,���0��z�ʚ����t�i�P�����t~K��6�0wW�h�W�q8)�B�1��bg��Tf�`�M��Ba�oo_oS�ae5y�)06�K`�����0�.;����������׭6����{ޭ����\{��D�����P0�c
ƳS1A֍U��Q4����v��ʓ�
�V�)܍��@d��N?����5�<ɶ�s\4鋜�QV��&��Fョ}�I�Q�� ��A>R��)�%��� ���-'���T������-+7<�u`>-Ђ�D�mEۣ�a�n�9��^�6�ڞ�qw��&%����yʌ`��Ƿ3uD�o�����{}q�u^z�f1/��
�'3�������p~�:ߧ 6(ĩ�� ��VxM�=^r�fC%p6�I���)x*�(�x�f�t�����x)�|��FL�J�*��۵N[`� Q����K3ޕ���G�Yk33�$VsD�Z'#O�z�����Tݷ��.^����-�e��d�
��Cj<�Y�Ґ��� Y@�M��V3��ۗ�B�9��b�6�v���)w������������hz�٧�����'��l�� ���1?�5Z��#R��jΩ�O�7��W��]k*�^�Z,�N1sM�k+%�:}�R��,9�2`Y�T)��+E�-�]��^�P)�!r���m�,&�*?&l�bF1D�"��N��l��
�(����'�~*��d!�A���"a.��qQ�Ӟ��:Y�[�y����ͻ�/~=��o�ן���=6EҠҌ,�P ��x88�4�>#)X%���]�@iozRLRo���3���H�2�o�!�t�d��r�T�Y7f�����������7���?�=�>_C�Oi��~�[���j�S�����:L	�Ȟ"�D�h��E�{��
9���P15�n����4�f���dz>5���p��EZ�̔�:���?��X
ȉ!Y�J�F�,��/�o�� �s��v=������lټ�<\�b�=4!�B��Q�G�Sb3���Px-�#��ο{f!["���(!:oG/~�|��,��`��|��,�̬:�|��w���I��������1ED�
�(L��\8��`��dX�MR �>�`D�<Bs޸�G9��l��+��v�h�M&ކ��Φ���E!��%W��f����pM��H�����>��N�u��R/x�����<D½0�G���1��_��+P��7jy)���7��
xe�;k+,g��Ez��&Ȍ;�m�]�k- ��%�1s7A�bb�ݴ�ǀ}��o����ݻ���O��Z��Y
Q_�	�C�ڀ��l�f��f��>�����x���8��!>Y�����u���6+���M��Y�O���T��͹��	�oK+�ؾ�r�8����y���}��v�i2�K��Hx��A    IDATu�͡g��?<L��47�)Nas�f����8�1����w($s���~|��RD^]v����jfi[q���
�$-��a�)�FIL<p	��$���jW�r@{�3î~T�y�_��U����[0֘�D���ՀC�~�r�����;O�h�C[4Z|��Is��r1�J������7�-�˙�j��dV��$}�YG�m��vGz�!({�|�H�K�u��1iH�u�/�m4k���9i=<]�(��'������� �B6�E)b���0�L="8*�2E��]ь-�a�
�0`���@�'�U������3t���O����	غ��6%U!v�p�N�k/��'��b�'0�F���j�6|1�wXV<V���9�ɉ; _+�w2�����j����~ی��z�K�׸��L{V�~q-���qNx~�q�q�?	7og�'yb�S���2z��%�y����.�������$l���)4����=�\f�=-W���?��|�����/Jw���Q�Z���b �ɶqh*��X�K�bQIC|5x�S�.D��r�?��] �ׯ+��(��o� �&/ۀ��I���W��rº9.&��W�/�1��m�ٔ�?���]�$������?�_�ms�x��kj�(�'��mB	�=I�A;|B���%��1q,��ޔa�%�9{�gy�d�\H��x���3s�o�6�*�Fd��.�Q&)%�������ɧ/��1��������*��ń�`�R�2�(B��ˊ������eU�M����7"z�0LaK-pE���>�� ���[|��S��- �C<�2#���šAa�g�R�R8*�0�Ȉ�Rd�B9r��~���Ɣ�ս��g�_�*������@NL�a<R��=	$&�H8(�d�;��hB�]�E��@%Y���Jq��(랚�%�5+'����� E�EãbE�,F����_��߈�D��h��"P5�k�+���%s�����{���h�� aө���H0h 4%lqJ���%2��*���|��n�[�1�Ü���'	���E.`�>��4S`��d�0i<�)���m��k�f�q�YN��Z��g翾���q<��z�=N�?\)����(S��'h<J�|f"ސ����L(��!sJ��]�ճ�2�b���
�K������C�M�T��'^�)3Ə>������#�#�}�8�cf��JD��U.���o�Od(�X�z�)��f��I8ZГ4-�Go+���8@�\�_�G��ۮ{�)8#N,��Q���˙�$�x�޵4M�d����i�d�
>�3|��6f��&�%J\��E���#�&���y�lx"�,�N���A����Hq�#����U0�TO��F�>n	u`�d;��zp�L��k����~��:�s|���?����W]
A�]Tz���H{T0�?��X.%����_��Z� 7P2gL}@�bg�
�{���.1_ck<�H�8���&p�7��+\�������8�����PAFh���'f�n�K��o��v���U�h��%o�Z�5���y��d6e���k��H�p	0�_�,_�N�-� Q��,5I��C@�sG���5a��]�7�����t�xܬ��o�1�M���@N�"*����M]Sߪ?0��nñ@5�~bn V�`,C�nи��a֤p�1^�t���A��%�Ϣɼd�a��T�,#0��M�<%ǫ�U�,�V޲B��7�>�����w�ۻ�ō��R�q�j7΄S֗����\��	\E?*���1ˋEt����1^x�φ��/ 4��ߓ}�_��z��� <�ZW|�i"8e���~��c��˸�M�o��~�_�oM�i
�,A���p�r���ѽ�[��Ō\o�a�l�WH5�·G�M/�kE���g�kS^�Ɵ�	RyODǬ)-3#���Aϱz�{�w�B��Ъp��P�|X�gXK'ܤ�k�gZ}�v�z#1aR	f�r^ng1�+Z��.s�j�2��No߲T>6Տ>�=���mn���`xn�O�#�!h<�G�ʉ�:�'**��l9�~6i8%��17QB������������\,l�z`�E��4
Sd�YXB_*�ozz�7~-U��Or�vY�u��dT�=xW��ԡ�7b0�Y^t��z	�r:`��2M�+m\����x�[����=�G�/��(f�I���E~���A9�������}c=��{����]~5�[�������P�.��S��u�gz
Q��uݺ�q:)_vny�*:m\)�{<�4��;!�Ŏ2{�z���p
/���دMkD破gC�����]�Bx���)�\���Hߙ�-[o�I����R�.F��d�.��` �QW@��EW����>�l�3������a�f%���k��w9�Y�i��W4({���x\$��
i����x�[�?��S.
����/	8�Bw=bHzp�g����vM�&E��'� �{���v�ӏ��'�}j�eɥ3����O��O���G}d4,�n��I�iA�|��j���/�N���_��W�2����=4Cϟ';�G�[z�`��F�Or�h�g�8ʁ:1���������\�U�
�jO�"�SP3�+� .�_(�P�k��!W?����}����"-Ϻu��m��g�����W�1*�����ѐC����1���$o+ cË{��U�#�%ޚ��d5��$A�?R.B_�mx¢���Ө�p��ݘ }����T���9��{��u������s����Wrx ��:0FOV�F�����u��T��~v�0~�(O��ݽp�%��7�[lp��V�UBMP+�|hq��{Ҭ�z� L�Į�w�X�0���w�t�ϖ8�WW�.��w�U~o�'��R�J zʻ��Aٛ���^��t�<��ß�e�p�|�*�N������\��X!98���fU-�K�q�9<�j���o�P���3� N*��Z��5� �A�"aY-���?9g֔B��~��n��Ի6����o�]Wn��vp�L�b*y�2T%�Z�}s?i%`��bMp�B�Y�PAia�������_~����:�I�jc�Q0|��ʞ�Pd��q���e6=�[����$nW �o	��Op+��VNz	U��ƻ�#q mb� �g�ް ��9D���R�J�D�~��p�e\!�n��c.�A(�ϻ?�hvR��o�O�m.���dGMޚ1��tz�����H�ׯ��A��2�Zp�ĺ�g
�N�}���W��T�qh3M�
����+X�iTY��� �P��J�4�=�=|������Ϟ<?��>Z}��x���*��҂��D�/�.�(��׷��o���y��݌NH�>���W�[E+͐�L��6`d"2 ��[����q����W^�1nJl�{ܑwo~��χ����զ���$���]U'�7��~��p�|��/�����8~|w�r5>�
�$��x�a�j�y`� :.�,L�jJ|��j�E1E�At,�3�_�]̮R1�ݱt�o����v?��F,�O��æ䓍����8d'>����j���8碽��8�'�1�%��2�:_�b��]��72���D�@$NTi>vM�B��O����Kܠ-�F�1���K�(`�sA.k�u����^�7�9�k����f�Ɯ��`]�
���`��!Ǖ���5�6��G���N������׊���Z���g?o
umw��\:��վ�l����!gu��kP�P5�IC�4��b*I�RHޑ��h|�?���PmK�e���t|��g7�Ww�x%ST��l닆�N�>XŘW�G��ʙ��e}^o����տ��o�����ؙ7>�����u�i��_�L�U"��B�ƵP�����Bt`���%=�A&��9�I�I:���6D�b	0����59R�ek�D���J���D�E�&9vw~s�������f_�b(�x���*`��<<P�L	_�vv���̖W��o�(�b)�!o������.4S���@;�A���d:�L%'_k{E��\���۔���e~��~��+�t�VIoa	P/r$V��Hj�-k>$7�SH�u��DU���cRT�I���8�Wp�R�6$Pt�v�Ml���4*������_�����Ұ��aJ�]�}v;��A�X;Q���Z�׋�Ճ}�*S�_6��U�������z�����7'/���nN���e_⼻{~�\���pI��ŏ�M��F�6@)HV��O��vҙ����ޏGlk��=ƦCU��e²9� :`��r�)\��������P�U�,)D��⡃����Q�G�^�ܿ��!p�J����܆�@P�3~W 	�
t����**����'��S��T������{1?v�(��9������?���%�7f�c�l&a�W�\��F���F���|���/F_-��=�H25����Z9�PҢ� d�3Yy����rC��(�n��ܒ�Z��as��zvQo��0�Oݹ���yx7�*�]^���\�?~ї�y�8����0�<�z������j'�:Oi_��E��<�+�)����f|=7�i��xE��/��do�ɜUx���8��r�w(�����f���T)�V�����Оo�t�����7���t�'���[������6y���@�`i�ڽ��?��f�r�5�:��r{?��wߐL���&+�T+�^�"QP�j���B�u��~�1Qu�0lH{�	�ѩ"M��b:���N/��s��-F���A�F�S�~a7�8�j�H�7���>��}��D�O�1�?K��*Ru�C�p�#e��fw_'ʊNF��?ӈ�l&���_hx2����6A�� h��3����y	dױ�y��*Q��p�"ފ�D�:�[L?[J��$���$����eYj���̃콧���՟��|�f;o�{ ��*��Qi��0����m��zoY�x5���|�b1~��V��ʷ��ޑ���N����'"�Z]�|)|��P�i۠��$�x��n6��{�}��'�\О�ul���C-b�M��W� W>�|��7�tC&��h	t���¡� ^K'�E����	�����g]�F���2T<��ۇ�D0'̕��v�AD礟���~)q�!eQ�T��+�nUR����Z̙t�I{28�gJ�I5�N|��o���F� L@�!��2�|?����7�2`B�&y���ZdUy��k�;��v���?L�y�-�u�s��s�|�{�0A�A��8h�DK�'Jv�ر]vR��?)�|�|���T�W���R���Keʱ%�% ���w�s�<��n���o��ݻ�^{�5���J��X�M[$�����+��jko՗*\��\��/W���m�96�B�<�!�ʹЍ����E��V5-ضe�,�aőS�32ʶ���d.&�L�2<�,��H>L�L�O�D61!'�_�
*l�w���8"�e4��+;�+�'�c�@�X��x���2S���~�>���}g��d���@�7�:��(�#�o,+���&�B�E9�-r{
��m@���.�H�tH��5#��\��V!<�
�^�T�U��r����@J�<�j�Z�PK	��[8�h��o�����397���;~��.k(ژ��~��X���yH����逅UX���7�)$�A¯G�.�y0|��0x�Y�r���J��=�5���44��&����2��+���M#�d7|�J�I����
�Ey#]�>RD\��W��_Ƣ>�1�<��AZ-y�H
�o櫫��1���A�`�����{�AI����"�oI7�����͡�|K��%{Z'�Qd~��+��1�S"Q(�p�;�oY-K��!�רd(YH���Y��:�H*|
x��ߚBD��g�`��ɮ������IB���.�$f)��B�Xx�`�Un��p,�#��Pl���诈��$'��Խ�ߵ�����á]�z�\]/ٜ#aCx�]`$=�����6�ãݽ�z�kK@:��M䎈B��ð+��F�ʽS��������Ȟaڑ��=}��I�:l���TJ��|����l~�{e��K%]�����w�]������ 
I��k����ܬ~�)H���.��gK�7�9�#�#�<Q�$�8�PȮP��.�}`�&��N��(w��v'��Oƪ�p,�06	y�.�Gw~��w��>z�2[�Q>4vh<�'ٽ��a���#h��Н��{��2�g<��:��Ya%&�<hVyh(��h��ō`��fYh�[�x!�ːPRd�ɯw8��+�ScҦ"M��&�@}�[ ����P��P�eֻ�Wg9� ����$M	�>����) �P��v���8Bwd�e��ݢ0�y	U�TD��"�*��8>Q3�̖��S�9&�
]�Or��#�!���������|a"�����Nl��"j@�
q�@P��e#��Q2��eY�k��;c�xEq�	J� �[nX�d<!�0"�ND,���H<,�Y(<SP��U�&S����V��ҍ�Kʮ���#��C&��C���C��ó`>;B� I<f��,;`��9@�<�?ᥝ�1L%�aJy�D�Mr�-`��!�����\��	�OO!#(a��
t��7R��e����������ç��X�xC����$qe]�o'쇫�Vr%p@T�Ѫ�qX_]p�T��Ew.MfYS�'����>�u��.���j���M�$b,��F)����:?!Mp����雟{�E�q����n����?�b��
�M���A�*ZO���8H*��eɟ��9d�� C�3fϢ��]t�u����o�F�-=�Dc'��?m��~�B�Җ~�����u宖n9wѭt�]t�E��;�6�I���
�-��g��~R�hH��s���zN�~��ҖiWn�3�▋����Q���4��)�������C�9B�L,�Z�J�e&�`!C�e�~�Y�r��`���\�#����4�;�[k��1��P�&�o�$�j�|�禃ԏn=b8�`�J���*��i㴍f>Y� z~1�dO_�$�7�M�����JO�'Q�F]i�?��E3��e�]/�/�ߌ��-I�Y(?~LrqK���#��	f�7l}z\�X����O�]'�zJ��4:3��ۙM��/��/>��G��z�7�5T����{�>&��k��PDwVz�0�B>u�����vv�g�s�?��O��ٳgn��LͰ:�Mc�>��ε�q:��Jz1i��è�	y#]�/�pO��u�j:x�����=�C
���]Jc1�<{���e2���m�vB�TN���ZE�
"��0��� �!"E�Qp뜊���č�Vo�/_~�ك��LCb��P%���Bю+�4vcȤq*WXdQ,>�S�p����e�+��W��v�=��$�+$�h����-���a�9j�%$�Hh-�X��6�_�m`"ݵ9+�f�$Fsry=�ƏO��6I���&U�wYO"�!��ځ�-�8D��X�&���It='��7��t��,�31��J{wӖN\7m�r�:yл�t@'����[���L������u����O��=w���'�şڤzЫ�+o��r�ɧ���.�UPNSkn�(�^�MI��;-A�������j���O����h�J�'Xeod���d��-?��̋45����?���7��	l<���9��ܜ���)��*��U?'�4��2)v}���������f+��/�������rx�,?�ࢃ����PQM��s�|�tz:^q��8p�K�S�NP:M)��z�pb@
�kʼ&TjA�ن�~,"ﻢ��(��d���g��N�����
% �r�6�P�K���Z��9�{��{�Vw�i�_����Gr�z��T�,����Q�R�*!��K���#��Cc��<������V�@�;�D�K.ϑ��(i��Gk?����ͬPĕ�S�NصT0_~���>8.eWUV�М��6�Q_OMC�վ��?���'�G��!;�J�2®���^8�L����OktQ�8p�L��3P�)�.mh��aui    IDATm�'�"6=,�6C9����#���z8�
��R���g�GH�|߳�Ik��dO���;��z:\�O��;���tkުթ�CU}�d�Q�J�E{�@��=���29�.�daǑ��F����",j<�	��������v��Z}����~��/�vP�����VGl�HhqP9"G�9�!�ANy�����Yy 2���j��H���+D?�V��W� �R�j��)&S�r�C�R=#0
ˡ�,��Jd\w��w����x~1؞��_�_���V���1M�L��)�G9|{2m �(lӋ���W��o��^��{������ɃҘ����/���4c^�僚`��q�'��kh�hi�v�L謩�J�s`�]�ږΥ|vy��i�7�<4�O��ˑ�����p�(��/}��߻wg����z88��a"C*N4d��[�P��z:Z��g�O{�\�K����ݗoTx�gB\��nޤGJ�~S'*�Dj�=��Fʹ�~�� �ԥ�A�)�،(T*��hn���\m���C(�_�Ô�In�qp� ���+U����;��>y�,�(�>ͳmEdfUS�@)��6�|�6��v
7n܊�>�Jnp+J��b��A"jpr+�z4�p(A��^���d�&e�lN>�T,?|�\���~�ލc��7ϯ��� ��j�K,d&�Du{z"f�B��3[���?aW�p}d������6T���i6�zR�:`��%�;A�SP����E�����v��i$I���ɋ;x-���JB��1_ɀ�����鉛�|��i��+��Y���SFXub��]������w6E:[n�ֿ��L����t�^��d���������0��d��*�3�!�h �0�>��p�j#���"��7���[����v{�A'���Bh�N�Ri2M�:T�}�n'���FD�Qʢ �!�����$�R :�F���5b��l��8@h'�$_{( �*2A�5#��B���'�e<�ߕAw3�^Xլ�p�N�P���lU��ɟt֗|����f{:���<�w+^��h���[U�؇=��ѲT��V����4��W�x��r��Hn��CIW;X�1�7�K�N�JU>"�4E`�uh��]��(�p2�Kx9�y�ͷn�VF�+<H����p.J�Ԑ2���%!������X�C{��і6xm<.���)�';Ȓ��ݧ����D2O�J��~]wŤ�Y[�g�HVA�Xh��]R�K	.c���[|�B�`i-z���M��P<c"�upp�׮J�g�|f�,��iE�j��L�T�M�,D�ވ;����J1�E�$M�l��M3�5�	���$�WQ��~f��ґڈǲ)P���؏��(P�f�u���7������M�(�l��ׄL�(s̊ڴT*4���N?y�#�H�.ރ�	�!8!\��m�.a��/\�(>@&����~�"%���h
� �vO�m(�fP`�I�wuI��e߅�R�`����r�)G�1��1^җv��Iy�?2˓�����ՙ�a���]b8� �P��0��a��aQy�n(���b2�<��G31��Vqw�����y��/V���pi�3x�X�X��]Xލu����o|���7 �f�6�wv��;��R���۬@Ћ	%h��PA	� �?�Jq�p= �88�'	�������Z��A�?Qr����h��& BI����5�b@�*�A�D���I�A숍Ɓ��LV�J�s����j�{�=�������9�qpz�}�͘h4ŹA 
Ԩ*B�ȥ�ٲ��[�Z�A��p)�@3@�鱻+����Vm4"A���]��e9�c�k(�]3�)�_ۿ��H�EօĘ�F�$��>Y���Xq DB�i�gruy6���煩L��B�-Ҩu|p0dK�x�[�IL࿐z����vh�-�9�?�V�@�R2��3�K�H"�RZ�JD^+���y;oy�֚ʤ�ʯJ��弖������>w^���(�VU��V�C��Z�%�F$C�u{c!0����E<���ˣ͏��\�9��J�-�Rͷ��Vo�i!�S��?��|�g����nk�k_{=+�b�J�����S`��-�x���NO�a��x{[�,���c۠��զ���x�C.=X�i��08')���0}LV�Đ�I��FjF~���W<�"��H�LN��JC1�,S��O޽�Zv�Νh�]Gx����"�^���ȁ?�d��w^����'�?����ļRϻ�miZ�A�����b�g!6������FK���p<��L��{��z����f�����D$'�]Iѓ&�7H�THݲ��V��(m*���q��j�sc�rQ��d����8#�)F؆b��[�q$������EDi�Խ�O���{pˡ�
����X�i�IⰎ��3���k�Sz�zz�[,�(e���9eB��V5եQ8-+��r�Pȹ���4��;�������3��e7�%j/| �֘�2��ҕ����fS�3�+�1�0�alM����qt}yE<D
�J�7y\�'��*_�Ћ�+�P�w9��s�ww�oD,�>I��q�M�Z����-������(-��(:�c�
�+8��t0A��,;�����q��A^c}F�t앉����`��WK�f���A�o�DD�X���)[Y7��H	[��0�/� ��J�n�-.l���7^zp1U۷�*������;��c����?<����e�J��g#RJ��3膠�zs2���=Em����M�zh���s�;�Q�����r]�G���N�oݽyLH�:�[/�n(sM~�d�;��m0EQOT�X����1��lp���DX%�ׄ���uX�h���'��9
"�l��(�髹����kjX$+N��EC�>	�E�P|�� �k�A�Hb�)>��r�U���׿���OX�+�mP���A#�V��yx@�|z��3c0� ��WQG�i�]����%w��\�B�{�`}����E$,��x"/o�%y�єZ�=Ed������Ha��7O��ҫ�r}<��I��pR�����$x�ڤw���s�@x��%�U�<�H�� ���, �iH����Q��'Y��3�=}�+��i&���\��zݳ�"�1]><,��O�����P�8�Nh��hG�O��=��$:ѽ��`�א��R����­�P*� BC�g+C�h��0�]h����~	"�6�5tS��.a����(mR�[e�f��PS��kB,F���H�k�5p5b����$��ph����Z��1&K���������A�'�&<l8F�����T�f�����#�z\O�:q``�E26�8�,S{��Ǥ����N�w�W^�B{�I���Cj�Wc���]��2����#m��Gҗ&��bL���.�S��g�8ק��u������O��m�u]K��5� A7<v��>�5"_͵�S3��$�A���gT�faB�/�!Xi,��
o"�>�wBۑc�7���Y�� ���O2�68E��d�P>�f����f��+]�@'>9�?/zp�6H��ٴ=� �B���Tz�Vڏg�΃�rxc�v�����;4pE�z��.��P�z=\d�d(���#��q��qQ{��ӭ�O��{��Y��a�,S]�A��O�#��vPW�߽{���^c���?�#	h��A��n�u�t�����;qQ�K��@�~��bu�ݻ�p���P�A늕�+=����PQ�n�3�K�a���u�祩���ޯ�b`�i@8a��t2��	�>�]8�U���� �����iq!�$<K�JW�3����B���.`�P�����3�VF}����	MM��s�����8䞝 $t)j
'��q�RH�/�y��P��_�R/�����%Y�Wk"�ppv��&bK&�ஒ�Jf	�[$��O�hƊ25���}#��qD��Ι��?y�����}c�MN�=�)1��h�c5NHX�v��D��X�xӐ�2����s��x*��t��c���괥�:w������y�0Z��C�I���zڹfiO�!�����]�B^��ӵ��j���'�G�$T�%sS�^�Zƍ�^�	f��7�%�)��z��6��p{��>9k�����d�������?����I�tRVPjS�jJ�V�Q�k6�����$\כ�|y`�<�Q��S %D���7�R�p�\hW"␞¾+N��x~%"�	1�>G���wvZo���w�w�q.�}��_�G�5��+a��uL�g��fҲ��UT��j�-�m�`�v��ӟ��J�S����,�2'pl=�����k�4y)�UX�,����]F�v�x�Qn<��ƹMN�	1pC�ϫ�nZ�r�D�l��
oZٲ�y��@����}��\�ڹ
[Ķ\����ɼ�$�K��*�i��#"�m���C k�j;]�2��겔��c����@�_$B}c)!��Ո]c\CX�[���o4��^v��p+h�f�pN1�F1L!��:��@>�ڛ^-..������l�r�v����r�!��)�s���p��
�j�43�f�̣���L�.�,FZx�m��u�f���g����jVY%���"·^�̷��,
�-�Ө�k���ҽ��?�f�M�gW���B����B�ǅ61c3I��SPߋ��� �G�/3ӶL6:���\�b�s�E�*WN<��-����=��}�od��=�����;w�����U�%��`IP4����q[�h�i��\Y���ӧ.>�O-���5�wV���F/�#����D��V�֦�����'I���
ґH��>��v��s���Fͷc���̲���7�����0/n�\j7r� ����'aFܖ7����A����u��~�'�I�ų��u�2<5�e/?ΖE�rv.�충�֨���cY/e�#��V�z�D�d)���[<w�-ֻG�]���-3[8��ԱY����3��y�~��߸sl�}s-��ń�r dcC�]E�d;��P�p��gVh؇K�l�pZ��_�d�]��b#��u�k�7,+��:`TJX\A�A;%�{�V��$�d�3����F�vi3�^R(T��zK�@��	�Rt|q�kv�3�ἽjUN���&sʨ�ȼ�w-�$y�"�h�r��󷚩���#��e=�.{��Xa=d{�{+�h�Ma(f�cs�n۪'�����=�綋15�$T;����t�������~g��p99�=��*x�PD���Z�Ku��W�!� �����Ç?�@Ά�tB*b{R�5cW7 �L�Q�0.F�QH#�1��I� �ϐ�v_Ȧ�\�������b5�?~�����m�i%l�N�O�a�0 "@ݿ;쑐�j4P�R=�j��J鿹�zxwT��_N��������Y�p�t��"'mM4V5�P���C]l���֛�IT�G\�+*r�{(_ғ�'�����	r&��S�X#(c������ޝo}�;_|똴�W{4�HV�Ǒ�e��S!��kd>��"���l��	h+v�
�g�v�@]�0܌*5�8n�K۟��'�P��90�o"M�=|T�x���DY�e02���p:AbSCsM���Z�g���y^X�T�8��N���u�Q^����Q�\Y;��M4����ԣ,�t�f>�KNk;��f���3tk�dIj�@��}��ɞ���W*IX����D2uN�V�f�Z�Q ���4��G����g���`Z^1f��=ɇ���,P�XP�r�G~g,;|�������U��0����S{s�N�_,����YVɄ�� |�J����A�vd�#Iz^W�!��;���DC,�rA�h�Y��3	؉Ill��{�W^ݎ�q�����F�W��/��gC	���`*�f���d\���qYW�a�8Ƈ�x��SZB<�r;���lZ����;r���{NE�S��5FP!����6�X�]�����7_��/��wrD2Q�\RgQk��<e��#O`��!3a�^O��O���hUv��5�W�˗#��|#��
1����f#��`��ٹ#�*��^��Z
h��|��|:b9�^�ՄH�IuM(3��O��>�c~YXF��~#_}��7���_\uo|r�]^0�L� �}���g����>�{lk�a�'�<��ݎ�c������$?�߭v:�R��aN�kY�J�=_�2bPR���\/�$$�-{�o~����7~��>Z���	��	l!�Y�>"�{�oz�{�
I�] ��T���@��n�C��bt�A��?݅�)H=��?	ݮ[��	ǲ`(f��P��OJL�:Mc# #��]�������ϊw���U�`Y��s�|��h���7LP�?�H�LA*�f�ʗ���]^�.�FA�	�_	Q�q&+�p�X3���Wx�2�L6�M��^)=��
�'��k���.Ϻݫ���_���2N��af��(�������Q�؜��Rlx�����t���@Y�f�8���i�a <WȀ)��܉/r�x&�hc����j��.	bur�`_e�}8���`0\��j�LA{
R|R�Ӧ�W㇓�V7�i�k�w_|2>�`8�=���l��'.3@��ej'{<��{}�^�<�"�T�N%�%�BX�����Һt�ޑ�)L�bn��FDKx�L�����E��n������x�����W_;��� vW,ץ�������{�%�p�4���ғ2�b��zZdĖ�*�r@qRL���	�ӈ���XG	8a�b3���K���p[���K�v��iǸ=��pZ�Մqø�X`���g��W�6U��u�����s���1pYAd�27�Պ�`8V��{dZ��P	]Q�����v��!\{(�m�/OC����:�H/����l�1�̰]H~�S]֫rxn򴃿����ҫ��fL �ut^(5�+���na�:OpF>�S��p<���\T�7r��7����-#5XqQ@N��hǩ�~��Ɂ줳`j�k�"a`\�ōOG&� #���	�w����w�)tT��c���7RR��>/0��z�7�����?��̯���u�.��4ݴ|<�s]��zy��BJ$8����x�
�73lo#d�R�ux�5Ο�Q�F�P�$��I� Cj{7R���#
�j���/.�����WN*9Q|���'B釕��H `b���M ��@�v�.�IFIH-4s���R`�3L� 9A��o.����C$�g�PO�����I���W�b��$�^������i�,a��dtH^��$E'}E
Y��vp����\9�>8d.�-Tn�m*��-Lo3�OvSR�l��Lč�cw^���Iq���.���n }x�D4[
N��'I���V;B6����j<c�kTs��՛�v*���ɚ�\6�[o��2bFfr=�l#�m��D����3I�*���HI]g>�m�nc���t`o@Ҫ	��_�ӊ~���7)�o�n��2���#�� ߊ�M�ݳ�	!c��!�	B���މ������](K�Q#���o��>|�{�_����9�.ԳQd]�D{��f�� �X}�ʢmr��O���B���΀	�yh'��?�������r���Kg犾DW�19M��$5�v>�����t�r�I�8O?�G�W�>H�&�zA���g=z��tW���;�R��T�(IĊ�ǀ�(d�J�&�T�������E'�!2��]��Nۘ����h8~򬷧�Sn�s��Rn����]��#Hř(�O�t�??�;l�=�8�P�E*��4,;�5}�i_��Xb*f(���T~Sp���:�!�l\.߹��r`^��6�ȉ���-�z��a0g��N/.D���z���x��k���L��v�X��j S���V�BI�:A҃���xc�	�l]�3�<�8�)l���*���y
����͜�ps+�5�j�����G��$]b:)�w���q��Og!����{ͬ~<�O�rџ��G4p1}�m�Ճ�i?�t����<m�v>��R��ٹ���$��+������/����Od��`o    IDATA;��y�.@�E�3����H�t.�6���`Z"APp�A?ڃ�&�������u��f���������ݤ��br��:�I�Fx�>j�H��s��q2�0�9��o
O�`�l�tŹ_���n��x$����+��Om:I��?��`�׹+Z:4�мhO�Hs��}ڎ�`b}��x<��t �LAL<��~Һ���5�(��ѣGz&�`\%�e����#.
�4�����"��F�K��� 5�c����8QCw�a/��VK�����,��?�CfK��Uڃ��#����?Հ�6��� ��`4:L[�T�sŉ_���ҟ�'��h@� ���E���@���ޅP#�����"���W�Zt���vO��v�Q&쩝�#���)�L��kb n�����Gwx�~1\���L�@�H��W�Py3ĵE'H8�"� &le�Q��>Sۅj��]��J��12��̓� A��G�2
'�n�:����@V,9+�{t���d�4~� H҈#��*6���
&����y��E��zt��f���>��gcl��bv��������p�*�kN]�6&%E�YРt�~ҋ�>�;-_4�I`@�)b��ҋޥq�~�W�H�F��ٕdHa�ѳ��:�:����Z���8y�.--!��z��\�"6�:{����;��H�X�2���.�v|�jI�ZP9�t��])�����ï}���hχ����3�|-�-��3�17�]NRl�Y�M��z���`��=��{�F~5�ZX��#���)*&�F�ZT,EqU�+���+?��?z��m��L{���j*�G�hp!����H�C�D(5H� �"п�_O6��L�9h���3���@��6W�t���v��2xJ���ׄ_��`�RJ�/�²j"�j���Kw���+1
#�����G�����{Uv>|���zh](L���/lU0��{�����^����o|�;9�ߚ���O>^?�����
��rQ-�k�(^>{~~Q�3�D�k�8Z�#Pq��J����L1xv��
{�aU3�R�{9'�;�zSńi�e�j>�YR�0>o��7^��?���+��,n����Y0ؖ;�{ٮ���@����{4��~bAi���Vw��|��P�'1jr%�\8���nO�����*qK����X߈P��'�(����RO�`n!�@�-(��o��,Ӝo�!ǃd%4� 0�P>�`#*��ڥ�٩W>������;�1��B��x��Ա�dѥ�Z�(������s���6�l� v�W{&���Y���`9� �
ܳ�ӽ�G�j���p'[:�m�[�����]�"����/�|g���'[~�L$:X��ַg��6b�J��f�k���|1�*cf�	�b�mC~��'��
I��Qc���<��GBPrk�߽����S�,D
$L��l~���#)Q+���ӫ'� U�'wK�j�+�w���`5�3<Ñ���һ���d���޷����{/=O����#�Xz/C瀢��s���V�xp��3vW�{3��h( C>|�!5����5ݹR�j��*ڱ��<ZBp��q���\�g�R�֯������v{-k�l:�@C�fY{��R�/�L�21�\�.��/�EսL�Cj�]ِܑ_,�JP�xH���ГG.��2%�~5CR��)V2_����IF|L��[Y}��g�O�_jFE�M'���Z#[^3	�7��PY֒��͝[�y��wۇ������+?W^�ب &s)-��a���NVd�����s2t%��'aQ[���̼�TD�1�"	����id�f�F�6����@���`���������B5U/��L�|��-4��^(Ey!IB�NNa��>�R��;.�J�e0����<�YYz�`�����?ۀ�m�4�쿀3����{]�K�|
v�yJ�I�mM����7�>���盩,��$��9ҥ����CfTV�p1يG�Yd�ɣ��UUE�Vݺ��Ȋ:果c:ߌ����6A-:=�;&�l�m�@�lɱ-[te��`2�,q�ǁ#J���s9��F"�٭/�;�����W�����W�gZ��&Q+� ���!�k�����U���b��� 2P�x���Έނ��u7�S�7�X�-������]$j����XIc�a�x�P�(���z8�x��Y縃��䡚��?4.z��ߋ_�U٩�����6���?���wP�|���W�F�46L~��p�E���r�c�SIf�]9���td0K,�{��9ޜ��ٮԂ:��������!�X���+�J�Q���g�/��W~�_��ln�S)�1)^�<�$��w)�w
Jz���VS^B����'���d��f��^�A��PvV�%/Bx����r[ߡ�E@
������$��|�D�'����\Q��e��ܓ���A!�MD���������;5����ˋ|��o|�[���ͪK�[�ኛ+y)'4���@Ȝ@y9����QL3���&6��K���t;m��*�'x��s�Y{6 �H�j�Y.�$�w|���h��_�ڻw�v2��\0�I��V��r�&Hދ���VK�\�ը�2��fo@ݲ+N�3:�i�k��w�8_��/C_ ��ӵ�T��d'/��0&7��m{mA�cn>�ί���{�=u��c�V3��i��
�e&�e��#�Mm����T����<��[>�֛��_lX�%�,f8�p�%(!�Ƽ�R��s=�ֵ�
ݸ�Hm�g��O�N�X,�iS]f�>���)��n�>�'���浳�Ĳ[-M����u�y�W�T�q�31�O�ȅ,��2
n� �n�L|Y��Z62[�yq 7�6�0v��mK2$n�t��<�_��̃��u���~5#���$NevPJ^�(S���z�Js �l(���!S,A��$"0?�!r����I��R�+�[�?oe������U�*��Yd{��_����^�Qe��o��v���#����	��!ry��p?
Y��R�A�W�u����0�`	�W�J,_��"�`8�N:��o����k�Q�k4d3���,�Q1_#q�}��I��p,nb���������r�@�׈�L��:l/�{�i�!C
v��;d`�OT�EXT(�����gh�Bt��A�k���Aa�2?���,nV5/N/�o\�և�#^	QJ�ǌ�"�}��Ea3�<�ݺ��5
�Khu^/5*�����e��2��]_�ޭu:U$��R�EIL��Y�U%^���q���n�E.�t2��9W9�+H�^��2G����,gQaZ����o����Sl�o�=a\KRZb,�$ 20�s��Y���� >�;X�]Bq-�q�ȍ`W�)�A�'���< k�e�dn�	x�u��2R�V���v��(s�a���#��� 6�˹}ܸww|�p1|�f%�rWt[o���%5��4;����A0��d~�x���q��/����W~���o�4���<�&/y��U�C��R��뜊,t3�if�n���Fro�YM�[�D������}^��j	�bw'N�_�lt��@���V����7����.���r���/���j�<�n-^Φ��@~�{DLTD��M���zN>�YI�-Tq����ͷ߸���n�J�����r ��]�������_��ӪD^"{Y9�t�r���]��doӠ{�J��~3qV0pF��0̎��R�Ӹ�8��wk�������,��I[���$��Ն��n����fo�A3����a�N(V:5�rXavE����|d���h4�|�b,�<��*n%�F&Lp��wWA�_�/��F�����f��=ϨK:^KJ&1�C
�P��吖%?��pY$�G��R5��3�IoQ��<��JBfA����b��&X���G 0|PݥtPC/����n:r\��� ���)Sr0�����D^O'�Ȓ4�@i+��"�ldZ���Ε��;^l!�C���!��;�+�k��i��d{���JCčbc��F�g�τeJ.�#01)�g�����)��X�7���}�y�"�fX��������r�хS̢Ru��dd@�"fa
�K�]fDL�P���_LI���=,���>��@���Ҍ�2����2��VH��V��vZ�e��c]�F��.k+}�u謹8<X��d�w�w��q��%���Һ�R��}x����~�+����ϯ`�Q*�1k99�	��%'֨�U�ISA�U�W,j>"l�"i� k�Q
5�̥�X�m�Ђ%��]<�M���ˌڽ�M� r2 Ӈ���6jvL^.T��n�^�%���0<�	)p�|>�6>__���"/�������b�Gj#����I{6fLh#��@�DTwڣ�iK����N���Vi�j+�沿J�uk/_W�����m3�$�.-MsG4�����Ճ��k��T��r�P��,�[�d��RN̥*w��M���7mȊ2d	����oVPg������ڌ=4�,`s~%�Y��T�L:Q�W���Z�V�BM�*ݭ�f��=.���+���n�>�i2x��| �,roce����,ܼ۬x��������� �_[d�
N1�Z��T��pN��^L�΋g���6��, u�I:/Hz�O:/Zz�[z�W';�?�+.j������{Љ?�z� ��c��-#�+��I��Ŵ7͜��փ�����[�r�/�l��+�d�߃~5v�I:*��wu����u��P9�����6$A9�_\�A�NގFӭ{|xd�D���|5�Us�����0)K��̖r���O00oL?ىè��p}�v4�t
���6.:I?3���̦�u��=��?=��u݉��.z6p�����٤�DS��y�#"��&����[:Ig����c`�'L~���wW�:���E�|��x饗~��3,[nܸ�V�Tj5�Z��t�'GGG�2�u��ɓ'��FºI���u+�޺uK�ZZŧO��5�3�{�����\�y;���믿�ϟ?7�%>@��г/��ԡ��g:������4>�A*=5���ĭ����d䁯���#х�w� �"�!���t,�~0C�RjL$��9J�HkYE ���v�;,�q\��x �SxH�ںP⊪A#��I�{c4E.j��)s��s%�m�(�օL����a�����㳯��A�,�6`�Q�p�U/�'�������h��`�mOD�c�bܷ%K�V�Mv2]\]>:����GO���1mv/��yY�f�n����}��t8�|n��xq��f:.��g�M����j�ӧ�fn��&�0�i���X�N�M��ޑ^�� ]w������SLK;wş�i{{{��)6��"��i�^������0d[�̕�� W�-��_�R�E��h�]@O-�o�S�xw�o��]�3xm����nv�^��YV��Ƹ֨�DH�6�g2��S"c؁O'���]�wd��Ƙ*�fo����a�YW�|��`�U���U�F����������lvw�y��z:c,@��`DFc�4�h��'���^w����)�R���p'�(���p���B�|p:G&AA�V�l��b�A�'YL:d-@�`pT���堨ư��tfm�H2T�wٱ,�%gl�C)���l��.)��ds���i�O��l�����kV5_l��W_�U�d �s6dk����/�2\p`g��XF��P�3̈́#�A���fR,��E�H�Z��a�ɚ
+��-�ɽ���/��w��Fn���]?�Ť�# ����'�a���tO	 �>y>����r��dE��)5�:��:���%�	ᓩƪe�^��d|�����Ku��D<�b�K����x(�#_b֒�]�M�!�*X*���a���oG��"�*OL���R[~jE�|H/����Hfn���v}��řW� a��_��"�<m�C���:�'��e��xN��D��.yE���bh��DDJܡ:�,�t%D�"�G��lu�����V�Z�����/���ڭ�Rq����Ř��yR� �����,"8�\u����?��߾ߝ�y�PWq���J@&m X^%a�K�X�n(�o�6���M�G���
Y�Qq{bo�k�a�Q�u5��?�tϸ�R�	���JQF�F��]B �+�4F<t�ڌQ?�6t��oڔ+��m��������p�QU(���K�x�+%d1>Y�r���n6�*�F�S\��tr]�P�X����|$�iԹ8���,GR�%��ޚ<N���������ļ����ˋ�����Rc]أ���JH	V�u���_<��̔/�x�e��{K�ґ8p�CO q�A�vk�A����1H�p��Ce-Q���>��j!tF�_���ZC�C0�" 20�p������:��=Q��4@��wv��[�Y���dQZ�fRTc2̄��K,����3����e#����㼾]S����Ʉ�}I�:��`']�Ҁ����k��B�M	%)sn��e����w�����d�lz�ˡ�2b�YQ"��Xy���qۧ}�����}1�~����{?y2I�{�"��0abZ��coD���(���!`@��r
!I#�dA�?���)��:n���Vd���P�%%qZm���`a�[�O�������Bl=熲I��Z�����ۏG�f�ivh陖�))7���ۊȏ�P��5#r*Ӡ���4��0�X��:װJ�^o�ȴ�J���BWf�3߼r�i����z=(t�Ϳ��~���.�������u�)���}%�9����7�Ǐ�?���\��Z=a3�	'O%�=�<�S�#��/�v޲����C���|KL
>vͲ�/��kF.8.�FY�
^�m!�5 � 
�	5~Bꂕ�&pU�G-�f�`[mmg��6��Pr$nC٤>�0��e����b$��ӟT<��l���e�(��؀�tgr.�p)� ��݉�^a~2~�������j��]��������[�nd�"�/��X�"��z-V"��1�ְ��jQ�U������'�ȥ�BL�Sn�!�)o|zf�[ێ|?�$,.|9�Ԥ ���THI���G��2��xup�������� �5��O��e���!7�<��e�(TX^kyvܣz���;��^~]X�k�F1����qc��c1��
�OU��
xR������)�x�M5t2�(շ�zM`���l�X�`.�A�"a!y.�dE�LV彯�?�~�䦨��]�&�H?+><�Q�%σ�Dp�k�?w�y���?���G��W���f{YC
6uZ��j�����ߠ�e�AK���Hm~a,����-��Ř�$�V�� �9	���Ѿy�H�R~����˦�'��FLLD�gK������V�:t�7O���oY��)�l�E��D���nvv���h8��t�>����/}J�PaHd�ܩ�����w��n4[{V e/B(�Vȫ�1|����*��w}��[?����zw���lƛ����J��kYg�P�9�
���pe2,�g�1B K�;� ��DN	ڐ�٠�0s�a��د������y�a)�����1�1�Z�Y�K�#?��+2��l�6�}̌�`cvhn9L����>΀�������Â�>����CNlȉʭ�ܨ2ݕ�M�*�ł�p�2�s���+e#�3pFYYKC�U��*�q0�������`(��T��Q������Ϳ���WW��r]���Bg ��P"=6�D��kd��t���<�7?���9��7��(�lW5�F;;�:�B:#)l]g/���|U�ϐ p%�~���a�@ �'�SWݶ��I3	�O��!�@���	����	�F
������r���_{u7s=}2��sl�t�Jp-���\��v�IMl�D�(�)��)>��@ԣ� dg|=8��j)��^16Ov�yF��R�(F�`_�A)����o����ů�c3�������,,��pp�1�ة�<,e�(�ht?��ٟ��'��)�L������䥗_&�'3������  ��o����?���1�6+��{��ŝ�    IDAT�V��_kV�/I|Y3r�[��w&�˳�� ��.WOřJ�]�~|�H�a�3Ro��Ӫ�W2�f3��I��b��^���a+1n܈�ݪ��; ��'p�ܐ�&>Uo��D��B�q�!#��B��v/�d�Ђ;�42Y���=� �ӽ��I{2���5F
�ǖ�����w#��]�����8
'�0{V�Z<�Iv$/��m2~����jSU���L����y�Փ���Tn��F�'���>��N!��ٳ�����H4�A:��I���OB�\1�H|�$��W��t|��"׿Ĺ?���j�a�������`ԣ��N���t�ˇg�4�.tw�b�ƣx:���C�~�J�Y�����Q�Yo?~���A0�>�z�^��$V*�H�zF��,3�ׅ��<���2�2)�W���6���:j���ڝ����暻\B3+{���WT�"R��`^����:���>|��da�(U�N�;��F3�G
+���4��a���H/BHd0	�HD+��7��Г��pX�c����O�l�X�p� ,z:L������I�$_���B����W���7�	�D�A��x���270��(�r߸/�ݖ&6N~>�3�]pD~�i�L*�- 9��="J��썅�O�q}5|�����tG�j���e����֗����v�����f:6F�a� $��Q�=�!���R	�I���O��%讆�4�#��|a��"N)Q����O�lT<	��4�� ��b��-Y�� �K���qY!����t��m�rؠ�~LC�B��� ���Q+�a4w+�݇�������(���ߒ�_���P��ocl{�c�,6����a;&X6;��xv��z{�Ɔ9�$1���U���ߛ0����JEi��S�lw�ջM���_��~���V-'�Q�4�ߓ��@�8`�����I2gF珇~,Ic��n�Vk(�}�(�l�Ct�6��OJ:�r�3���>�b�g8����I�����:k� �+OE���NP�d�:�:�R���(^V}���vq}��G���Cm�l�Q">
�~ћV�yxx��3�a<��20�EW�V�zx�W�P�h�9 �h1�$�)X��׃����/2`+���@,9]�%/�	-����J����������ޗ���l0_=��Ș�p0�+���L��H;v?y�ч�FSI8��,..P27C�m3"॔Y� &) �tR\q��0���'��E`� ������ Z�jE3O�܃���]/~?�2�b�O�t�^[��3�$�<^ڛ��|� �!}���h�܃��G\q��z�6�-'i���[���#�'m�>K~y�ɮ�8ҋqŹ7��zWz�\8��uѡqz������������]�f�x��W�'��,җ:w�a���~����6Z��Yz+�N:O���u������#����8qŹ#E������حtr�[�%5}֯�)n��EǞ�T�w��'���K;���g��q��11��G�Ȩɾ�7�G-���ǟ<yBD2FM����o�-tW�۷o��Ǐ+ۙ�.�6�y��8�Z�5u8q�h:����޽���o���F�M������b r�[�ܹ�k�<e
��	NטG���һ��ڋ��a�7z�\I�du��d����!�{���d:���?{f[��ja4
����>����+!ֽnw�z���}i����Ɖ�3CJ�䂺õ�n���6 }�M7Q��]����K��S^�2f2Y'D(�
����݈����u	�W��0��V��V&�N1��|�����/��od�}[�a��ȎK���@�a�ʨ�z~ѻ���Ï�?x����ય0�झ�6V+�)^��W��k��-�����f!���|NL\:w�-O��~��Tz%������w]��-~�W��ʳ��bڛs����\L�����7�{��ЊJ��?�GzKK��p�����)s$�do�+�T���һd�&�z"�F�VS�Vئ�d@�z�٨�Հ�m��������ZÞX�ii�'j8Q'���d8�V\�}rԲ�c�䥋���0U�e��RD⬪z�h?&�˥������9�=X��{���֏��?�/�~��;ۚm��mX�	��)���Wi��Ka*�r>�������gә����{�i6[���k( �b!���B�tJµ�$К���:uq�^�)
|lC���dA'�4�n)��O��kX�c�K�[h�K5A�� {,o�G�VV@^~�`�(!K7���v�P�{�~0����;���~��aAR�<����>Xf�����UF�����q/"4[a��lR�0��ewXj	͘Z�=< oHiߤ�sF`oV��~�������_�2ٮ/gϮ������<���ҝ@�A�7>���U���/�h|EDV�
︖�o��;�ܸwx�]n��s�D5�D$j����\����.��sD��v;B��z�� 	�F�7=q�dYEL�h �Ԓn���k%�?BS�1{{tT�*R���I"{=}Z)����om|5��φ䕄@E�d�1�D�=9i�mQr>#����f[|C�XR#k٢��#n,�������a�3*S(����]1�������Ϋ�{#������'�!k7�t�	��B���^m#�����g�3W���4J�!2�!��*�������<	���R��k)+��l���ZY�K(Q���( -^4�����p�C#^S�/�2������A8��R�b�����<^��j������L�+�ճ�տ=of��d�s	bYKߦ}GnY������jr�|@�E3ί5݈p�^O�U(ex �q
3O��-�ޓݩ+ʸ��iM��V@/����������Գ�ӳOF����pq��#$�]3�Һ��Y�n_��?Y|���N.Rc��
��/���$Dݒ� %#f�����g?�&=Hw]�*Y<�c",ڛ��.��)�	vO��lD��7!�ԪV�O��3�O�<u&�y�D;mBm���媶�y��[�r�xQ[��BWzO�|iF���I%

�B@E��lCx,!�V!�'F"$�)_�9�jIA&����3����[&+j�c�����_�k��)H`.�h/3̨ؗݴ���`��27��?��1/�$6�����z=!]�^)��^�� ��c�~��X5ԛ��c�Wh�%8�0]���������xJ�V��80BK�4-�6���VpXX�P�%���R+�΅)w�-����\v~q�/�݋�#�L�3��� �lpp��kH�>,�����2V�0�D�W�_W5���Q�z� m��v�N��hQ$�CE���W��K�l��������'��+_��6��?�������Ap�R"����VIװ������e����|x9�j�R��T�Hb�Hv�H �� $��)EH�m� ��؞���J�k	kI�� !��CuL���`EZ���K�d�@�xĚ@�0���t�B*7������[���a�?}6fb�ȓ���w[�}D]0�t�%�U�M���f�QSoX�[���
/"? ������!g�1A[ӂ�3{���z������~���������g�)�H8`��E�Mm��;��"�]�!ќ�����/���!�Ȑ3ä'I����~��]TU�ZF��`���ل����"�	r����"�H�'�$a�-�`�����bo�HU�B	��ZHa	�#Ռh����pZ�b�E2��"3.�f��UI�մ��?���R؟�#<�U�����,f����~�^f�G�+e�KU`^��i!��#tC�Wu�Ye`�x��づ���b��[o�����[��&jz��t%]�Z�/���@&���A��E�����?}�ӏ��ے�L{A�|ݽ>���q�.�'-��P�N��qJC�����	?�t���>���1Q6�l^�դ�%B�vya�E!�  ��_�P��0�[(�(d����'��?��O�6��~Z��q0.̢��A��ȁ���ʎ䅢��B��urtrs�xO�|��M#e�2�]�$��}1�:,���g=)�������0s����^������F6sog}6;�`r�XŦ�|;ۨ���	N�U0��è��P��F�t��_�Q�5s��8�_m�t&�4p����%QƮ��c[�{!����;</&�!Ϗ�]F��<�v�����ϞҪ)��E�`�����z���'|-�o&ن���f����ށ䨥~(`mn[���}�(4���	D���6�'����i�r	���H1���DM�NAw�ڍ�z��^����+��lv��>w�,����Ƽ�*"}����/X1�JM����G����?��ӟq��dWn`���Aխ�ׇX�8`�A쇉 O�O�^hl6�**��y����؊�z��<��{�wQ���%���޸?��7��*m�Z�7RxE� P^�ðe����y��l�x�-9d��׳kN�U`�df���G�Vp��Q8L.sH��ډ<+����k��m� UH�{��~x'`��e����las���z�(w�HS�J�����_�����m�N.���l=�z}b��I�GB�!!�:[��ѽ�^^��ٓ�XyXdw@�,�'OnܠG���;@��%A��\����O������'j/f�I�կVh��	�&��,�\��-Z[�[�F�.'0�-�ɢi�'G�ԫay��3���+%�UƔ�� �J2�̲춊�;��F#�<ۓ�]גrJ"��0{)d�SE�$%dd$�P�nw�IWK����'�1(2�ٙ}�7B2�i�+e��h����٨�D��x�_�]��|����w3��L��3x<�~>IJ�B�W�:�7GM�E#BT�''��g�>�p|�^F�c>�;_|���n�Lsp��������N���>}��FX ((K�'"/�	2�ڧ$�9������jz��xh�&u�=������X��.��
�	�����[�l��F��������ְ*��3��x�s�+��Tv@�3�H}H���r�G8�d4�U�X�D�i����9J�鵸
�6P��#B;9t���lؗ���ۦ^��~�o}�u��Jl��R�D6|����R��R�WcGJ�����~�������c;�j
��"�斄�h��ڽ�Hcz	����f�"�( Mfl�>��є���1ǻ˘�+�89�L���6:t@���A�T�B�3�<>�4�D_[�ɣw����T�6� ��.S��1�)��TlI�$��L.��ͶQ\xq�Ш�vQ ����c����&K������T��J�Ķx\��j7dx�_z���Y6{C��z؟�.��s���%�~�+���cU���4���dS�K<HSc��sp=�j���A��\se.͑�� @����$�<ހ?�A��I<�`e��	u����Fs�:�1[s��O15�ńjY��+h���ja��~"C�O(�p�]�`�U�)>�^��p�&#>TR[U��:�F��*���j�x��� 
�+nd��&�&���l X2
��b�>;��[��ޮ�=w�����<����t�ʙ��r|u>Ek|F��}G !3��X�H��>���_<��
T�i�P�%$q���mD��{q���#@3�/B%p�f�]���x�u pP��e{w��ɾ����>D��}0�/"l���,�Yʃ��l�}���|"�Z�~�9!���׀㙕���� uxi�0.��+��d�I�2fx�A R4 `�`���
��`q��m��Pu�Y�wr��k{�?����/q��^].����x��\�
�} ;�]ǻ%�A�X��Q�����.n�#b�����tD����H����Su_]�-ׁ�3�*�*MeV�o{��Z�8� � ��Ar�0�!5k�K���0z���Л���(�I3Z"���ۦڔw�3+�2���6��ݧOƉ'Ύ;vl�Qi� Q�Q �f�R���a�g��d�lL��A����*8g�(u#�u(qvˑL���돟Zv��:�o�JϦjw9;\���Ծ�����ӒT�ݧ5�+`c�Д�w�𸷤F��k����=oIb�T���t$ґ���Y�8�W��u?4J��Mi?UpV�[jzD#.𖱌f���lj?��w�g%q�Nzcj�7z�KӋ����T3=��;���J/M�=�ޫqמJ��B����R��^��z�:T��`��w�FZ��x*A���"����x��)/)5�f(8��H}g�N?]k�u���+<�����;w���(d0�e�)�c��z��y�ƕU�vvhԵ���vqB?��O=z�<�h��'Ť:��BOB-xD���J]t�ߖTz饗@�{�)�^�x<u�=}�m�1'��Л�X2d3ر�sM9����f���b�Y�rd��iDCs�?9�X���!�$��5	
B��1P0)Bo� ��C^�M�M\h���dh�2)�����z{Y�T���.�6�ɼc��z�tF����5�KI6�Y�=4�M;'��v"|�6P�Ԋ ��ay�y
Lj_�@9��|��û�w�n�=|rpt��g=ᗉh���H5�Y O#�"�}��X����3��3h�ʾ�顦jp �$d5�Z0��x�a|�+��R	Tt7��S
]�����ʪy�:I�hʇ�y�[�)w�tW������V@5{���^-hG?�=;�~�І�O;ͭA񈨀��5(���9QM�Qʣ&LLq��#7��_+�?_}��ƍ�gpb����E(. JDl�f�(eI��ӕ����iG>6c��������f�N,���A��޾��C*����խ:-emu�;�_����)��;�ݳN|�ot�5�0	h��)@D��y�|k�wLɟ�����}��g���aU(9�/�*�;9pa�u6��ґ�mLs�>���X��M�3lo�k�m З4F�5Vs$N����3�&0c�MܠMCRry����Pv���V��6.S1��rF���NT�#�ߐNC�Fp��Ҵ���R�oV�]VH`=�IB�9�K�M�,_KĦ�[�SJ�z����g>����b��5kֺ?�y��C+X�x�)�:L�"�^�;:>l=��Û�F������v��W�mܼ�µ�k5��1�;[�����9fPz���7o�;�m�u�c���,!&7˰Y�l�����H��d�qbB��V��\�Z�Mui�2S;��^N؜}H��j��<7][�YX|u������ӽb����pѿ�f��D�"�E��*���+k+͍�A�f��R�����n���ݐ��k�S�5#q��\��g\��G��_���_d':�x�߹7<�G�N��%b�֡]�'ќH�;ó�����igZfg4ӧ��+��cHZ�_��[l�@\hM�B��;����Hy�'����ˆz� �7�F��#�q	�λ$�S(4�@�u�~�O�U��e[>�`k�M���	��I�M��2/�b���.�7�~^8�F5֤B$ٔ5jKEJ���3�g�㳽ݝ~�+�����
K�Q����;���<T��dzz�E����?��=K�2���to.Vu�r냿���|yn~5�F�ϞlZm��= �V�ER!��Lg����=��G�����$�K����j���X�E�ѬŪ���{]��hb�����H�O��D���DjTs$��c��c�~ �c�VE� �ۢ{<�FX_���#1@b�v�r>��&?��76V���X�\�_�X���Ӈ��yQ��̍�"�����SSt����I�	�ʔ�<cO�����k���N�/B萮ȋ��(���pqV���^��w�<_�Plyƻ�ӝ����e3�&�lt3�c}�+�i�msE��?>�w���������m@�R�`��YV9�?!&����zs% '��
�F$��B�~�w��5mgn��E�|�b��]����&��9��,�U�b�@*��Ml� SO�1z &�#�|�ś���v/Q#-'@$_&O���S4b\�3r�	|Uc>8P�8W�$��r+�����{C��G��G�#�X���_�Ĉa��������W^T��    IDAT��K��;ã}��k��H�J��լ��A,�������{���[ݚY�,?�9|E��NPJ�Y9��U��Ȓ��ͦ9�@H�cy_,�DDĤ���m�M脰����}V&�~QL�Y���hY��C��XYG��b-�BK�gO���p�6�\,��I7��rYU��Gg���@�Y9��j��O#})�?K"�� b4P����h��� 1R>g�a��O�3�[�������_.ן�j��;���,���
�^�uR���e�i��?�������(Q�6�;�[BA�ʺC�%�Y���ZK�݋��a�Û3r�����VM��� C�:Q��X&�5(Ь�Lm�JI,�v?F�IB"�N���c=�c0�aD��jzb��곳�++[Ϯ�޼8���e��yi8twϺ�{V<cF7u�%����� tϢ��6'�̘("�5so	3�����s��un�����O�b*���Օ�~���|�[����ǳnkt��#�q:O���:�R�}��Z#�6���у��_�N�����-2��Vd4f!��q$y2�YAi])5]'x:g�~W �1"���)�'�:�Xz�t�c�E�qĩ�F�KA#�?���s�{S!l:l����ԙM)�p�����)����@�潇]A
8��JӁ���d�㍣���ʶ��m|~�i���z��N��+e�G^Q�G_ 4����������e��47/_��+_e����|������pO�+&�(xGl��Xq[T�� vCV:�����sN�����X�1�����P'"�ع ~P�wi��e������c�D9�4��Ɗ[="��4ۅ���G�zu�OW��]&�Q��dl���M1݆��ҭn	v��?'��z�\�Y��R�{Rp#�]X\�b�T��;�ۡ����\�m�w��R����WkeA& 91��w1l���mT덥�p�G{grϾ���	m��o�巧+�g�P�Y��4f�����ulNH ��B�<q-������7��O��E�n4M�@�_���iZ�-F'Q����g� ��+�\6q�دȦMd^>1;���12.u����q��C��騺4��Z	�`O���78\��Q��I>�+fϡo��sի�+׮n��Jl%	 �ZdϰRoo�1�9Xk>UPH�����'f�`�pE:���䎯s�|����,˝�=�5�4+����/	�
�$_]������������ �P�����>�EQF<QH�4/
��y�฽w|v���������p8��޸����[���ʘ����J�����7~�t斲҆�H�C���X��%�C�M��+촽@�e |f���v7ׯ6W��D�C��g�i���
�Q�G�+�\yU[���Ǿ2$��X�1�a�s>4�x�A[ E�,�������)�;?Wk�)Z�@�s(g�1��~%��tG<��U#��3\���Ln�-m4�^[���Ya��5׻����	����x����
h�� �(�p�x����w�#[[v�H���ڳ7��r�zmĦ׼��<�޽K���$��D4�u�-Aơ=r��_�[���ؼS�3�������&�2ű� ��LH���jѵ
V�@TZ��<?߼^�z}y��郳i?/ ��VK�G�#���i��(?��M+]e!��T��hF���pҵ���CK�`����i���	�y^�CV;�耳a��e_��b��_.6$������N�p9�W�u8���KXt�1V_�İ7h�{k������kV�L��bfk�) |
1��/𨖉�Q����(������x	/�@Ĉ��":7I7��K<���q����(�*�)��F����˴���ظ|��|��nuT�6�1��Ŧ�0;=#�
�"��|��Zcyg��WÐ�"�=�'����@nM_���U��pџ���_B\s����py�)��?���������������&O��	-���c�o��$E�8:�u�Dh�������x�7���zA��5���X���(B�{���K�]UD�P�#{��/�y� ^عI��c���U�S
���l���:ᴁ�r�ݒOP�h���QF���ue�Zn
rz����>蜅�v_6�DEb!�
�F�f�M�����gH���F14��׹�tz�Bvx!D�T�W�db�-m�4!r(�` Ѷ;'W� ���S�_��O����u�M�ڏ�i�4[�e��zl7r4y�#�����v���f�S���ޫ
!s�3�uqV�]��j
S��{��`�P�l�����i����43������Jh�!kV���,���ܢ�67�K��rmi��x|�r�;>89��;�[�X"��F	&��vL���k6�/��.6��'�I	!`1_�ؼzN��׷�7��7HBB-����=��B���NW���ˍI����|�֧>9���;���v��'��R>�O��,3=ۣ���~��'�Ҧ��݋�ł��A�ɘ�F��8�]���tdw�Vpv�u�~:'*��q5���O���?�ή�AL�~�ДB-`8��Ԭ�1ƙ�P�*��ZVߑjz�|^�Ԛ����Q;+�H:�Tӡ�t���ש�ޛIoLߞz��R}5���:��q��g���=)TM5S���ޢ0��>'���;�_��Å.y��.,��R��.�'�@Z�Uv��.R�N}�:\{$���:��Ѿ���E��GR��FTv���Z�t�0P�/rNL�]�H��e/�'r�L��C0�x� �zС)��|�嗽B�ނ�N-h*vu�^���V=��K��^���9i�(5���u���֭[s���獇Ë��Ú�K>�����i�E��S����T�Is�!��$�G�L�*{�vޚ`�+���S��g{�.�Ka{��U�zV;*�$����(���:�w�-�����@cd,�!S��>�O�'����5l�_z�<�M0]���hn@��И/�	�e��7@_�,F��
�&��#*��Gb9�aC�݆%�'�k�%� �ɓc���,҃�5y%:�.'�yü���m�X�p�	�#�`�?�8�i-�����ف��6���Q0i0뤦C�F3K����w����>x�std�I��mY���slvp+�j6��5ޝ�� �[R!tTg�h�ġ�
Zs�v��Y�id�W�-�Su��0�׈��M%��g�S�ew���Q�~j'�Q�P?�/� ��4uϋ�TG���󕫟�>�֠`i�ѥJ�L�ll�Wֈ�t_a��l͂��"dm�b|��&�\/�Ҝܠr���|����!�P��-ha�]���%0��l��<��q�;��-ҟ��"6�M�%Lc�5�hwf��j������KK0���������O���N��<x�l���z��qR4����n���a��s�<>�i���)�XSQ���-ͫW�\�v�	BAp�Ѩ"
!��|���!sW�t�y���HZ��5��A��uf�JNL3���ho�>����>&�2Ǎs�a�
���}��x�ê` ���6==��?�%i���_�a��f����t��Ң�)�b~Yd�E�iyKk��rz�\'�^V���p	�-�V/�N�Ļ���b�VbL�^(�=-���;_��?���(.�����ڇp�Ե;7� �]<ko�h��	�'o?x�����\��&,r���4-^{�S{��+/���E���3	� �h������~���^�m$V��,00D��P�C�6�Oh��IZ2��d4��h�R=�ӰG�ػ��2��-��B���ZZ�2^�$5����or?]d.��'�e-M}��`̄�
]a$���`q�?'��#��}� %F�C##O�)P�I5"@^����9��p�m���[�����o4�
�����ѣaO������G<Ha$Bi��**�`p4nv�L�>��D�����<l�L�X�,�2\��u0��F��?�/%2��^S�_�.":�Ml
rA�B��]&7��Fs�z�?���|	
�n�1MwIH;�����m�U8��D [�`�����Ӫ�\&P��>W�da����*�.����y��%��݅<�N��R�e���;[m>���,���֓�i4�0�k���X��3�8�]!�K�\�χ��[��&�Ec��?��kשK����㻽Ó0��Z�ZF��f�$e�ꛪ��%6�u��<�śg;4]��wZ���Fsc���+�j����}�`�����
A�X �IALM���(^P�����h!Æ
�p��nes�$�I��$?T�jj���+�Ь�H�����.Jr̪���W����wWǝ�3�"�y��.�~I
���
4�x��G�>RA��'<.j����\5��a?2�vY���խ������9d����'��ڗ��+sF.�ޘ�G'D�X��)#<��o��&/���gǏ�~�No"#��2*`��&�0�6�DsF��E
YJvr�Lt�! rm�0ޢqe��l�?̖܌+��@qZ��DΟY./"���l8��Y:i-����YK@���zm�zqn-X��Ҡ��P˟��}T>א�K�Q�����Pd�ܨ6�<s�e^8������B�������s��M���'����Fb�9N�Uz������s_����M���^w��1�i�d3�>��<�@�8��e�Eo$����ѣ�֣���(��e�N�4�c���9a5���`$.;��m3�X������ļ���K&�8*@�CQ�������0�A��s�[�6)�Z�"W��~�7��d�n�q!+�7��9����/J��R�7κ6fh�$�������.a��i����0t:�~��9�&}�_,S/��h�6$~���W�pVc ",�X/"�ի���?�U}������h|�Dϴ�����eM���4�*�We2i����������)��"!O,P��K����,�Y�p.�	2`��ɴ��7(��^%��x9'$7R�X(�fH�R�T���˗�����7)&��$�A����ðx�\����Yek}��?W;K�I��$�r�C��ؘSF���`Q�_��z�^�f���ޘБ���d���,���i�`kb�N;���I�0��1��}�5>��|�_��]ϋ�y�?<|�;��< X�M�8�L$p�`��B��n�u��;�G���[�b$NB�a_�K���&,h��2"dV�{ ��Sґ&��(j���~� ±]0Z�7�)���N�O�P�UY��*��}�A��쌙�aD\��(	��	힯l��]\����٥�f"�A5����.������ĕ�����6�����q����6���fv���CC,e����G�{�Y��jbf��E�._{��/�ŏ/?h4ٞ�m��9��!�Oi�Ρ&Kuw|j��qT�)߽{׆׷؆ n�J-�v��ʁNM�y DITVW��I���[	۝q� ~F����_u�gl֥������k���N�i&�RZ�����i��Pʩ�@J�Wr��7�7.�,tJ��m�e����с��L;�T�bϟB�Wf	�
5|m�B�M!���.Z�Z��X)��b���N��ly~rk�)@�Ƴ���o�?]�Rd��Ξ��o�s�o*�<j��K���y�!Dp��A�ɝ���w{ ��ʹ��B�9Jl-���7����7H9�@5�9�.�IPlK�
���qɐ=0o&�k���Ƣ������7ε�g��uyimC�װ��X����B:�2D�,6�D��5�Vr%!s9tO�_�'�q�����cć���͕�˫V�y3����{�y��Џ����eK��2���������?7l�N��׊K�Yi������W�[�ɳ��������|Qx5ҋ2�q�q]ex�'<����}k�i�);�&x�R2#QER Ia�-
rJw�P惖v|i����zW�����G�-.�z�/�&1�j2�ـb��+�
�b�I�M���8ϲ�3aNp�6A,d5�V����W�ؼQ���|7�2L�����|�BQ�iN�]f��bOs�퐹	��w�š	
�������;���'��HZ4�ϸ�?�l\�p�����ai���3�]���'�N+>���u�_��vNX-�t-"��vO;���t4�O�X�N'����W_z���rU�<�)���#Y
[$�޽{�u�%�O�1,J=AL�I���(��(傶Q��!�D���H�X���(a�q��oY�.��ƶ�s�����Ë��d��x" -"�C$s"�-F���]���;`8�B9���u$ki4Se������q��O��f��
�!`��Ϭ,oUVG��7��w��/�8+�ԣ8h
�i
��!�
�_�5�!L���eO����7�<���\�H��#���f��b�i0t�^�48q��8�~bDlC�2K���(��f�m6|�:u��f?K�>�#ō��1�Kp8������K���y�Q�JW�5Z�݇o�vx��%��/-U��I�s��	�j��Z�V1ŅE%r�����ܾ�a!W��Q*G@�p)3�g�B�Rsqщh|R�$��O���x�E��T�z��W��O�Ć<w88|�9�=>��D@��B��g��b��(r��s��7~��#1��a�87��S��b,Mb�An`O�2S4�3��F��`�p+E-	~6���,lҦ�)N�}��pkkckm����2�=�ak�h�0WS̎����f}e�֋�)����!Q'bY����fms}1�p�����|��������홉]!�P��np�N*rqz�Z��l���>t^m
 ͘�٬K~P-I,���g���K_�����v��mk����D�W�����(i�/�˥u����nw��T��Р�&�o5�ъ@�l�t�Hh�" $��gu�GP��O �`��bJ� 憈	��7�Q��M�҇�I|����j���s. p��n/ן��c);��$�	���0����W~�0�0e��q�:�s�+�L6��C�rĕ��{fZ%Y�p.��"G[�2�<s<�Q��Uk��_�����蛳����g����#�O5$�*�����K%�ѝ�ѝ;���QY��3��������M��f���W��<#��o��JTN�wz��p�Zs�����A���f����UPd?s
􈚩�t�ZgR���tK��.ҁ�Ҿ���-�MO�֜ӫ�R����^%ךJ�.��-��O�oQ�u��FG�W�v+5��E�v@,}��F�Xf��5uR閳�8?}*U�ӑ��"V�.��-�A�����k�H�J��-��B%�4@w蛻
����T?}��t�9uR�Re%ʵ�.R���D���S7�E}�-gn�D�RM՘`��Tǋ<h���Ub;c�Tݿ�S�R'��U��x��?��}�ktԎ��)u|�[~�$��p�*WӳW�^�1��'>���o�#�I����<�]gO�g�=�pͥ�O:Nm�`ZLmy��2�S�+m	(��Qj��Շ��w'�L�RA�F���`��{Ka����:�;TP3�Z���3��@�憨�l�rH����4� $�B1���.a�	�����|h�������]�H����ɰp�4�[()8�rYQ(5���4l�%�ff�C�k�e
���B6-�ON����S�]�`����bTP���I����x41�K��Q����(k�ȨEq�Dg,L���?�=��W����/߾�`�h�F�[	G�e��	��c��p�G�����@$�W� �^8�	5�0��UsK;�%�ւ�\+L5}�B���McF�T�.��H�wŅ���k*᪗*�0n9Ң�"�Jj!��Yyh�2wa-@l?S������Y�:������� y4��r��I<�}:�l��Rl6�vF#�I�������������5?��[+���˳bu&a O�FIb&R�J>%�Ek�!L�E��$�-��0{����Vy���3+K�kҡTo|�#_�����9�����ow��Rp���$�K�Bf��P0��*    IDATV��p�����Ɉ�W5�4����[��|>;�q�2jFd@O;�� ٯ��w�y��0bF%�'vb�9�-��i\=&0<�W�'>{��	;'n��ŉ�v�l��Կ�HϘ�{��IT�����A%�8/"I�A���C"^����M�g#�R��z�� ����'�7�[W/ۚ���l�SP�|h,�t��U�S��xk./
�Q?<���?���O��m[
�^�����~h@d���Ұ�F�a�����>�<8�rh��E��ы���W_��k�]��U��ظ�=mJF�=l�����G��z����}�2'�%#xr��2�dC��و�hi�e3�� ﮁ�5J�c
�yFs1[#oMZ�#��"֎���4ms_Y�2��.��)?���sw����*�|�UKD��x��Ç=��;0}���.��qg�=�=��cP���S$��������x�Z^�NT�뎊�������4&�������J�^"-�P��hl?c)��7:�����F�Zp��^FI�M���S*�V��wЧ���
��<GW��Q\	$	ȇa81��}y�Ř�-R!o�H��ID|4�=���2�%aI+K�r��	�<xp3#vh�&��PĪܸ\h4��5f�S	1�V.�3�.�]?�(���!�<Uv���ܼ��JC��H�"�.���vOƏΩ���DH�y�Im��]]`��YO�BL�v����ځ�}}�����˵!��u���gf+Kg,J��30�����M���,��{��;��6����ds��b����^x񙵵�zD�z��F[�%�EKD����cz���`�(�u@`�	�ӂ�����|�K(��P�Iwמ�Ǎ�J}�̅�� R�#
�#�G�N���D���&�����I�!����������"*kYq�kq�jc�%z���|'Gv�gG�ሣSZ�!����(2yY��Kt1����"�%��}�;���7�1���sǣ�wz����A��2��'�"�h�'���wFau�ួs�����޸)>���A�3���� g���ey8hOc)�&	,�5�s����4"�«	��u|B��x6-�,��l��
Hq[��ʅw,�B�6���?d/vx�)a���;���I�Ze-7w}��߽򡗯�v:����C�:�*��+�zS��
(���K߼ Fy�py�&_B�-k��ԩ��dW΅Q�/-��l�Vk%��h�^������I� �؛����U���E�Ea�X�q�d/����=<j1��s�>�
$l���~���x�q�I��A,!p�
M���\�4���b�ep�A�ā���-��T!l&�\��u���xD����.\*�W�P,�h��ِ�������0������"w�0�/�;����Vd$4A���R7���d4�ژc(@^dE�Y&7e7�&�q�ͮ���Z���_�+�=�O�\��,���~g��o�]�wq�p�?]�s^&�@����U�4V�帺8��=�������L��P���=�u�����s���԰ȴPg�A�B�������#q,��N��_�/I%R(�ݷ�!�����A�
�\<'��^ô4�f��.� }Oh&t���T���}�v��Z�s����D~��*r���i6�Aq��*����KW�^����������Aw8�Ա%����1<jp�E��j���`��W��])�_�r������6���k���_��_��:��n���T��{�x(1�Kh$F���d��M�0>$����/%D�&0��[�,,��.q|���/�j�#�60�	����4�8C�ȸ�٢���D���z�f",�ݠ��S��b���ɥ \*C>���bZG�A6�,5d(f2Q� ��:ʅ���}���].֦M66-���l��I.�� �Ujz�j�
)�Hg�f7x|r��s(g�H���¢l�}bt���[���G���\zߧ�����E�C��\ao&h��i�bw'ro��p�^��׿k�&��-v��m�q�00
g q (���>�j%z�đ���@����i���Є$7
������,�ݓ�k[[����k�3�e���>8u{aQ'c�E��r=B��.j7��_��w���qg�ui�}հ��%X)B��c�'>S�p�*z��6�ߴEy��!O��x�w)f<-�da�oײXxfE䈅�?x�+�����-aS�n�����j�`(X�Z�0��00�(�0>J����������=)�+P�|v���9v&>�� �t��{LEls�B,K�xA+#�f�ʖp���`+4m$N1˼�.%X�ٸ���7���4n�pkmu�BX�}7�SP��`c�U˴	n��P� 9�8VF�R�b�+7�P��"C��P�0�0��u�Z_�̪��K�lS�γ>Y�V�p�f�=�DTb�K��*�i��p�艳	8f��V�ԔR|�������V���lo�h�{�1;⦏�,�FS�sb-��Mr�sU��t��������̋ oc���7��_g1�B�L���֌�����<�>�9�	�[�����wח�4J�ONX�i�]BCH�,N�'{���dT`�t�Y_�Xpw,{EfXQ�����5�u�Fr��ڢÇG�����fp��c��g��-�����Z]�6�V�5��P�|54�܇�'��&�#l"��X��Msd��a������h��>f����Rn�V]�f���տ��ꥯ�ʹ�Y�L��ΠH�(kh�x���dV1�͕̒G��w�B�4Vk��1/n^[�u�
':2!ao1i���aؑ�'O�l��<��$P�p��	s�����Q�
��J9i)E�m+ח��Jq
����h������Z�*��|���Q��;��եQ�č�eVk��F��_���l��uڲgA���3����6�]l�M^�R�a�c�#��䘓B�f�V-s�шDc�x%G�R�<����G���q�#jv�3>��O�p++�C����	jE߈��9=y�}��7���j�$VVc[��s�D��1���>��l$38�\HFcA>x>W�˅7#�&�3Ad7F�B�$�:����R�2�eӆ?���!�s'�N�}<[��Ja'<_j�]�ݗ�כ>9S���[��3�����JE�+�G�~[�[�s�X�l\��v�����@ZJD�����rr���4�n7�.�ǝ����kKk�W���ߜ��.�3��x�t�~���@}�9���n�S'Lg�>���������~k�ĉ���,�d���Ⱥ�J�|�c}F�=�~¸L��g*IX�(��0܃6A�t+�֓����3[6�k�\{��`�	�����3�-W�̊	�]L"&O�AV��b ���{5�g5Q�Օ������Ν��Iwcem̧�n����.��h�l&��g��__�7���߈ڡ��z�N��[�0��v�Z&����2�\�l�Ǉ��ǿ�G���B�5Nwn�ǌ�����`+獖-R)o�=�ů~u��ߞ1G�H%��a��z�6���hf���d�j
�ye�K��p0'�e%P)�����B��!��&Un�d����Lߏ�ó�Ȭ�0�5����~�U]���g�ۯO���ËfMD[�A�î��5r;#�P|5���E��b���0\�~Pōp����)����jC�k��S,-?|p�M�9�\��\Y�v�W^X�����旀u2>��v���
���;3�� R��n,��w=z��_����FU�� x� �=�~x"�	�~�Z:'P;��a����T�IT=�jڌg2�柷c\R��U��S&3=�P��wS}����t��ҎOi֑�~4�:�"=�:���T�Yk�n9�L���1yX�Y�M���
S�[�l�(�9TЂ:.��Ķ�]��4�=�:x��u�R����P�t��.<��sR�)�=?�J5]���t��p+��Yy�N/J�^�\ORW=�W��5�*+q���թ3�w��$|[M��*<m*]8+�O3E��L��۷i��O�1U��ѾÅ:>_ �q�a|�R	 ;}���H��w��!�R}��W^y�c$%(����"�ݸq�ZB?TպRoM>���Z��j���t�>JQm�ko�-u���?%_k��Y�I=�8K
"J�"�v<N���ʕ+ �Y��%�����L����j����`A� �Y��!$	Be>``�@�*fk�,�@Ɖ]E�&��2�=qw�����kG����NM����DHɰ�Ɛ�c��k���E|�Z?��I���x�[�!+[>	�}[�m>Y�W�Q6��l�G�03���Ȳ%��j�������!&�&V��9������L$��ވ�ǃ�ݻ�߾��Ν�w�">��5-#�à��$���R�N��%����(��a� ���܅��x����E|Evd�����tׅ#=���>-I
�՚��y�����az��.�����S}�����C�ų~��^�⟿�$l9��A�0@aKhU}�� ���n8����":{]���r�)�&���T*���x;���9Q��H%B���\�v�Y)5���2,����C���&��\vڕ���f�ƕ�3�j�UNA��/���7���'�<?'=m�:?ysx獣'G�����,v���b($�1SL;o��Ab�������$e����7o�x��������w�M�N�N�X��է=!�r���DΟ�ZȤ�Y�K�^�$$8w��7�@�l2dj�Hg2��⳴(vTu� �oN��P��?]0oX�&�:���VJ���R�����7׮�U&�X�d��L�d?y����nV�-t�Zg�:�/����g��,�o�I�C�-�U���H.���������#�,��r�?��������07kza֟����2r ���L�v��"���W<o���Z�ӝ��'�m�KuA���I�Xi������W�փ�LO�b'���X;��޼��[����#_D6����q�J���)��2ƺ�?�r�A�\G�{=3O&c'��q���hl:b8�I5�5�h6�J�+^~�^[��j�U���$���5�b^iXF������g���4����C��$l/��%�����Ǔ�l�=�l^�������%DqTl�����~�3J�R���t����#^�X����]y���0B$�;��c|�i�t�n�vE^^f�*Z.�ZK��Ņab�k�&⵱L� �@�V��l6r9�vH�F,Uҍ�},#Z-\�"vS��о����`��`xv0��e~�?�C �<K8$���RE�҇�V������݃�~;_���Q��f>���͍J��Ϸ��v�(X�\yY�l����xVE�_����	������:>� @迭}p����Zc����ԋ�~�?���gM�|�s��[A놧��R��X.u1 <"2,J����y<��P�|��I@Jb5ܼy���k����8e�<�j�g���;�<|�в��K9Us����~��X5ש��� �pH.8��{=~j�6�ǡGB����6��<*b����񜟴��,�*Ey����+��ѥ�̿��/����B��7���K�"C5nT|��7�	A:E������;Ov�A��T��]�DKaJ<Au��_��o������]�!R�{[X���ٹ�(�T�rb:���O��t��	����������bmyc��m@�mX�Ě���%��	��������y�� �1ı_��{{����F�pϮ1<�B�6�汦L����wϧ6������|R�*��ˢ�@g��7Te&Yiem��κsT������R~m%W8�k�ϕД�!Y+��%�+���7
�	eh�h�8��ȁ����Dl����R�/lUk��H����_����������d�^g���g��z���^�R
��W"
"_���7��p�ëڨ(�i9K�!����;�2�J�Fޑ
A�k��
����^�,��L/���s�1��&+�?B�B�-�RW�aL21FH�����iS(eẌP�C��Fo�v�Q�g��l�[��#{syV����s���`(
'��c�If蒳�Pؤ���ʈXG
[=o`���['i���X�.R9_ٸÏw�%X^���\^���W���4��G��άt��y�!MC�V����N��������l@?�}��O�vJ#$�F"LȤ�<�uD5B��`����x]v$B�+�Rha��$�}�B�c�9�g�,��SN����"?�`q9�W��#��y���b?����W�z������ݢ8� �a�DgG�$�)G>���{����o�6��f��I�CtNT��������a����Qy��`t<X/U�W��X�Z�����?��\�UC?�o]lO[����V�	�|4ʁ0�>����������Oo���.7��L�X��`hF�3Y��6#�@gh����*��Ot���#�]���t̀���ɐ_�.�t+,
E)�����j06v(V��H���(ڡ���
����&�����=�?��Sg0&wÐ'(�s0��ǃ���qg<�����0ï�<�>��e��zB���1��=~��������s[�$Ц���O���^����^2�h��w'gG-�0p�b/6�,Lsܶ"v|��@0��ݻwI��.�]��Z]p�t�6�V�74${:N4����~��`]?���lT4�ۃ�Q��m.��O��*�`]`��#̪��#6B������n4��Qg�����W>��^,�N���Z���/q�+/�m?lǦ5Ƕ,�P-��d�����+7�ӣ#z�K	u'��+�����F].nI�>��g~���ʧ�G J�v���4�fz8+��b�hb��`���R������������x��r���>V6����=��5`*��`F�g!'ڤڔ�F���T\@�A4�\[-����a�`2եե�um�6/���b��%#�Ͳ/�s�
F`w�����Ed-���魖�ݷ��s3�P�'�>����k��� �1bcF7A�떨ZPYYI��PA3�dپ�)� y�w�v�̴ӕB�Re��F��9����p����,���n���<3�>���	3��I��Ys��8��\�{��������.T��@�;&��z�*m=�ؘ8c �>9�1��v�����B	W�ӹ�4ZZ޺��7�f�$��$�LNFQ�08g{ۏO�{TL��XD[9+�⼘��"b��~��#5"��C�� 37��A,�5�|奅��ϫ�%yK-.v@�Eqe�>��z��7��8���߹�P�g��n�|��&�-�u�/M����.l��;��G�4��Q�S��^Y�\Y�7J���?��W�/|;������FG{�NW�vx�R�X�BMf�E�3�}}�c��޾ӹwp>��,�%����������^ZoX�.*8
9ࣥ�g�A�u��G�!/U�0.1��s���#���eTM�q+�G<���x��t,B� ��:�k���jo��D�m!�����T�6��5n������I�~�0�=�VY׀ጂ��j��t�61���.2W�1b�d1���Mn�'�'�ON�I`�HD�L�*_��Ѓ�~�K�}�0m���i�h[3zS9��p)�*N�լ�d�o�*�]�t��ͷ��zԕ5y��$�C,��0Y��Y(E~�7��9��+V(���5b�`�EV4t,��@�3��#; H����bM���(E�7��[]�-�sZ�aE����Jk�g2n��I�аH"�*�/�V�V�~�}t�w8��j�-���HVV7�_{{��1��� �G��rݼ`2 ��{�iM�+����yQ����w{g=��KawH���ه���n[�X���};��R�{z��ڇrm\;Ȝ[UďA��u�S@
M,�}�b����/_��E�#6�� ��'�	�C0C/�T$����`C&�Kh �`��&�Z_���eE�@�"��5o|��F�+�U�옉O�����!�Ѯ�*�!V컪8v/�r�ƫ���W;��ܨ5=;��aLC=�    IDAT���GG�^�M�l������eec���$��
�`;�"a�'���q��c[�3r�JyM���U����}h������Wp��a�Ƀ��Ña�G,7YH
 AM�,|<�Hf������p�PoX΃��bU��le��[¼����
����I%�A](�a�T��XU�G,�nN��,�5��-B�!чH��\b�E�E��H�&�YK�i�Xo4�OB_N�!E�j3���G=o;o����rN�K���jEzR�F�_��Y�,�$-�՗�����m�LϳSf,�Z�i��Vȿ�DiƢ(����T���b���{���~�MM@���8ĔlmC�W0�!g:=��s�r�р�`Ƚ��d45��5��Tp�w�$׎ f&xG���t'$����+;�yZ?jY��-���S:�O���
Y>�u:��^�JTւs�t��^�t7=�QA^�"�W�uRˮ�|���v�Q�oq˵���H�t�����r�i��D}���)�:�t���T��9�ѻ�U�ި%/R�P�+�hG#.|��L�J�q�:����9_?L=q�³ni�#Oo�GR��K�{�uzܵ�}�.?UKϦ���sG�?�'}���Q��*=��
�S"�:U_?�se�I�OR�^Q�q��}�.��/r�"�����5B�r�޽_��4��F�#l��xo�Cj*�&ݥUtׅu�7ޠ�Ђ�p�^�M��H0M�����?�6�"R��{��.@�����(�:�V:�F���RS����1s�K�
>�#@ :����*h�Y�Ԧ:^��.db� ���U�U��<�D"�*�SI��0��~�6̙l�1=F�����ŹL{G�ӓ�Ó�����V�?ߗ�s6�<��#QL`K�maf��vAJk����/r�-�F�+��'����;c�v$�q%��ƚj�Ԫ/��V�eٕ9�ɿXK��B���<�. �?��:����ɣǇ�����o��֛w�S�iGg"�X.a��b��Q������:�ptͩ��!���K�f���#�ΤY��Q�S�ӳj�r:k<�]*W�~j!5�^��EM9\��.���.�<���

����=�U��#�w�o��$��4m�h������jBfg��x/�S�|���@`�<Iv�*	\�s���lЁ_��gV�{� 4��E��F�s+���Y�K/����k׶޹��du��F���Rr!��yQ��F���TjI�.��bqv����V�y?��j����3_�����`au�-���n�}��S�~ʼ��r8��+A�F����r_Ӟ<|��>*�h��ib']�������z���O)C�$�D��.�a�s�r��!mbb�.�Ѻ�l.�Q��0�}N2���K�O_Ԟ�N�g0 &ݛ��[����4��͊�T���A��V��X����PN2�Y$�Sh�3%/�����Z��\� 5<�?�]��f�4[g� /�� u�9���{^���w���<��Ȳ7�X��4�/\����ݏ|�vyxBY.�~��9x�g1����G�"��X�xұ����Zo��;ĳRċ�ן��6^��=�K���+� ����D���GP�}��ۜ��i͉hb0�gc��;�I}o��$�M�"���h��5;�d
���#;3�ǡ�\��"L�郴���UBs˪>(,4h���Z!��d�#�}b�������b�>K����<W�+�r�0��P�hVךeƍ�M��śW�꫑�(d3�d�\�����|�īr\eμ��W�ÿ���/bE>8�y����XM��6��ý 3��W����������;o�n��+��"�Ja���I!����>�]	3���I�*��Q`@"3��wIMH>2�oae]���j�j�]�������l#�4A��¤5���	N¥P-�ENW�L���X�����c�ӂ�[ >7�?m+��j(6m�
����l�z�ҕ��h�"j����s�ج�@���JyeI� ��~>"֋�L&Y���2$��)�.ח���:�����~�+�?����3�r.מ���f]��	<'��M��6I�b"�0l�X�ݝ�Ƀ�V����@������K����k��`T6�~[c�-X�,�7nAC�5=�0Q(j��WI"A~��ʚ��u��T�j�p0'�g�9x�R6�DW��f]�(��.@�Pc��v�7�l�s�x� �!>ט�_~0<~R�o��J0I�CƓZ�
��2m��'���WH��rye���Xh�A�����y�\+^Z��p��W�򏗞�v.�Q;��}x���WL�Ĺ�@�а�x�m���q�� ёxs ���;�����B�hà������dx�&p��c�J��M%3�B�t:�;[��V`Z�3-�	�� �]�+5k~� ���,�2Č�ON���u�=��be� �D�
��&,?��F�/���;Χ��+������/_��__}�������R)�>p��c�n��>G�3�����ϺH��?�҇��|�#��/o��.�a0f_*����%��?j4�j��W��_��4_3S�����>�;M����f*���hx����;{G�����P^��0[�� (�	>.�یgH��s:�6���w!�
�fT�����G	�,�<Q&�>�QF>�rXUc#��4�QL��7��
�V���H"�a�0V��� Ζ�xPX���,V�7��������K��X�eiiդ&���0���L�G��K��N���-5W9��m.�iЁ����O;s�γ�o�����翉�dl��o��c�asD�0����#
@lPG�����/���[lW�c�Z�e����G��ab�1�u�9�}�e�� ژ)�_i���ߙ�>�.��iWf��q���غ���2�0�@�5��uN.)���>��d���U`5c��)���+[x4���U~��̕����j;ߚ��}a�9$
���r-�c ��	����g.���k4�DD]�ݳ��� �G'G��?2�o��R�u�ٵ��Χ�����垥�,�'G�9�S�D�Qڟ�U�'IlZA��Պ�U���G������/�88����(�^�&A���T�H�8p����Xa46�o@�lǒQi�[����k�d M�B�|%�@�H�>�-(!��h�rP�=,�	���,w�t�ƒ�>�T�ao��j6�������՗6��~��ϯ�O&�PD#�Y��TE�5}�����D���ŨO;�֨m�,�U��X��\��3�\_�W�IS��O�����?o��7���C>����;�9;9�bF),�]1�δH�/��Z����x[�?~�Jؓ�k���C���D�:�D:�T'��"��x�
~��]?�'w5���&����eo�ͦq�_[s�T���[�`�
�U&�!~��ؕ槂*-�s�.4V�u�m�­���"��W6Dا�lKwO��1�D�eq������m�v��BI�Y�M䚴�����/�ب�5J���KXߪ���_���/|nH�0=}s���>;�w"Y��G�rqC� ��۬� F��:'G�o=���G�5k��tDY�DC��܁܀D n�A:d:�JHcL���q�_��)�U+�g�C-�����*OK1��q{�h{�������}7ǧ��K��=�� �h5�\~p!�m��%g�2���$�~����^���_���⒐��2�wpp"s�"z�j("6�-(�rY??`�6��5%	�������:��J��ҥͭ�ŭ��u�����G�c.���������\�x ���Z�S���! �h�p~��dtrzv{���G�y�>�fcu���_|Q(Z���@�+�ğrB�8�w>��x�<bQF)[(��V�W)�ˍal���h��;A�
�h��X
�5q���JK��R�.T+�=��'�jȌ+l�b����2l{�KM�*��� ٭�^�6��AW!�,Z^�B��pKk�}�Qk�L,��F�wZX��Rm��v��%3����ܽ���X�F�oV矻*�O�|�������-�����X�Y��h�l(�̰����28�NQH3���9�[>��e�ջ{w�µ�5	w0v�zy�ꕛ�k���,���Od�����{{o��z|d፥y1&.�W��g,��pe�6�&�+��O�<l�_�/�񫌩�Q;H4�\ޥ�у�Y14�<t��+�\��qe��0n�ݍ-�ɳV^� �T���~^]\ǈpf��$3����C�0�x���2�$�`tog�#��V\��\a�������������|5��E�����c�G�D��"�fP�*���pV���'Eb��������<<aB�{��X�������sH˝-��(00X�wYDk��'��_@� 3&<�6Hv0ء��2v:$M�G�cܣ9Z,[�>���DƆl�L�(q�N�̹ì*W��B_�b�l՚�럼���������ޓvi���}�d|~x,>&2�>�&X�½����8�Q� �w�>�fo�bҗ�����x�t|֭��*�ZO.U�o-/]'�i��/-����I~�-���\����Ce5<g�V�p^h'�!�i:��J�gȟo����'�O��\W򈈋@R+APU�
���k��B�h�2h�:�G[�S L��f��펋PSCVb��N_��M�����Py�*5t�͐����\����X�ml+rm��s���/{�Qi�G���ȉi*U�u�b��j��f���R�z֥��?zr6�K��|eaq����ƕ�L���b�kT�D\vs:'��|q��k�����7��W�O���n�N���p
��33���� E��0K|�o~��ƣ#��$֚����i5t�@2���@K��\_�~��(F��74�z�E�]��"�Sǂ��~2��Ś��Q�Ī�v��b~��N�<d	�رί�_�zkS����Z"� �����b�J���Z
�Ҳ%�ZRqb�M30	w��2�<9�V��~��եj�w4lӫF����3��k�fiVnn��W����r˱h����m��p�$�>�	�+!�����`�솓��'���>�[�԰��27��ѝ�	�EL������P����(L�&�0U0@�Sө�ÑJ�T��õBg��R�W���U�Y�9'�����xj6�Գ~��\��)Gj$���)%�Lͦ��M-��S���uj�-���L焖��TY�%��.�^�Ivj?A�-J�3LO9+w7��g:jDe>m���]_���)u���So]��*�c7B�S3u,=謚�[T��J}K-�מ}����+�.G����(q�Ro�l�����l��9�� ��$Y^jJ;�ܷ�z�R�Wk��|�~&(i\���\hMe���.sO;#5u դOT�ʕ+>�ۃ�E�觷X�u�s�]f���c.��l�֭}�C��k׮�k�f<��s*脍Yr_�z�F�JŒ�#���^���:*���Ry:\{���q-�V�O-�~�Ns��y�&��}^�I_�fcU{Ͼiζ�s倷��)p�P�G2��MV��0x��x��$��ǂ7T>aޚ�L�Cؤt��<wK�s^睳����u�����s�	B�o��o6���V,��� N����$�����ä��������p�*�`�9�I���
r�v��"'��W��3��9���/���x���������w�>x��Q�+�^����z��ڐ�_1�@��($2�	tv�e��4L>A}%�]��v�UA;7�~��¡��T���Z������~�N�h�Y��rv���t��OGj�ٵB����EjV]8�N���h�'�@�h.��^�:�Bfh��
#&�s�C����%9"���,2y��-��N�a�}�d��'�����¬�8�f�s�?^������'ɒ�@�yVfVfUe�]}_��3��  H�\�K�rI�j/���2��Id&�7}�Lf����qIە���0gO�G�WfU�Y���g`���ud�x�"<<<<�=ܗ���K�?�lq���N���P���R~�ϧ<�L��j��
�B�^~���z�W�[XyḰ���̱?�VVaT06�8}�`���^� �,á���\��g'��Gfh6g��zx;A
�J�y>���Ǡ �ˌFG�#��S�4"��Sm7�s��Uk|h8�`�D���h����sf�2|��y�ĠP��R��x&3ïi��t��-�1�1��6b��:=1D�r���b=[|=�������+�����r��Yq�|�=)ИP�ԋ�RW<­��Qs�P^��7����p��a����˯�_]��y��k���_���}�~�-3:��Av��g�b����̭jt9���b���ʰ���k�<:y�q�`T^��$���TW.|����z���z�2 �"�ߌ+�I�oES�{����<�k��"����3��6��|؂�a2^Қ��J9i��)��U�u�L��ҹ��))D�XB��Z�ȑ�4�_�Y�1U(>����������Zn~0�i�:;R,�u8�!��-TD��E�F��Ϭ�2�!��;0��H�g�dWS<�m�-��_���g��7�І�Qo�G���#�i8�4�M��iD\0ձ��A6حF�q|�^��G��H��vF��g����hM�0��� ��>?�q�_wCmzA�����S� �˂?%�5�����<��BSi�i	Z��T�Cgn��@�)�97�"�ʽ0T���h��!*��!�� ���dv�N(���3�����Rm�W{������BѡAD,s�;���.Є����{m�V�Y-��;,�G�C�siav�N�>j5��y�7����wsg�A�t�}�����:�>��T_h�#\���U���7����?��vJ���"(�0\�q��W>��7H@/�q��V���VL�����S�(݆�
���ȎD��g�P�?1.2%�T���>uDW2Z�@��)��!�k�-D��ؚJ���y� ���L:���ύj�+\�,|ct��o��������*�~��TH/�k"�Z�̧�Yf�k+s�7ז��*�3�f�ęK����xԋ3o}�So�k�O&�/���;�n�;|�=�Nda��(T�#U17�H���fW�g��Z�w23`C�i�9�@qB�N�-�-6���HM�H�Ȧ����t57"S~샀��H姟FD�_f�������5g�e0"Gӊ|=�8��w�«C�/�2 ��K �U
�cF]�/!��BfɁ���N��K+Ùa��ˋ���dL$拵l��%�t�wnN��o\��q�е���΂	؀� 4��=���@��T����������w&�{6�z��`O�J����zɔ�X�M���:��s�4�H(�jo�胻����Co�b��+��� �FNX�y<�@s)��=� �)Gj�j��l"=���j^v�O�t%t�g!m�]�!��f�K�2���)�#�*~�ޔD�\�!����l3��o��7���~k�ӗ.ܞ�P>����=���Ys�@(9��e� �8��GO���/PggO��w�����ŕ����L��q�lv�q����i��׾�_�E��7c�g�о��z<������N�E�#�4�F#��\��8�~�����?�ރ�y���4�r�!>b�P�[��y��P���|DȂO���x�)/:(�GC����4^��نŴ�?=UR���NnCCD�T]̢���6����n%C���V�`��\�o�2"�x�ޘ��r��+uZ�C4yB��;SB��\+�gy�f�4��J�����ݝ=��x�23rve�VZ)�Wsyf(/��ݼ��\;?�4����_��o��wsٵ��<|<>x:8��c��}�>�۬0k0[����;�5��GO�7�<z��l���J�c�j��Wk-�IZpѝ82;0[ �E$��'���;�:�_[�s���؛��:��M`�1P���р"���v1���4u0�RPd�RT�Bz톘F$Nd����^?�_�_�U�U��f�H���p��#5��7���,r    IDAT*�.o�v+׭fz����/8s\,-���j3k����::����ү\���"��Η�_�lo��q�`��<�$�L��U��$��\�-�!��#,�mΙ!��� $LKtZ�LP���Z��T@]���]��G�R�=%�n�۷yQ���+�Sk;�H����Qو	K�Bw�M¢s(�ڧ)�l�H&��X&�,�}p樺���V�����˗�7hi;�E�B蓄d�"p�p/\cf0�ٹL��	u��l���Ka�R���I�<���]��o|c��E6s#8�Lk�w�����|	l���Z,^���@Y�	8��X�bw�9�e���~����Y�d��j,*��PpBCzMzdP%p��L�K�!�`k*��W��z��r�k�V�����|�O�Z��{���|pg�Y+S^.�/[ÝEaH��� �@�1T8<0��"��Az4`��!C�qw:�Gp.;��xf~T??���6��ӽ��z��=���Bp��]�l�����i6ڇ�4��κ�fg���f�:��מ��7��k+˳�I}n��B���;�/�=qh#&;�'Y����n$��a����f��
f��!��f{pp�x�����!xXGt(�e^~��+W�$Kb Oh��a"�ó +�����?����ۏ�S�a�;亥za���6.����X��0و��s�u������ӧG�a5s�:ֺY�'�&%�0�>�Z�hâc1,`����1�=m�쟶ʥ9[������W�/]ڨ>=�0�q��K��>��NK|�?�p����q��R���q�y�{��ɃM��Gǭ�6�����zn�^����ɞ[��啯��?�,sBc� �O�;O���D*���Lg�$jY�!!``L�=,�{�ۍ{wO��w��\K������%�5�-��ϔ�#�^���eb~�d�$:������{hK�iZ馢U゘(l�]驟 ��{�rb`p�,2T��xD������>����O7/t0�0�+{�Mx���I���a&s��~}�(�*6=Ix:�r��x#Y�p�1�X�hR[��.V�y��#�f�᣽��힫�,]��A����q��o���7�2��n����ΐ/�N�َp���.ֵ�DG�v���e}r�w�w7��Z�13�4S��h�l�e��Lly�g$��S9v1A�Q��<��8�i��L�o��Gs��/&^^�a���@�Y�o!^�t������8L���� .	=AM(}���]
��'e!c��u�Ͱ/$ `Ea�efBm�����z~c����k�:@�M��{��r�6{rxr����[)�Wk��
E$}����¹����������t9s��|�|����.r*��*1���nMZ"[5�Ik��������Ğq.�HQ�\1a5yoKf�ӍEo	�ꁛ�r�`�,wQE����q�28��i,���4t���Z�*�A[!�����^r�<�T�i)V0��(�w za>D#Ʈ3})�&�o-�r��Js��7�/Ԭ�N�=�X).��p!����d�(㥱7SU
��~�ڧ���q��s'���zq�������p�s������L::z����6b�ѹ=4��<<�0�bȣ������{�wx:��H���t4��� �h��I���&&L?<a�DJp���TBf����?��/���)#.B�}I��$�+�H@p?�u^�NI,.���+��k6��Ծ�-����?�\�E��jضU?�ìa����tL[�3��ր�2��V���1�*Y~X9��-��{۹��|q9_Z��JK뫅o��+o�I6�k����ͣ=n0O�Cr4*� }��A;��&��Q��h����]�˼�%*R��)��u����Ǡ���0>veF�)��)H�<�'�R��OO%R�yUJz�6ܦ�~��I����/� *��ҧ���Q��<}�n��ݕ�>oIjvj��1�Ґ3]�1u�
Ei��+�u��d���aI�������>G6�e�ƪ�며��x�re�6�(}+%R9�U�12S��K5��ӇR�)�d��LW��Z�wSB��-��{7�E��I{*Saҕ�+�
x�6w�2=r�oy$-_HX�~u*� Ȥ�)S��ӏe��8{7�U�G�5ݻw����`��)}��$��ipU��TIzˎ��h���,^'���j�w�t��,P���F��H�8x�
���m�d�_W4�c��VuIӸbzp<�{��'��o������2�w��/�@-J�a��v�h�^�O&�S9�Vo���^�Ȣ�Q|Y�����ju85ɋ�QF�����]͖�yr��~~}���kM�����2�T��n�����BS4��Æaˠ6"D �^��%ޥs�s������L����I�4���q;��c�D�à����~��A#�á
#��ٷGD�!jK�a��_d����_��R�b,m����ւQ���\��!5jvF���'�v?����̏�=������!���&�E�ј*g��	 Ճ�%ܒ��H�e\���])S�T�݈�$����N����.�>��+i�S���9�ˤ��Xj��%\��JN�������i� �hdJ+���-�0�yD�(�E%S=��"o)&�LXc�f��b���P�OC�w�V��>�[[y��P���2(+�^�{,�s�3??s�U?�O.���^���/n\_���Bgca�����VF����W^��ڗ^��7�|�W�`��_g��T�6�?:x�akw�����~[!�u��i�$<�r��5�)8��9]���v;w��6hAX.3_������kk�p� ,�d�a y���Çէ�]��|*����9&;K��%��r���#���u���	s9��tbu�ǋ��
�K�������1�) ��,�Ɣl(]x�F��d�c{��r�����G��h˙�|!�B�6/0ǘ���,�3k+vSݹ��Ջ���'�#1�fW�_��[_��?X��m�m��ս�ͻ?>|�zb�����kx����Rlt�X��lN;���;?�Vה��篝�s/�q�|=W�-�>���?���7'����|���q��2 ������+A^���c��e�<�P2MX�~z(hV�ݞeh8�}�WC��ZF�x��7B�Ӎ:���Sֆ��lթ͕��/eֿ[���<o9�3�5f&m�2��+-I�������V�v��r�3�������I{��q���_��G��/�O2�zl�b����y������d��>�ւj�j�l%�ȶ��g������q{��-g�h�_������=�y���Ip>6�6Ӟ$�!��X#���R\�7�b��@��/�ؗ%w)N'����-0 @�y"+J�v��s<8�fz�q�a7����J3No�$��W�̼�'��CY�;e�Q��[]>�خ��OGy1;�����7����^�^���zs��Jy~v�D{̕d�� ڀaa�P!o zc�8]ن�Lic��^�����յ��?�W߹��>3�:�]j�ɻ���1W����tf�&D�zf�J��`"�Jy���n���I�`�_\�<-�i;w���|��%VW�^���t��~��O���i<x�좦��5�ӄ�	�E��w!�QPRN*�^��ٰe�:S���0�]�3\��k
�u�^` �Fd�Ga�B���g�9(זH0�֩q����|�0������A�oGO�3�owLB������<�\�粢&͞�Ϯ����n��;�qe�����~��o��`��z������OLFbKGd�>;:ˁ��ب@v�O#�n������b+�"�%���9�9���Zݲ��Lx$E0��4߁.Dj�kJd��H@�AUB���)m'�	�F�!���<g�s��j��&���
3���B7�b���*��8T�0�%{K���I틕V�ԭ���n���Df����'���Q{�oU˹��l���`wo���Ǚ�S�旣n�Z��˥U�?�jk���ߺ��$;�R�{���������A�j
s�i`�I��a��D�,g)�5�ݚ����ݻ�j�� ��� ��D�^~Z1-�@d���!���FZCA�[�^�� dPn-a���35�����ӄ��C�I����)�ˋ���LEP%�a7d��;a\(���Zj�:�_a����D�!s$�srh��l��|y>�.�����g��Z��
uO;-��<�������&�¦��ꔂ����������.�=p�Z�����ۿ���g�6n}x��əS�BPH�k!��u��5v�#.������w��2|4�����vό�948�p�C����j=
��ňƚ`��χ�p�y�G��x��T�܎��Ka��|iG��V��t���E�9��S���ٱ�Jt1�S�#����K�d��������������{���8l�vZƔ'��"�Z�u��O�if�Fc*�錐��3.*�
��������닷Y��g����}�w_z��iv��&Y���zO�Ϻ��n��P��T��)�q�i��R����{��s����8�1��4��s��X+J��vd����F��W�)<�倞D�?�O,7]`.Gc$<�T؋F��X�����\�mp���
������6>]B i6��A*�LqB��_�t~P�U�r�K�_^�n�Y�~~��|{�u��r%;S/2���2�D߬~�ǣF����>m%B�5����֍�o̾�{\�g/�"w:<y�}vo���2(�BT7���ج�D�:�l
t�6�-e��> TK�!��' ���V1;Y����1N����Ka�T�G�,�	�*L5�2����Q�%:6&}'Q�ĳ�hƬ��Z1�&c�|���Pr�N�Y�E>78cq�6�n6�LƝ��Lu�*x���2�ȗH����Y�̭~9r�x�s����g�򭗯��?ͯ�VnB���Nwog4>�az���h�iJE3u��h�!	D�{��䃝�{o{��Si44�F��0�8_cb�I�p�����$}H�t�8O����8�)-/��/�i�V0��0H��Μ���l���T��D�[�3?q��F(��"���U�`A|C=��09�eW��.D�$E(2W87)}~�r����k�f��Ɯ�br65�A���qK.xo�k������̙s:�ɶ����lnp~�t���E�z}��o���o�a~�w���y�d[�m���؆�g����ЂX<ؕ���
S�QyT�����c�x�I[f� P5�7n�x��W��'����Ŵ���n1mN�w?��������#T�I�_,U�-��ϯ.,W���������sQl�;�yt����i���L�\Յ��<"��mp���P X��; @� ����O�cZ*��>�M�\�U�Vέv�*y]��Բ�.�Kfѧ.=��D#r�ܵs
~&�����I_�c�3�^�G���P[(!ޭk���֫~��ǳ߄_�Jwv��Z����&�6��e�n����rxN��������?y�nP���j���g�.]<f:�nqB%b���Ex����ӱc��w��F�y�7e�AL�%�t%�m.�
�M�@>�k��ʘ�֚)iRB'�i��"�����Ɨ�we�\nr�l���Q�q�5n�����m��@|Q���,G�E�|&N�`�>�HKD'�#���}P�Wj�V7�.pj�����l�Q����\���?+�R�!7;�ڇ��w�O�:Ⲱy�-�/t0�h]s��w���wDfg��I���[<�nsS�5�aZhG�H�:���]M�K�tX�\���N|�)�&�F��#N��� m�0�L
�bsˬ�,�./_(ghn$:�ѠB�|���R%W��c �CR�gk���\���7���\��R⇜�t{�(_�-/��0�Pf�6rX^��+�e>O|:�]���
3㋋�s�3+��J�"|��/ܾ��7?���ތy)']�S���o��U���͈n�L�K0B�Z|��F���o��}1��E�+Tj�S3=�@�]L�T�� ��d�z�O�)n���%�U�2�lO\l�ز����#��E�#��BU
�XGH�,����.����Ć�Ղ�BgQc>h%�%�)�mv���2�~��Oe���Sv���PZ�JS&	\JD%2���qXe��<�u5�����-������֣g'{�g{��i�߁z.l��W�׫�����K���ɹ_z�6h=9z��1f.�9ʐ����a�Q	ot��ƴŷ����~�уM0gt>�t��y��S��[`����O� �=�M���L���.(�Lá�Ĵl,��,��]'uǢ�ת�Q,����1<�>_��V��ݦӫ^��E
Wr���K��?qj3؊� ���LḲ�@x#�h',�Oj�2^�/Γ�Z@�$gg#ⴀ`�x���~��ÈM~��P����063S.8�<{���7����/��\�<�dMx�s���A�ṳ
�aS�k�m>j''dƴ��A���Ï�of�Z}�'��z	�	Pχ  1��yX��+�%���L�W�8�¾%ᑄ�T'�%���(��J%���Q?�ݥ%T���ue�ϔ~�'*L��<阇�����ds��&�UaW�Pj��r�Imp���O+�
�ޥ:夏*)�uż���H3�S�<��)_m~�!}:������������Hզ��G���6/��T��W\*q�G�ڙ�^L%SO�LMRXU	2N?��OT3���3}���R�S7SSH�K��H����f()��s)�>�g~��	� ��|�P�$$}bڢ�[uz�l��� �xyD�(�|�R8R=���m��2V;:�z�xKy��u��O�<zѥ�Լ��ok�7�����M��i��0�˾�x����Ҕ;w�h�ަ��Ɨ�Hߩ^TFUޢq�<UC�YC}.�H���RQF�q�`t��&~���0��|��J@D��;�֭[����#���&�Q2[*��x/g����y���&�m�BD��kgi�g�a~�����<F��l�%̎z�*�}mavq������
X��hj'oV������ϊӺ!z�?1b�;<����<,A��G���"�G B�y"�t����!%f�ؑ0h�y�g ��r�F[f�o &힀�.�R�X���q���й��X�~z"��%!G1WBO���_���qy}ڿ�*��jS�������{j���i��
���t���
�GS%<U�{zK���*(jO�'�P�W�GS�]6�2�I7���L�����ep��uBff(���5��Fs���Ƅ���U���wh�N�7>��Zk��ժ0��<�#7&�뙫_�^,��wi�6�1����J}"�Ki~�=��R��Q��H�a<>}����Y����;!����J�ƾCaf�S���q����.;�mg��{�ǧ��ynd����x�"*#���$A["�H�q���i� �.��"�5Щ�(H}P��!��g��M{p�VZ�ν�zs�{���q���u�����{�˯_]�̓nfXʚ�<�	�S��l7�ݣ�h<:i�66���:�.\�[�KoU.���_<���a�����ֽ��F~��cOY53�1[*�*hX�&�2KK��/�~��ҭ��_�
D��.c��^c�N����վ�(��={g�ۯGp]ĥ@�q�kw[ݟ|t�`T�//�Tk@1j�����W_]���ե��,�NO��&�jp,�d��͝���C�L�g<�#�F�Ѐ��� �୯���ل1R�X���H���۠Ô���A[Hu�.��� g�>7����q���vᬿ����Ly��a�������s���g�=��l��[�?rP��+�h@ ]�Ɠ^#g��aO>�^�6�'��7.���ko|�[��_�������;�g����K�K��\�&2�1>��qvS�=]�VR��~���x����K�a"C����
�H�2'?���#�_�E�Aڴ���m�'�D��&B��~vEan�쎹̝w�u�bδ����-�fJ���7>^y&ҥ�kC����;}^u��Vg�3}3';��l�v�.    IDAT�r�iQ���hf��J���DײW��nƙ���w3įo}������o�y��w�sW�Ϭ���LM�>�0:�Da��ag\���z��ڗ�k�W��-\�	0*�㝭��ݳ�Q�Yc��БB�a�l- �m/�v��6�Bk�����lu&3d�R�������s7oި��G�?���n8��u�+i�KZ~��j�g�|̔D����ˑ %�\{��i�����>��6�&������>�_\���?!�r&�3�Y-q�$�E
�~f\��m��ՕK�ϟ+.�t�oX-��o�q�����Gû���y����������g�8en�l�:�!p,ί�_���§�ʜ��qs�2@ԟNg�.a��i�U���uF����N�m_\1n!{zR�Vo�Y����?:��V�fg��S�YH�h<'�S�����iԈ-@�4������J������08�GF�ǐy�Ow�A�,�`P��p]��E�d���o,-�8��
g�^���6A#��p��4�x�3<Tkc��0��KTW�������nܮ������R�������fw83�ݲ-� H���9��wO֪���A�᥃A4A�@�奅7��r�_-d�H\�ը�������9���Y�V�x��' ��fA8��ݭ͝��}����'�K����:+]���+�`&H���	��p��)+�S 5$[y$��K(�DT��2d���.�&Y����\s�duqu}�o�z�l�eB����G5��/Uv2����~�����l�V��Y|�P��׎.l�o��/Oe����f�/�ل%���+�<���gG��e���̸�����s�z��;_�_]-u����]}�;�(,�*�U%H���w�o�����9
������S��N��J먹w������3sK�zV4T!4�(i�l Ex8�c�1C���5�m?`{�a���9e�K���à�UX������Q	g������j���Jgݡ�!,5����r2�AG4�����z�fǼt�:�)A��o��o��臟��w�w�v�>�;�k["�1��8yzg��lD2\�D�<)�f�B��y�S�/]]����U��x3���Σ��3�a�p[�F,���0C�p0c�e7CDj�M��������>~թ�ҜM7V��z��������.R��1��ʥ��)s�.�s|��w튁ڻ	��.�9��s�3��xϥo[���##r��jH���\�图���s�5�1����g'��ų����g�(��>������6w�������}�'�{�Qm,d�D�CF$6�=��
,��jw&L�n�Z�xa��~}R�e����D���}�?�t��;qKT<���jy7�e?�bo��F0�6��5%�@�(@�`A�2
������(�tzQ�t��S��a��0�I-1d,1x���j2i<z�mT��yvu�X&b���@���+XhD��@�_�>]�qP��|����V������������׽�~���ڹ����lW��v�t2��\W���]�	# geN���/��~ji����|�6��+D϶N�>꓉��3d(�L�u��q_����>`;�M��v�������Vg�.�*��^;lj��G -��[CH�	x�P�#PR���O��U������!�)L��p���n,��i<C'��ե����57�������4�[� �}��g��a�ڲg!ߍCШ�tu���A��G����RU�_�f�e^�]̽_�hk|��=�+�uJ�b'3���Y@il"Jb	���w0�X^qܔ'm��O�:[;����.~��I�W2����y�I��ӏ''{�3N��3VK6���V_m\�3ŗ:J�򛡷�ok{/�J�@�1�M/���@��&YL07��v�?�s���b���s����vO���l��/�/���v�Ma���Q�膅�	�'����G�?~*2��,d*��XLf%D�A�P�Wq������\[7E�F3�������;_z��y�����z����(�][�P�������$�g*������EvW�@/F�N�R�,i ���R덯�^���Y�}�� 7�r���֓A��?�*�t80�rq�`�}��)�lj��ѽ��^�9}���1�A���ڒ��<���i��4~wR#$����9Fq���@ ���KiwMBL�&i�Ű��E^lFy�p��p��Ήdޢ"0��:��a�=�o�P�<�Xn<ղ9vj[q\�u
������^z�˷�C���>�^����fs��!��l�oj���8��n 2OnxJ+�U={�뎙ܼpӣ���]\?�"L�ť��ο���9���L�2�q<9����]a��8l@�m՘�qW  zڷ@-���	W;���Z^����2�1ӗ�2A'n�Q��1 RI�jz� L!A��������U�I�>����ix4�)_���Nږ�*����W�7H�1[˄Oϰp���aғ�o�E�v�Nu΋S�˽9zm����d����\s~sg��C1lcD�I�?���{<���,V�e��N#��5+�Ӥ�ta�эϬ}���_��ɘ񟎒Eo>9zxo�ᮜ�>n��#��A�]�s��C�vc����z���0r�N��9�8i@@ͪ�O��Eh��cSe�,0��Li9iD|T���)�K�e#�Ȇ�)J�>gd�L�׽탅E�YK�fA�(�z�^�*���D�>�Ϗ�ݣ�c1��/*ŵL��}嗾���w��/�����6ۙ���XȂfeҲ^:;nӹE�ȔmL�n�����]�k������Z�Ruei�iE��������5)|���G��l���-Hauqv ��5S0K ��E��u�xt���ޓ�O�x��O[N\w�$Bc���O����&�N�Ş�m�9�'lO�V@~Z=S���JMN��	I�cu��`�����G�F0�-�z6z!�Z덻���3f�Fܖ&��/}�_t���o>��r-2��3�I�Y����֫?O,<�U�C��������Q�k�r渄��f��BHم�Xo��s�B�Q�v��������D��l����ݏ�?�$]�RZV�:e3I}1I��#ǟ�웟!����"v$��k��D �@ U�@O%K+���L?�{K:���?�v*�rR�T��^�N/Ԝ��*��G���ȏ�^��lK�y7=�Q����69ʻ�(�p�)�.<�����O�T8�h9#;�@���JRIm��ʫA����� `�T�b
���^wO�����Fʔ�T�kV^ZIOA�#i��I�O�/*槖�SJ�q�-��=�2�I�3��:}=e*�J}O����(�|Z��ScR;��)q=ئ:��[j�YW�b�w
8�c��I��f�?�A�>�Y�գN�}_MW��.��T�v&.�n�G��%�+ޒ�������`T��
x���NQj<U�իW��T��iUj����x�wp>�Kr�]�������M�tLO47K�4��*� �K+��b��n��j�&,��Ǐ}RO�	��
p`����ZIUi�?��O�qz�'�$�#!��&�V ��x5j�W� �S5O��M���.�Spj�l݋xļH�"�lG����3���,#*�cr���й�}y����;p��$.DZc�Vv� �q�ch9
�;%�2�Px{�6�</,��	��c�g�lF;�/6�����~*J��	<�N;�.�v}\�Vk	h����.( M"z>E����F$�Sy� m
�_IO])���VL%�$�ʻ�Q���"*���T����u	�H�Gj�3}"_���Sm���S`�	OS�]��;�W[��=5�+pۥ�3ʰ�<�!�:�L���)jv�G@�=�x��װ����X��F��q�$�K���sWj� 'ߩ�*�B�k��fF�����R+�.-Б�H8�L~>��r뙹l~N'\I�`{��qB3Ė�vs{��#�v� �t�X�g�h�����lf�,��C6�=1��=�<8hg�����A�!��۷oܸ&�	h b�S:�i#XE �GiXu9���DR� #�ӓF}��.
+xxRP�Ɏ���I��d�Ve���z��E�ZS�٭����=�H��r��A�4�Ë��o�*�Y��y����֓�^�3S]_�2�\rN��\��OHvacRoU^|���v�����l�������U��:m9�ӈn�^��p�����dS8%  [����w����q��Ų'j�3D>3�g�hr�Q3z��F�ʇO�3�y�\����h�
�s_}q���jy<Kg��b��1�A�##r���ÖPa�H� �����h�A�+��	� ��ё�@BcOe�A�g���2�:B��5^�u����:�go���NC�0�ȝv����e���+������3�k��/dW��s�{�r�������;=:l�p8�c�-
�P�y�\}��/�^�]��b������SA\������A��x�x09���	�!|e�l�d��_	�x���6v��}�@X�Ne�~lB�oS�����L�#1&~?��Z�T "�{���j5g�Ar?��H'$gw����<�MW����AF<XPψ�f��ŬV�]�[�^lz�\g��-���9��:\��Źjo�����l/�go���M�P��t�G^sv4�s!?;�~n��X��Mu3賙�/���ٍ�t������|�y�{��������CK�0�ߞj3�Oը�,�]�<{��o&�U{l�Ѭ��?>�~�9��w��}��|�B���`��suӉ�V��������~��¡��[�RƂX�D�s��	� �������7HV�2�#�s.�O����Ĥ&�F	�[��П)�X1mqěտ��������\cca}I�<���F�j@��M)wgM�h�Oz����,/Tn�|C�=;_&%3��&�_*~��s/�m~pk�~sg�ౣ³���+sK�k+W
�7����-�箇(�@�=�B3���G��mX*������y��A����x�Sp�d�Ӟ��[��Ǎ������hyqm�Lx,���
�A E�x������-��¼�@SB�hڢ���L�A�l%�A��Kk�X�9�����1V,+;1N"�3����MGck�*���� g=Ti��3����s�Ȇ�I���0W����?�ϕ�ե5Z�rnR6���kkv�+�j?�<}����・��I�r֫@�us27
G���������7�.��s٥/�?X6�K�;����K 3�&�f`1�aB�e����j�,!g�fs{��40�8��>�,HCB}A3�呟.�����O��U9)�� �is��%O*TT�fif�Z\��?]	�k�/�IY�����/��j�j����r,�S�'��iSؑOf&8��x<b'���8{!����ߨ-l���;�O���"��IchtyΝ2 	f���R�lvv�Q�B���j9������+/}���_�f��n�n2<��=x:t�'z�̰m����*�ɔhCB�ַ̠��x�GO�����׬ټ�[mE]���s�un����o0��L3�X`^���`΀/�R������i��J�aQ�`Ar5��'�w�ni;����ۏ~�|�����"�����JR�ZY����#��ٹ�>v~:��bn5S��17��n]����G��ҏ��{|�������L���|u�妎BW��
�b?K�/�g&w����D*�{嗲�/�����6w09|�=��nzB�Iul"�,9V98foN��Yf<��޺�W�����滛�g�/Ε��cX8�L� Վq��nK�g+vd���M�sS8K�G����c���M/9�� 쮘'^w9{G���4tI��2ۿ�¶e��̜�&f�}L���M�东8Ӥ��*c��Y�Y�Wh=�/��8��S��8ɿ��Է�^��s?ys�����~�m>>||<�2�L�{�	JaQ�v����/gV�:�l��r�g����n��j��0�3�����$��f���wc��L���M�l� ����L8� �%`z�P4S� $�L1�*��R�V2�8e�R��i�f�Ȼ�n��&fQ��r�[KY5O��>�k_..���?8Z�ح֣ ������=��N;��7Ѕ��� �X��+gk�3_~�⭟,��w�;��d��X>��t�U
N^T�Ոf/��,�sX1^�un������g�_�>�^��5v��w���#�S(����A9��c�mȌ��d%����w��):c��Y�c�E-�C�� 8��.�Jit^'<�5�$�y���%���~������A),�ȇ+��k׎����=
Hn����F�0y���5��
�&�>X�@���`���'�ZA��ܹ(we��Uaj���^����=ݘ�+<�������|�r�\v�g��A�ܢg �5iH+j�}�/�糷?���翜��vL��]a���h�9>������%�h�⃲:����X��i����Njnmm��QGH��,� �'A5���~0!�G�O?��?��OY����Q^8R���Qg��w~v���'1��Ǵ�>�����@q~��/�r�9a���h�aiy���LaU�6L��I��K�L#H�V`$e~�=ݻ���[���,d6�}vx�pa����w�>-n>�Vx�l-*ggZ}1��1\�P�q_'�(�����o�Z�x���/~3���LvՄj1�G={2������؎��u�-H� 
�vcՆ�*cw{����G��
���*7�aw��~�k�KQe��(j0��VP�VU2���G�)Y"��4~*��̋)�H�G�J�OE�&d��ܪV��D�)�5]�d��q�1L=��I��<!)>M��N)0J܇���ɕq����g��_���?���w����e*㺕�}h����ᐛ�0j�K�
�3\�ЗS����<z�3s���gf_��l�m���q<ޙ7�15���6G+Sv$H"1X_W����g�p�}��?y����>���Ҭ�{š%)�,
C���Uۖ �*�����;S9D�1�d� 3�?��#��
�b9 fl���E���3Ꭓ�مZ㤽c��[[��r�C�1C+ڡ�'�\���_d�	����Y�˂9,o5[~{r��+7�z�~���凓�m��J��mGԛI��iK#B����b�>9h�B�g7,͇�����̱���_����f'��Y��(C<���}*ư��L���}J��4l�:MT����@���P@����YY��(X� a�`9bd�8=��t؈c����$�}(Fs�S�e܃��
�_K�5�?���4���w�p���A5�Ƥs��z��lp�ƄZ�2"'x�ʕm�@mVװ����&�`����پ��J痐)Qo��T>Ӹ���l�ü@DLO8�=
)����
��[�����ȹk8���쥹���L��3[.��j��Q@�����˥���s��1_�=�:;l>���;0W��"�V��=w�n��@�0�A�}��s��i�C8[�;����+pa<Po�5��	�	��L���� ��VK�����i1�7kK;��]���x}�=>j�l���c�X�V�1���W���N9kN3;�|��~i�\e���vv�����������g�vq�Zi\����������7��|���w�<y����9��QI�� 7[�Y��K[���6���^������_\���Ff�w �Z��<:}�0?>�q�e?-����5�fqu}���X�'[���ȇ͖hOF�k���M��	>PTP~z��''�� �Qo����L����9mI ww������i��?er���ԅ�J=���T�m~z+K?���:��m�H%>!��kjPa���uG���~��/ķ�Ju�bI�Ea�fC�Dxţ�Si��)�-�Sx�񻚧���<��/�>-�Ҿ���L�L��R���6xK������*I�Hu�z���T[j����w_IR>�V�_�2��C{��T����]i*,GweT('��p��#�py�+M�D    IDAT黩�$��);gN�����L��JԜ��[�4q&�O�R3��ٖi��I�w=�i��B	�oi'���ΤL'ДI�
��˗/s+����}ϰ�x�<�Pch�+�@]IU���CM�����+@�e.�^�vMa���H,�/����O\�����h��u;�Q(hkБl����
P��+-%���ݥy���Z�u�2���&`!�޳1���#ʂ�]�����8�11��Lln8A���=G��z1,$V���\���x�i�N��JM���'��;씙Xq�S�נ_�����OO�J^��v9�Dk�������Ԛz��r�΅Y_6H�W��T�I?��P�<PXSN�uQ�'$/��KTz�O5KK�lɔV2�k���
�h^�� ���Jc��Li�*��	?S�=r��LWz�S���T�����
(��_��t�ȋ��^��CH�c�	i��$��d���fv�j�������9�o�>�lmۛ��\~5_�S�`?��a����!�C�u��A�*Grg�0��f�$wXjl҅Fx�p�[���q�I��D��q ����Gb�vv���ٌ#<�p�����Ł��؉Dq��8�5F�9}�����'��'��~k��>�m�K�0�����t�U���с�zђO��A� ��5�
��
 �z$\^1(��a��uH�0��MAj�L%�Uͮ��x�q6�I���A�b}�+��(\>n�>�칵�ʀ�'�Y(�Z�����Cm�g�S��M�t~��>��XY\���,�5�	p-3Y�g~nbߺ�Y�E��o���~>�C����8 �V41f�
Q�?{4l�R�1��^8�n�"2E��'O�����>��ϣ_mq�i�j2�Aq�~�ڋ�^��xm��G��l6[[���Ůj޸�����>898�$�=JS#v2���A[SS���+�Je<M��$��yb_�G�����E�[�j�+��Q�$��9�(�$�<>5�"힜˴O��]�D�� Ч'���Z{�9����I���wV�W*D
�H���x)�[M���K\�	Б�������=2���8�B�ɐ͐�Ww�$��R'���6w ���?��k�/��*�F�L̴=��ΖlRE-B��qbSǁ���H����i�Jkغ��\M�z�����b�w6'֏�q��i�]34n&�&s�]�h>�>:�-��snz�>mn~p��̍VW���mtN"��1��=%�a��J���#�U~���T]]�u�>_�,����+���e.�'w�?�Ymm��Q����<��q���,f3qB=6+���z٣���nc�y����Q�!\���:R�U\�����^����A��''N$�hi~�nY�T����r����W�\b��&��`w�vw�Ö~h�{�w���O����Gjx��)`�G�۔����6X�4U�C�NfZ��f:��z���x�.�5��  �"K=P��7
��I��`�Sgv�mn�E,�3vPs/g�.^WC�*�5R��R��~���������k���ZhA�vs�ʫ����ѭ��f�T);��M��G�vr|��[w�<������e�DC�?=>5}�Z}B&��Ya�;ƑT�0 ��0���Ŵi�,�	��	\.�N�G�夁S#'3(gI�#��Bt��;i<��k������CR��N��Z�2�7��U���͖��Y�ա��4��X�t�<��E#	znfj7�/��RqÉ���̙�N�}w�{]3�j����n\;�+]':��P55̤a{�	YǖO�����cmD�c�#Hً�AH��! &{wwNaS�A��&N4Ї�z:�m��F}T�|Ţ�Sc�O�D�w��^���cV���N���1�f����U!h�3�B�}
�t����~��͕.͟�Q,3̘�I{��l��tK+� �o�3�qkw8�۾ӛ)�/lp1K����ꗳ+�����ˇ��ܿs��-J���@�%Q,;��>L/I�a<��R�0[��p��ʧn��x=7���~@]�,w{G���#�6�Ar9��S�hf��+hn�
�T(�Z�gw��ֽ��c&#=f�@J2QAԂ��Q�%�2�G0'�=l����P�Ѐ?h{aQFa�D�R$<u7:i��?Gri�*!�#Ϸ�Ò~������%�m2?�|`�ԳA�b<օbZ[,��റ�z�m����jey�.�]�d/�?����~g>��q��\�qf��ou��uOCL���)�
�s�V?�����|�U-bJ��.	|�[������'�6��B�����ǅ�<�H�Wx>��`Y����ݸ���O���j���h�a���T���$v��,��$!'`��,�`LȬ1.s�=�Y1i`S&�s�����Yڦz����񺋄���SB��O||��8.d?5[���F,p�r����k�X$4.<�ũ�|�k0@R���R��9k�ۓ��Gkϖ_o0/��n�p���d�HXi);s1��8]�pS
�9uO�r�ԣe�����+&�_�VG>��E(g)�)\��A?u�n%I[T����)* �` h$ j���]��&'�����Lw�:A/�e�gʔP�ݕj�݀󔩌�xX!�ִ����Qso�������#߇g�n+�c��Q��?4�d��D���ިY*V�������Ra�1.^�^�����1�^͵����ޏǻ����a�X�Cd���ʍQ�r&=7��(�f!��κ���~��������dy�r
`!��q���}",�v����Q<���~�t�1t8�P��t�\3�l��)`�&���� �"v� @vI}[�4��#29��t��N*�§i��6W�X��I1��J���qu�Xt��n�f֗�s�e���q��j��>#r�j�����z׷�
�E*%��␙��X�_��f���2�˓��Ʌ�k�y9s��h�o`;��*���|��0�z��e�-�tm>��8W�)/_�(]�tf�K��%f�Y���t�ltZ'+���ی3�1�"(2����Dr�UQ�-&Eo����b&��`н��RX&�Dd�$(%�Z8>��zv��Ǭ���YL���HŚev��{�'w�>�֪k�O�LN��������W&����b��y��6Kc���=�_��b��;#t����|g��v��e�h��Q{���ѓ�f�U]$�[�z��ys����z������>����|�p��3:<8⧩-(d6g�e���4�������ҫ��>�b��dK_���z�Wl�wOv�ZO�g��C��H�A�Ɯ<�X���ɩ���eF���o�n=n>$ �Ֆk�ŕ��@�a����r���+����>��8��DEa�)ډ�v�!>4�j	�O#2�>	b���#�����+rP�)inБp�k��z��(c�x�PX�7�3q�����D�A>�	D�������,�?c���,�߰���Ծ^��+���+��W������̷���+G��3�6Qe) �`���#=�I�#}�W���F�����k����1���[��L������o����Ŕ�=JL���������q�Y����3�N@�q8X/�c����nn��`�ؼQ��yV���B�(t|� <��S�T9�k�O�E�r�{rGT@�|�3<n���8R���c`�+� r���8"�u���k�z�V���=�����	{S��/�~������l<�����O;xB�T��}�����L��8�co�<�!��/W��3s+3�o����7�^z�8�=���r����{g�*�e�d��p�l6�c�h�?b:S���ݓ���?||g�8�5��C��;z�}#��5��O�[�p>�{���l��:�J�u7@��	{!;�˅�GE���6;G�^��L8��4ϖ0Ybb���^�S��N��#��l2E|���>�~����N��؀��jm�\ά|��?������}��~������r:�
W(V��]��˕�l5 3.�,�}g�f.T�qL�&�+�jĨά��u���o�s\�co�8j>}�;:��M,Ț������f����5[�̓��7۽��j=��O�� ᧗�MZ�HZs�sc?!�
x�O�ͧo��t9. wE���zC�lXf&�{���c�rv6\���a�υ�D���D�c�_��O���Uv~<d\~f�7~{����'��h�Ѫs�bK�t��)�Qv��ُ�n�qi�I�����Q�3|�f4I]!�%�3I���e���ٵ_��a��D�a^���o��>�������6���L��[R�{e@p�c���́����f�r1��p �B(>��X>(��)�ҠH��^��?�%R:��	�NO�ӥ���65K<//Cc�Muu>d�]r�+��z$Rm)_���¾�K��� �<���2����G�)��S�7��S���i��T���WRc����s��~��QI���Ty��Ԙ�V�W@�.?�%mh�L��S��R�2�DI����*L5H�����s>��ڻ�ez1U��2S�>�*?}KB���T�2t�rRZ�rr7��ן����+�9v+�sS��ì6O14��
��TE��f�i��J�BѨ��v�M~,Y
f[�*#�s���J�h���V�wM
�Fd����%�(=R�b��?��>���G�);�>*
�j�/}��z�*ϴ��:�h J,��C��+�v5PW��Ş?^�"޽s�w����R,�@% �ٮNj����[�����׮]S^��t��z]�>�%z�/�P�� '���TF��UeD尒0a{��|�˂Y������6T�,��V�!"H�XС|���N���;��� �b���vv��������x��L��ߡ	n\�4%��)�ap�K��ݩ�Fg=��eIh��S���keR��K��G*��2��i�i\�w_TR���]	5��'蹻Ra	e�����*i�ѕI�T�����2.?�H��m�G�[���������ha�AmiL=M���RR��9͈U�yͪ�	�H^�Q0�xK1��ҧ�H+���u�K�G����͵���F� �`�����L�MK6662�L�z=���	d2Y�Ј=�l� T����r_�o�����
'�Ɖ���������F��Tp%]�vYk���*<oWMGe&?.{�q4�|?vQx`�`�����9U&�i;�Һ�9e�P:Ō�H��X_y�����R!�[��G��8�XS4�L��R9���c�Cs{�8���n9�}�[�����݋c�d-NG_��,w��}���M�|N��� 4���!�h!8 �G�b�ф�oߢ2`���{�7���@���8詯�B�m[8�xF��|����A~���`|޻\-��ۥqn0s��l�� @�7Ʒx���t�o��\�:�I �Ӎ�\�.Nx���������j��;���{�Hi���xC��#�
{��m��65?�:B[d���i���w~T�rk���RâXWB���
$� (�P0n I��vΦ_?���ΠT�Uݴk��.�����n���B[�TF�*c����C�������_�=��BS�D�BJcj����m�'�D"L��'ec�R#�� Z��&��t0�Vj�����v?mm'C�^��
GU�r�Z��튊�wzѿ,�(�[�w���ܵ2����bҺP��?uh43�#C!�2��o|��4��ގN�����k�Ru8�P+乍cP�����<xC�XS�u����8���?�nn��r�ǆAwb*-�(�P�j��K�:�$��)WJ�H&���	aU	*4#V�j��H� J�A�x��ĭ�U�딫�*�I.i��{�B8�/�ww޻}��}6�����z�w
���u9W���l\�Y*lة�����H�kݘgk��j�u�q��5�͎��7�����jmW���;�L��]ר4��u7��U�,���抁6�u�.#�v.����=vq��cN��f���wBD"���3J,)���������/a�n���Ba�֦���޾�9�ӧ�$�,�$<IOJ���N��`��3C��nÑ(�,���7�HX�!���!D2c:�"6�A�3��g������x� �d�p���5��
+��� �+��]iX>h��5?�M��Uw���_����ڹ��-��jgï�/�h�'�DKd�V�y
��p�s��OV�n)|���J����!*غl��3�I�h�59��-�1���w��z�3�j�n�4�!19�3�L���(Dg8�rB��c.��:b��^�q�ފ	V��X3�)1�nF�O�k�Ҍ@�b�V�S���Ls���׎���|�m���h�W��j-[�u-��1,dW�xE�=bXY�����F��v����~"[Chw�cH!w;�4�M��8���E�H$�;����Y�:Ӟ�m��^lYL�r�,�3�Fأ��:Π1�����+���܇׻���9ã�H���0퇴��I�J���Ȁ�=�c�m�So1J�V��+E��-����:��ub~&uʁN�������J�0oő�I��Ѹ��p4��܌��2Im0�L�@ۊ�Y��6�(�����VC!I�����(����/����~~y���9������/�������Ï�wʹ�r��`��G�s��E��;_O�׳��{,�!AĬ�6�I�����3%}������_vN�/rܥ-د��E�Z�(fb�J�GB�	 �`&��ӌ���3�:r����Hy��x�4v�U�G��P��F�WÚ���p���{���<׼~���-�4V�����'��I��*��։&��_���]���7�\���lm�>�U��������v~���-����Z��@�tmn@.�~�^o���K�l d�?�N�'�iRQW�̄;8)���2�੓�#���ĵ�%O�n�st��:�Ǘ�~��hו�(@�E`h��gN0JŸG�qD|L&RW)h8;b
 W ?��j��	���H�H��p�Y�H�/{�a�`��f�>���;w�n�ﮋ�i3Xa�\�o��	'�t���]r/n�s�R��[�~���ޤ�7\M��=�>p)w�
ifHc��+��!tꯦ�Db��|؝��9E�F؇�a�ԡ��d���G��5���,�D�U�r`[��	P8g�JH7p�)˥ľ���/1�&���N%��̛x O�� P%i`���QG� ��H6���5��ѱ�whC�y^Ois�yq-�x����Q9���O���l�;R�8��W��f�Q˭�gi�o�֏mXr��ֻ���,�6�,�asT�A��,ֳ�I�z2j�ϯ����T����#[��m�mN,���p�#>c`qhfU�z2�:}�u��z�o5J���Z�X�`���2t%����6~�sb�T͠(?�i�R��FV�VL�W~A��ގ+�m��D���q	`u����?�x�]V��_^���k\�<{���*O�t_�]�6�1$�?�Ol�3/��Ք����r�-	��n������ҟ��y��b�'Z�o��8=ɝ}���G�R�>&W���z�޺���.�>,�wБ�!�,���E�b::)Nݕ�C���w�G���lv�/laεP����u���tҦ=cb-���Ǐ�<ͬ����A�L?��O�ڋ�s2���I3���v��e���4cQ8�|Nۅv���pYr�A��1��AX�h�zV7��o=�wyz�;*���qƊ�G��[�{l5Xc2_��

��#p;l���6閜Um���z~=��Qkk�e�I�Hn7����O�����^��Aw}���JV�'|�u)��J3�h.w?,l��\�z%�x�q���vt}H����ٷ�m.�V;Ū5�� �K���R�n#�j�r4���˗���Q��fsk�r��W��zx��S�_���~�!T�!��3"vv�l�?[�aiK��O�#>���$�6�iR'�n�Hc�B]\0��7����Ֆ�]���!{�rL[�bicgay�/VL�����p��:��}7X�Ε�����?���?�����Q�>�x���䳷�����i�;�G!��-    IDAT��(��vy�nak���?�������j/�ju�I�h�WX��蒓'bFC��$�&�'=��ćZ��S*��o�_�_v�4�Nk+�m�������6��ԲV�hQ"�`��[���li���E�9&-�iC�,�%?V� � ��"b ��kj��q%-���[������F�V�㋄�JP;���!��"٣9�G6�Q۰��de�7u3�F��]���۟��O?����_~������<z��`yݮ,G��l��w�Vu���V��W���>�����v]�+���n��[�oڗ��uD�0.[D��d�����^p ��2���h��������� ;�;�b-�Q$�����hIMژOAm1���r�*���2ǈf�O�=�%��\ʙ��W��8�L��2�D������ǘ��5iԥ�_�Y�9��4��]�|sG�쬬L��,%�Ugu�`�[}��M
�q8=�i�_�/���m���vq�×�Ƙ���^q���X�lǔ��斵T5�a��7�l�؍<���Ɵ��\�o̠y�_9���-�����RW�q(�
9v��QLbw�ǹ�x�.�.;���;$��$!��@V�f:��`Z�{���`[�Np�N�K&�+P'�! >�����ۼ`��R�X3�t�h��;<>,Wn��4Nq�[(���;N5�h6�����_��y���h��Σwv�	�֕���������_�����_��&����/G�ˣ7����_=�*�!�*���v���k���[w����k�a�<m�������_�n��L�bZ����_����V�E\/�〱l�&8\Fb���h��t(5;�癫?Vx6��A� N�Ʊ,���h����	�d�A�;p:�����+EJ �[夰��R^����ӧTx
(�ޔWzOj�,��T�pj��{R��Y�#F^�@ �)�O
�S�S��ŧ�;?��K���7���Jݑ,�T�S CcEɘ��O_R�T��7��^F�R{R�w��Wa�$����S]����Rz_�S�uY4Ú�X����+��B�mHuy{R��º�J�S	2&�I��K2o��ړ~J�|a1$9z*o
��H�UGGG|N**���@`� ��|)-M*M�SN�Q�Ή�B]I)��d\��*�H�-WuR�">��
͓1A�4�F����˗/U!��&��b�ÑR�k��47d:��Hu�W]��Ȝf���U�,b��W*Re2��5�Xv���)�'�
�@���I�M�$ ���R�O���G��Dz' *6�}��)�nKc����(u	�����9(��q�9��=-�c��L1�Ђ��Yj/C��S\�9��*!DW�SB��,$��v�"���mp�0�^m����E8�2��(jP"�ʴ�ڬy(�:k��g_�����x�hz��pt-���Q�� .I*6��Mcq������
�W�B�L��	�ڊ�I2oa�1RxJ���(?��y�,��OO*J�
�] �K����)�a2ʞ�*,�G�쾦B����-������>I/Yzn��29Ց1����C3����_�����{w�䖢�|c�l0�!�ȅ�ר�+Ґ:�Q,�3zx(�c�}BJD�V��;T�-�� �
{�*#8Ҳ�	c�I�
�ipdv�,��E�.O���+s�(���	0Úz���3;�~s��,
��l��t���#��1�ll�ii��mv�Ti�T-Rw�/��믿F" 6=F$P�0�O�@y傥HJ-�O46m����?�}���n��g���U�ׯ..ή� ��9t��b�ޣ�;e�Sm՛�%�]p�C#�L��'P�ews�j��s>��L����HNyIl0�j5�D��o�`�+���+�8���+@z�t���=�´��`�\!I�q��kœ�ې�7��	U�ۗW���'_�O�8�Jc�!�X�\�P��|��u�y��kr̘a+�����5�m��>������]f�t1�>��4v�L�O�π�H��� ��G	tPظx��ko_�*e3&�e�汄X��B�oU��nv���Y�ح�l�k�ً�"N��j۷mj�7Y[i����1�(?��d\ D�����ͫqoy՛x������b����g����=]��qq0��wt�����W����C�B���ipРΙ� M\�� �h����bIX �8��'D�m0(+Q��hOJ�~{�m7�����~�Z	
�����e&��L�Q�yZ������?��Gn�-߭կ��^�}��� �j��'��K��~�9o#rj}�e/d1�i�肽�xz���Y��ղ��7��B�G���K-i��M�J�
�Bij.���No>��� �ʯ{��U�vﱁ�]���rN/B�@�L�<�0
�����M��E?�f�sH>kh6TC�z���>x߃x��c 폫 �!��!�W7&$m�|10S�#2% ]��Q�R�O�oȜ%�?'f1"�Q�XM\w���V�,Ww�o�#h.ĹF`�&��B6��G�/��:�_^�׋{����jvռ<�K���d����fʵ&L&*��'�j��!���������o$���/7t��"y:��ѯ2t��o�Q\�uMi.b99����f�o�����]�
4GX\��:�F�n���BxI2��x�>7:�=��V"P*�K��������,��P��FA��F)|���P�����g* 9��Q~0]���t��؝��������>�F��@hzzE�ԕw�3���w�ﲸ���J�^ۮ6����Z��Z8�-��B洮r�E�~�5Fק����K^ˢ�`L_m���h�F5f�)�d�N:��C�W��f��������:� J�!KpS�4b��K���T���Jl�E$����8�c�h ꣎��B�!|�.Tu�A�N���WG�}ڛ��n�YKBw����BHl�H���y��Ao��q	Sz���5����f#<��������<,l�x5 d_�ɽ��3��(�	��@}�az}0�o�� ��Z�<��	y�*0}� �Nrp�Ǥl�=�?���_�N:f��F�{CT��BW��f$
���Hv6�͉FS-���'��3��k�˜p�3�&%A�i���H��+�*`��l�79��0��4� �>{�vk�V�ThL�z}�ʯ���CGR��e\�,�j�2˯;�&���`�sn=�����6����7�@�k�z~��|�!ۇ���R3�j� ��p�o�{W|�Of��)n��^\_�J�+�M����Ze�_L4�"�^�f������]���j�(�n� ��7��߭KCNA�;~᡹d���6��Hi#������:a;:��wU���Wo07}�O�D�f��d�U�y��:jZCI�0�|���;]W�[����ʒÍ8��sȭ�aQ�L4���1�}��{�cj�����-'�z��+���;�e�Ѣ!c]fB>�����l�͛�y,p�֤�f��5��= Kݝ��z;��^�i� ������1ߥ��v�>�!��O��I��A�@�np�$�	�%N�+�1H_�%�[�44���yK铺�:��@ �#N12�#������F~�\���u-�1�e؍b���v9�b[;q��QG��]Gh��]l�ҏ
a'�E�(�`c�ێF�7�]]�Gc��Ť����P���]�S�9���UF��bJ�S�S@�=&��Ɨ�Wߴ�gk.no�S)�5/�(�Ú�CLQ�'��%h�Q  F�� ����D(��ž�� �{}5-.�3��9V���2�<�a(�K����;�~�AN��˃��|9b�y~||�f���h�g�lC��p��+���m�)��@p��-Y37�M���A�p�ːZcΗo�d ���֕�X��F +�&�w���bD��@�ղO�9o_��q�$��\��\�Z0*Fߖu�h�M��}�Nz���Ͼnw��!�9�)3��F� K�#�d_3`�6��?�	,�hn��І�`�RZbV�Pb�eܙ�~ݩa�C%�1b���ӝ�Rm��'��뢕��;S]�3��h�H|��7�w��^X�)S�8c�T����
��@����&��茽�ɋ���ae�������Ze��,q�� h��k�,���#�q���dώv����8���㣣��E�`��a��/��T��l435�nY��	�$AGE��;�����7�._^��g�6��za7օ������?z��M�5&Y@�Pj0[L�Gl^���N�j��������r�7A�x�щ?����d� 	Du�k�#f�W�p����YW�B-dvø�i�ژgk%2ưx>r�XxJ�i���r���ڊٔ�͕�m�Y=-���ɭշ._.��o_�x��]��9����|���r���֏ )
A۽���[��! aW���FP1���(h"�N���wIț�����烁;y�FW�-��5 �%`���0��,�|��b�3<�R��&��tB�$c�Jv�Rlf#� �8�X��<�%P�H�Bx[
?�����Թ�u��;�u������"\�E1�)�a'g�*%*�a�R��ڮB��.���*�M�g���N�N���N���^��Yپ�����w
9V�&i(��]�{:8�v�l^�:Ƕx��ɼ����FE�L'�L�p�GTmX,G8������d�*m�Sd �8a	�[�x��D�F�̝D�C*�A8����&��^�~���Q�QA9,,��<�R6�bm �q?8�@P�]�R��gϞ����k�qL�rX��u�,�Z֊j� ����f�����yw��.��G�w�ܿ��ъ�K?Z������?�����7��_�N����b�c �EA ��MH�q�{��n����l��ia�aƇ�*�$<���7�ˣ�ܹ��r�ڔ��QsRx����ޖ«�d�f�U{�v���GoO��-�����0zAv��H�q{@KjiD"��$z�:�)>�� /��H�!�h�d A�;kȩ�� �y^�����^�l5jNts���U�:��B����
�� =ڍ|Nا��S��a�o�څ<ክ�?�~�o����_���;�����{�M��̭Ѳpo�7�����Y������4��[�v��ݿ�����=��!�����s�r:nW��l;��7c~Y���k�ڟ�N�|�z�I��?9�>�������F��Ѿό U8�ހ#>��y��* �'?���pJ���UX�4")��)��I��iȤ��[�4|�b����H.?��{˞J�im����ڃ�U�'�x�<"�U�G�;�yө�2�T������dL_ŧ���D��xk�O��$T)��)�,�1�H�gyU����Jao�'�<Z�4�"��W-)�&^E�j��Y���.��i��R{6/"�'��6՞:bU��T����S���2��X97��S$��)ej�2������%��@�ا('�!�1�����W�&Y��S*DO�A	̆��d)%P�xE=}����?�����O-$pV&I˻�K*H'H����\�����P^%+_FY|�S���L�3�ȕ�E7�:��
����;��)�N�'ţ��F��s_��զ#m�U.��}S�^�J=)�OH�J�`y��a��d��U�5	Ӭ�z����i�G���PS���]R�\�{눦궟_���Z�l��Q_.("B�<ɬ�-��l)\N��"��.w�� �`��.'XZ\�m9;ႵK��Ma��f:F���14^Veӹ�1NN������V�GlE �Md�`�W_��U A@��@�|����h��4>	��N�
H \�z�MY��mi��Zb�B�iR	"�EJ��F��
�I�e�N%����S�G���[1QS��J�S�O
�W��W����
iD*�#^F1��5�=:N�ɛ�P	ީ@�	�K���Ñ�+G:��j����I�}q���}pk���aa(��*�C挷 ø�+��[��"5~il\z���W��9��d��Ă<0N'��'y��
��� �g�L~��^fԤ���L5������b���3Z�v�R9���>j������?����P��NZ~�0�F?� 8�	��|��g�~G-H ���'P��]F?�1X� �*�Y�=%ƀg$L+�85Uh�*�i�θ���>�nu���.y�Ώ�lF��v�����^�y>|I��ږ՛�n�4il?jkGW�����S"�Xm2���W��|'Xġ��-f��񸅈��yW�E��Qi)���0�9��	Z����fr�������]]\����O����=f�u���i��[;~���w���K�A�L�4��N�����?��s��a�<T@�zM(
��i\�=@��'����N�4Y��@L�@��XN���F�����룣ho��흍p�m+ރ��8R��`��S� v-SC|u�!N����!�recZ0U��!Z����B;�*����5���.�o4���Ȕ�<F1�K��:��{ؚ�7�-��������U��rt�.��ؼը�&S~�Bo�NQ��p�/��(�/��h0"��=W*e!�[�D����O���@�����׭�j�۠$�7w�	[Z	Y���C�s�uu'��n�A�u�g�<žO���Ҕ;����r�x�Rڽ�ְ�t���%;��n��<n�	��$�´���O���g$�t�s�D[J-�m��N�d�i�圖�M�ǳQ�-���dtŁ�pv��}8���AKP-��!'��'��hȲ|}y�<��\��\$4���S����w�R%,�W	�:�1o��H��˗Yߠ�>�,"%H���~*��Dm���1٧�]�KP�[�4Hd��<�����ϣ�y���.���Iq�]�9Z�%��
��o�Z�.j����ب ��6酙�&� �1'�i2�+������.�5%��.�DS��� ���Xuc�ޓ�n�\��a�%,��x'�Qgt}�}�u���Byowo�Z;�m5��"+�EF[�VF�G)�$�����=[ř=�� ���Jd��8�7�<��4Qr��D��5�#& ]4m��
Ô��Z3�N����n��w_�ӏV�y�kUjF�!]iŌ$Vv<����Q7`��D�)m���<Uu�	�ǽ���$�q�04�Gn��b��B�_���8��ٜ���#�+N��]�]&���  G�Q"T��R�YIq\�Ph���e�4M�̩?᳟���@X�>I,��xo� |�@'���oK��i�$:(粖%X����.C�ք/>�3��%s��;C�Qda���x5��{wytr�B8��#c�l\�F�C.q
�p��УS��o�AM��^��Q�D8�k�h'-i��E) ���c���7���tx�*�U�4�@Nz&�0B��[��T����I�GO�v^N����]��j��l8�]{�-:�/'�'�r��q�<P�����jT�k5dOB�������+��F�$6@���i��E�����梾�j0��~��x4x�ɣ��7<,/k�]���d!�ggh�1)�s��Z��1-W�.�1l�)<��8��ln]�!�c�4�đ��mK��1#re��a/�α��S���͞c#�zK���'�v�m:��o2�����}��ѯ�:o7�{��t�n�E�loN f}��c���;H��8�g�̀{����`�'�|`���&�i�p^�i
H���ݍY�_�	������T���|��L|����j;�+N��^l˼-��|�R�� /������b�QBK���֌/�ql�Y�9���		��9��3^�� ��A��hcCo�ȇ�l]���gZ�X���٬�.�>����
��߄Q�oǊ��&�p�5�
��'$�'߀ �H�I,��Y8/��"S�����Z�R��R�4L�����H��r,L�����4P�j�!w"����wP��Y@1� 'tt��1ep��3�)�gkn�m�,
�ʰPF-V9;����`��>��dWS�������|=�_�?Y�P�9��[����'Tl4E@@A?��y5����o^�~��ΰ    IDAT�ˣŜېJ�u���!�P��I_Rx�y�q�@����lz �f����F߱�h��bx5�lwn��MM��p0���� ��s�t�G�8ޛ�ľo���MVWG�~Mӳx�����F�2uJ}	?��A{C���hJX�c5��jh�R���]���#��l���i�Z�;}h�=��V@+

U�Yg��lxc>��%{��r>7��`���Lv0? �!�$d�vU�z��`r~v���kJMS2�OA�
�)5?���í�����ES2��at���}{�i�b�y��q�5p2?0�!��M�7�B�����h&�y �liSQi���o�t��$M�O���Ἲ��ـÊy��x᭚-�2\�x��P8�{XM���Iw������W��+ͫݽ�;�0�<�_�Qa1fkj�!/���^�%���~g�ᴟ��:��!�:h.:�N+�dq=IX��̷��J���W�sw�"�ǹ7'�y�z��-2(��-��Vy�w�=||��o�@wHk��IE`�'�]��*��[��7�.^�#�Ǥ� �A7�DY�W1�#eAD�Y�w�Z����O���f�� d�і��}�cY!7�8�jY�|m�g���1+�κ���ܽ�N�N0�yC�BCP��.�?����|d��PF��8���Q���Z:�l��쌮8�.��906<n���+�l�Q`fX U�DB6�������K�}�/����fss��7Esc�It�Ƥ��;��u�-�Āxja0	�cD�P�`X�Ř�V%cD-��(ƞ������ҠD̝P�#��z�"�Vn��2��5g�����[��wnUo���Z�L'�GB	�\pC!���p�;������� g�^�r���쮲�G��=|��/5X�1τb����!~��t=����sӾ�KP�lv@�������Jd���d<T� �/v����M0<����r�:]u��GJ���؎X�-	�������0*�!�D��L�a�J?�ߓ�Ebq��+4�VY�����Hɲ��l�Zi5h
:ݫ����z�κUS8��#�i�K��R�冎s�¸��Jq�>�Aa{���i�%̂�N�������Y37Y�z�Y��M�30n�b�������?��L�'�5#{q�����{�owTX]-G}��"��X�,"�5��	t.%�u�����ۓ��ߘ��n��&)��
^:DvTǒ��7hl\ �bȂ%*!&�?�R�W	�#�!C��F��86F�|��-�\�\i�J.r�}��[6`�Oށ�$����|�a�1C�xb"!���t�x��阵Mw����ݻ�;��^��6����B��/����7G�������yx�m���V��m���s�����r����G Ȥ˖"7��:��W�+Ǿ�x��m�Fd���؍��!�H����ñ��fGg�o�N//���fܻ�y��^�)�Z3QW�I�+P��	�	�	����?C��~J��$�W�ȔX���JJ]�FGJ_�%�'�D�|I5
K�1r�6�Ou�$2=)qz�]dZ>�����*�xy%�7��Z�H]�_U�'u6eL�KY����'�JySf�%�JE����.��T��ڙ
OE�f�O��W<��d��>�����I�ĩS)�
O5���@�di ��I9Z�^�O��L5J���SO���[J��F0�.iLmomN�$q�.�>Y�����' �իW�~�-}��e�-[�h_C��ʗFQ���T�Ȕ Ջ�����Q2���=�I$H##��`�%t�J�&�M�~�xm���� ����/�tV�$Jqv�jR�:T��[J�&g+����c->��J���6�SS#t��O�g��&�*�u��ϐKs5���P�L�)��>��J?e�-i�d'�:C���S͐�ΐ�SiT����HM�L?=ڦ^�x?(����>t�a}�L���KvehT�H!�Y�Qe���0NK<$5x��a�QRƔ� ��$|d�E���'��Gh����B��ږUmbh^, Yb1N�R�d)�wj6����~�>JM��QX�*��%�O�kVdԒ
),2%S,T�7�H�ț4bd�B)ūBz����@��QX2	�����Q�4���T~j�x�H�-qj�O7�<�a��ҀLZkS_c�2��-R;�U����VQ�-}R�'u�[�
i �Q�Vs0�-�n71�#�E��iu�%�Oڮ5Z�.ۅ�Fy�����1+' ���a
�nD���al��M�94�|�� O�S�]�,�<$��"�.�H�A�iv��Er����Vda�N\"�D�^�a����z=��tt��Э�>�3�Lΐ ��"l�8�X8��uI���@$-���[䍅���i _�O҄�[Hu?�0����l�)�h�nY����=L��j���I������[X�78�e���*l/�sW.�`���N��\W8)�dN�v��}�qy� �w縦�} <9L`���/��&\MLY{�0�q�<n����1�� 6���.�������9����8�5��mq����O~��?�䣽;�j�Ⱥ���q�;WV����������/��M6���Pj���D�lj��f.
�� 5�'����H��c�z��¾*���-�h��h>6��$��2�i���E(acH����<�ݚв�Ir�(�)2�S�����m���n��Ǳ�2�<�WXX5����usx_�����~A��e�w&Z�����
"�M��o_��{�>nOfq����Fb���r<�\,!�Sqd�[�-?ס��04 U��
K�X��%�T	�D�~j��<i��8M׾>i���V�Ud�����Φ$.�Hi� ��n�[yg�}vt|0pLw�r��,yqpս���j�h�Ə��?�yf@����>�$�� ]NlZJ��f~��	&#�\s���+��o�U�a�CSV;K�[� 
�n��@�����d�2����F1�/zNbn�Q��?��bH�ݛw���pu�ġ�^�;��@9��;��w�U��	�xe@F��<��Tk8/�'����'"o_�t**��(7�ڡ:�H?�.��\lTC��O��ʮ�c�
�f��-�i�����9 ��c؜I 5�p��̄r�M
y���,ӄ_t͍X� ��R�:�pq����h'�nO>��L7(y��L�S���cd��[���H��_�~���Z���g�ߟ]�mUKBV��F΀�"�]��rY�_��n^��	�:g`Em�X��G-q�+�)eK�7�y����	k��Y�VOJ&�ݒ�%����,m
�Hw�C(i���GnԾ|�5WN�n5���b[���@D�7��̣P���E$h������ݭVM-�ڌ*\	᪉M��tښ��`�y��;&r��?P�d�E2A %���Q��2Pe;ca���������l�%���,��|&8$���p5pR.(���$p�Rz����O%�Q����3��B���8��X/ͯ0h�G�(sh�2�A�_��i��Yn�i�/�u����[�l�Vq�oe�1k�j+{w�b�N�q����E�Ⱦ����������7�q�QX��}��VА�A4wI]�О��"��+ӹ�3��L�`�� ����BX�a\�9��õ�����Ο�^�f��V��|���0;���8Ѳ�����p��'qF��Ѱ��Hp[S����$��d�/,�UU�LXJ�-�����OXQ��	z�-h��jn}?�Nie>�Uo��Lz���0v84t��XT����am���߼T�U�ګ�p�ja�J!΋	�%ƒ`R�N�#d��U\jGr��XU2���&F��*���h���qH�0�\^|w��~�$��h�U!#�$?ÿ0���s�i�՘pۨ�0����;�&��%o`�@�����X�:8{|[s�f5���JW:��Lc����m�pzO
?~TlV]@�@��%7���=4U��#)�
���$���b+S���ĝ��	lB�`�t�ɂ��cV�rƭ#��-�L܌b��p���7��4��ҁ��7P;z9�,5�� d�N�l�����E��3�}�	�DT55��n���2*V��xRQȘ�>I�
L�����x�T$Z�a�������A_����h�tk���7��	"l�����^-fL��u+!1%k&�.�u���khr�g($�Ћ�6c�1p�8��6�k�Ƈb>8�X!cD�i�/�=ce�z5��SN>cs�P�HN�燽�8�������[p������jp��1
C	���}X��Z�b�g���vc{&�^g���ޭ���}z�<�C���G/T�ĳ�Uh��y�0�6�wX�����6���i_pU/7�{�b��թ�+~מ�(Z��:�Yv��e�g� �A��4����0�J����qL��H��i!ph:�R�7����R緰%�g��j*]�����
��bB���-������W�߾1�w8�'�I&>"�a�nv�4 AXc�"5	G퉞�!�$Nm�Nx� 1���^O��vj���;Fy��Hi��)�fm�q�G�1���g�������zW��������?x�����53�!L�]=̛`"k^��1X���T�W��J����N�A
�Su��iD#��=�-Ayi�E,�KG��Ny?����
!CX,��m��Bg����;HH���q��4������ni:�L���/����Ԫw�=���(�N�R�z��?���w���LC��Xc�9dX=�@r">8�Wt9�!�=bjg��xDI��&�6�=(�H�%��ġ��f`x��)���Vs#�&/�/j��;"�&.~(i��Ȭj	d0����`t��tF�F�zf�Y�i¦��Fs�o�|���X�ܦf��e;̀�6��N(�XQ�Ya�[`8zc�R/zVN�gd�H�d�_��OOg����cs��<�Q�h��mQPŊ��9l��"�DI��I�������a����M�hN���I0����M)5$���و!���/]���7�[�n"{��o��=b�����r
�(u(�B�H�[���Q/�Wky>c��3��Yصш����(dµ7��23��׶�F�^-�j���3�lJ�In�oBL\rn��K�Z۳M�����O!�t�]>�%$�!q].گ�\��'v���1�^�Ȅ�R��IJ-�ֲb�;�~�(��:��E�2�M`Oa)<���?�N2�^Oi7I/��ޛ��d<s��\L&29�`׬�G'o��F�}��E����a�
��d�V�fď���q�����-���[<b��hm���Z�*w�d�
�6f�aI�ʀ�A	�3sr?³=�&yE{쿳����[�� #@ܿ[�9H��v~��f-����ߑA��P�Ŭ��jg�=:m����z�ֹn���<bR�2�h��������o+2{4$z�-+�b�c&�xO�;��d� �L�@	��,�b�� 
&�r\�~�w���N.x�/-����T:�� [V�*�-��I0_��\�^�W�Ew1��b�f�-B�
�ϯ��o���O����k��\������|�]6���;�և��G�3G�=�f�TV��K6�����I:����9+���@�*�:��k�֓9iɼ�e�ѵV^v��D|lM�=L^����cu
uOOb�QW��sd1�� c
�4���)l�H��GY�x�E�b���5�j��b�/�*��yRv�R�靪Ki$���#J���"�f�Ha�rĀ�6+G����k�O��xo�ʨ.op�NúTrjO*JJ�|���"�Fai<JH�4R^a�I��Le�)�=� ���©#)F�r�L�իpi�4�(	R2a��T�~I��"�G�<�H��aY��O)\i�2��������O%��i��	+����m�To/^�888I�GС%�©�fnk��$ j��C�Fl��2�g�HU;B���p���0�^�޽��T��կRQڦ
�\
Q����\d�JK����|KH#��{������k�$��������Z*Z~mJ<��4��b4N˔�q7�+ݣ�Z���k4]�rhn�D�E4C���ki���bO�<�tQ�� ���N�P�h�����1��N��bŤH��L�ў�5ի4_%�)�O�R���˫�(+K&�M8�H�Q���`��`ln+�WN��@�T��ҧ^(��d_� �1ީv0W�rd�K��р���i��o��XQJ�Ӣ�$ئd)Wj�b�B�9U����\"�=*�%;�j�}#+ F���[��[LJ��%V�\�Լ�l]�I �'�)}*�O�G3䅖�m�
W�I)��@85^�J3�UG'y�\\/ؕ+�!)�ҳӷ�aw2���՚ߪ�7����!l���P�p����	�"��� 7T!�D�!A����S$��i1�wL���$R��8�9�Jq�A������%(�W���Yg:�	���p�S�n=��<z�Ęԩ�z�Eb�*{�D�%��Ն`�=�x�ϔ�fR���] ���%0�I���T���b�渱�����W�!�em��S�9 �� �) �HHa��`č��i=W��/f�E�E��� P6:��f���Q��l�oֆ�F�	tq2���`�nw����;YBH���,�����Q�w��Oۃ��{���7� F�|}:��=����g�û����Owd��jC	��D���ݫ��_~��g&K��[��	� yp�4R���.k�@t��F4���#���ӈ�*;_�a����)�]��85z^l�z��5nrH]Qv��n%a���E~\��N%��U	\Қ�K����͚y-Z�|���4�����#F�./vVD��O�:��:=ꜞ�=�<���.o9�S�%7��8���p
��&�5�sv��O��X����h��V���2��Q'��1�4F����vyWL��Fϑ� ��M�s�X`z�g�l�w7ooo�z���/G��G2�Ba����4���{�喋���ԡ4rGqڣ��O�ba̂=��3$Ϗ���z�DDf3���+N�X�L�ܦ+Ciz��(�t�Mp3E�~��t�y�r�Z���?�_�]���R��S������C���0'�ЧD$�3JB����a�l�I	�Dc�G�j�+A�JK�\��RQ�!�"���@W�R��R	�&l�Uz_��7�-����C����b�Qi�(�)�P�O�t��W����f�NJ��DCܐ��[�j����F}�\��@��kq�Ja�kW(���jk#���l�)���ړ�����O�FK��V��ɛ'�/��`#]���%�kgQ8�*�و��@��g�Ň@R��| 05L;ċ��Jb �|� i ��҂�O��c�u���ũ�ZCk>_=>�{��{�hc�*��fa�^	:�
+O�gf����U�-���2��Ԥ��]�l�)E�e��Ν�7���N	ʤ=���T��� D!�N���q�&�o!a&F���K&	��ڣj ��Wl�`=�x	�"��@z���CFZĀ*�f|b�C�Qv���/$![��&����������jD]C.�ӡ��k�p�7�\� ;N2Ul�Ûg-d�hbfH�����@��ʹ7�>�������O�7��y�:�n�q�[j	��P��
`^����d����P6�h)!���ѧAZ���F�g�C�K�/��U��e�/N^��N���f�b��f��c|X�t�$|M�[��h���i9� X�@5!�H�H�xdL�+l�|J���;R�ї�u*�րj��%C�������T�A@^�|�ɽ�Fes9�+�]3��=��h���b������<���t�h 0)Ԇ���"�%6RF�5�HȜU�ӓ2�F?�Z]Z��[D��K��C/�� 霼���G�j����|��p85{\�<��2��s���d�l�A����6_?�����y�̉$P��:�3b���i �4:YߣA1�؅���,RzĀ� j�FAXJ��(�O�Ea~~qb;ǁ�?��w�C�    IDATRF-f(p���)���)��(�4���
�+D��������2Esڌ`��@"�Y���� N"2k1F��8 ���	��H�=����6���Ca ��(�2�S�aٽ�~i	���W��F�=�mM͕E�Wi�p�IX 2qz>�Z�VO%�B�p=�}8��Im��9}�d�Τ٬4�<�P�Į16j��H�C�Hr��m��
���Ķu�jAE�I1�A.��t0Ӓ�kP~&�B-��G�x�X+u-_�]���%�6�m&;����|�߼9[�0�����)B�d�f���Db�>"�I��d�(��>i�nުG�CW�,8�u��q������&�H��yg5�� �K�Gg�w��������������;��2K��pvq��j��$v}��J��8���i��*L::@ n'f'x�0ó!�t2���t}Rm����>h�4���)��������ۈXV�bC�Xb�M�_�a
��1��Vʖ�^3d��	]�����������4�wl�.�O�O?��>���`I4A���a��6��`V�j����nI�n�.���/�6v*�M���'��]2n�A�N9L�ç���vΎ�L�t���Z�����fn��]k��k���Y�0� �i��P&�%��!$��=�0,M������h-W�������^���i�J+׸"��r^�]7��Q����7�F��$86���D�x�6�B݄yy}5��]����/�[��v�;�Q�����������p�<�	 g�@�r��p Iy�����@#5�'�0_������R���T����GᲤ��+���ދ�|��'�=��-�2�	�� �p}
��~q��C����s=XYp�;�+=RdpW�����q�9^H��Zp�m�	�
4%�Ά�,�l,��u!� �45�?0Q�Ê"��nopu><zy����ˋ���vu��'��ay��R@�eу[4�x7OBc��5���f߿�Y�W�x��H�=>h%z���3��Q�! ��HhpT�IPF��(�!"w�ק'h��J���u<��nW�	!�$K7`,�����P̸����S[�PJ���s��a��@�$���"G#E⬣�{�ubԍ��3w���ϰΎ����xXa�l��/���4aN�3��,�����zq|:�O�='5�\�� �	nTMC�i e�l�!���2;�(���&�d�si1>x�)�h�Ig��)M�ɚ�g2�Rj.ڇEP��v07���u�ۯ�'N���P�8���^�:���լ�g��neX���'�چ۟&�-b���L2#�="|�O(��b�n��3�W�Y�Ɓ��b6�����A C�U��3��Ko�]��ʕ�X6��h�<>w|���wf�H7�x�A`��pe
��:b֋Io����j��Ha1{�PP����T�r�L	P!�z|/�NF.�ß��7J�wv��MC�2���g%�e#��=,ӣ�"#c��r�n������fp��F8�/��e�W��:�Ea�/�/�_�w�[%����}ޝ�۫����Z���ϸ%7�WAs[�rl��+x�������6zxv~�C6 �΂^ԐAIǅl�7�	'����,�J�N`��dQs&���$�+- ��T��^'�� �҄��3�G21�)2�SuҤ�7�}���WK�H!�"S3d��;�h���KkS|��oJ�IpP��O��%}j��,�4�zx%�2S9���N)��O�y��Z
+ē"���S���i��Oi$PKԝ!��M�O�2�xE��&��?=�_2���߄uP!)���Rz��[v�h�	5��\q��+�[-髀�� � 0}ߋ/���Tlj������la�Sxj$�0�Q�)���J��$!��J�!��e��O*�;׵٣LmP��(��F�"Ũ���/�%�~�������!�>�����{�&�cW���soE(1q�r����	�&ՠZ*�@i���ÇT�f�Hp�A�Q��行��4�o����w�UI��L��3�+	�����<ɥ"?S�����
��#��*Na�Smtyu6��I�G˥L��S�#,��b�W�{���T��@�_ ���ʗ]���i��)!�˘jOi�J}�^L�T-��l6��Q�#� H��r���L�Iե�����mJK����T��z;}�@��Oj�&��J]P�M��
�� pV��T~��F	���h��'���M��+ALj�4��L��q��QjO`�^��J@bySw�L_�hF�!�KљU���9f�z��f"���C�!\4)$��EKdiB�p��}%�C��� R��D�s��OkmX�Ł?����=��pe!��u=�[������wr�?8=?���&K8[�MW���P<*�dR���'O�EL��?E�:�ypp@��2�9t�$A��-�,���O�iX }g���ȩ�l�B�]�oݾ�<\�}"�&]�Oi6����ȋb��+��|p��b�L��-X��}����x-<��( �Q0+���m`z�2�p�f���p�KB�S�G�^�D��熧���!��ƨ3<z{�峣��_^N����mZ�dk�]V�}�?��_��_}pw#|�)�����јј3��۽x��W_����W����g�4,�Im�h�z'dN(�'�J#��4@)}�"2e�W�Mb1��x�(Y	�=[K�#[N�	��W\I�	_�w�M�����1vM�9ǒS~�}�k�|a�Ǵ����Ph�����\c�"���r�B|��c��@��@�F�q�rй����u�|0/lmַw9�$G/��(EŹ����P�"�Q/W]�2�0ZW�Mil�l	2��%Dl2H�		�~�p�t�F����V��!'r����6H����������m�[�'W�N]�/4�&���EF��{lF�V!��Kr���B�h�Ｗ��.���g0�v�p-A)Ɠi�a����l/(���sS&�9�)�-։���F���؜t	�g.�J�ȕ�(|���C���B'W�/�yu�f=-fq������N�?��7+��?Wz�O0Cf=��yi�0b�O�H&K��"Sv�qH�d1
)c
��`LU�I�d���')���p����`���ࡰ�Z�rN�*a�&7���_���\�A"3:�A��l�3��ʏ#k4���5�k�"�5�EW;
�[@���9�jB/E�LF���g'��7��^]��쯛�H�Ц0TC�c�ҷƹ�w��,��J�b5&_<C@ ���;!C`T�=>xX|�(W�7���X/��I�'��4���A�Ϲ�@N��%�gK[��\Za�ʹJ=��3��i�#/��d	Ek�:8��1��\
�Z�@>���o�̈́�#&�e��lab[k�� �W&�*T����LOo���o"��4N�y0�ݫW��:l-nSOa�΂����0\�d0?~b�)AelOZŃ0��-<�'�4�ʷ�Aph�	������xo,�U��8�f��]!�ζ���-[�*�F�� 8���1��L�Z(�`@,x��!�2h1a��? �<���f�~a�d�f��u��&�k&G�!�W�ħ�`!��a�3p>0�������//���ߝ���?~~�d���p6fn-E�'݃��{E���iS����ao�ٯx݀:�T�#H�4L���t*YFC#�Mᦃ��ᠵ
j�O�!��r�8������ �e��VfǴE��3k���j�t#��\���>Ӳ%�*��(+�+�)V04����QD?��PM��eS[c�&E��z\�9�y:���}�χ�����>�R�جe��?�0����p��lln�Po�?,� ���z�b"��[dr��A�:�M��SD���3�T�͠OryRi�P�G��]�C��]׀��� lľ��؂G2k��W�S�h
>��
�nAj2��Us-�����u	f��f�f�����t q![u����>��kc���f"&�!��W�B`���~Rj��蚰%g(��AylxӾ��� uʫ�с?�9&X)S�*�� ���D�c����yRzi�:����8X�s���RsV���'q���v s�lB([��g���pzhKfD.�8c$BVk�G�b�{G�4�^�,ƹi7F'�,��(ָ�QmȆe>��6�iË�g��?;�Ε���6�����v��2RaQ̈́�x�O��H�31 �Y��B�#�X�yE��p�>9�R�Z[<p�2��(`��l��� ���,��bNf�9��x9M��6d����Edў���`�gi�R�D������p�
�b�Ik�:A"��6��,W#G�*N�b����v}��\������#�ӱ���*,�RՍ�K�����8�Y��]%�ϖ������o~�ٛ�� F���j�/�$���ߧ�$�1�c�^���7��/�5� qXv��g��~8P�<���X���6^�Ʈ��V6�q��	*L��O@���x��*~�瞙�8����h6稐��:���ޑۨ���B���TJ#H�M 
�Z}��_��$O{��c��e?��'�դ��b5�7��8����̎���J��2ۺtՁܰG���X��X��-;)�5nvuz�9�O���N�����#��KfӰ�o���_��_<��]B6�bnAM6"�~L���8� uF�A�i�q	����13�Gz%�'�ISJu�;�%K� �p�	6QCpږɠ�A�͏��?bkt�@��C�EQ7ژ�JA��gC�T�r^x��� ��,�]�"<�/���tP�g����U�4����rV����A���Z�׏�R}�	^dGf�'�Wߞ�|u���b�h�To�kT(�i�c�:�]v��"�:�F����:��>�� �O�L��	upĲ뎍^��\w<#�5.��/�b!6��Q����)6�V�>3bs��5)�6��P���D��]qCePX`��9w�Ȩ��%��8�	��ܡ̆�Y{�I���ɝ�8������j�$�����~a�*M�
ю؜	�������J�4�?ݤ��Y�Io4�v��/���vv��[x˶&C0�l+G�H!��݆k��a����d������	������br�\��ԋ�t�b��sc�3�dp��Q�����.`��|_�QR�����V R6�+��΂��JIL�=�<�����s~��ru���F���̙�$Y�ni$�����;�o0�x�{�mɒ:��L�L�f��Fu�W�B��8@!
�B��{KVv�_��Z������'���n>{��r����Uw܎�㛫��%3�'�u��=Mx.��8�{�����[v=�����g138�|�}���326��d6Ta�>��B>�Yc�~��a�ꀵ6�C��8`\�\��o����$�T2�d8���[N�z;�rqN$�^*�@��L�d�Gb�����ק���e�u����������i�6>c$����S�Pn��ú��3x�˭��kO��z��꺷�e��ul��c�vtۍW4.t�6���md�4ꥲ����IkۣY��h���$���"Pȁ��<�5�O.�y�{��]U5$�z��T8�°�l+�|�r 9�j)��d�&���4��⑐@V�r��7=ݜ@0P����e�X?+79��$BT��$�k��xD	/`_`e%V�0�GHQu%���j;m5_`�X9�#P=+��*�2�
��[!��+�@~ \eR``*�`*+��(f�'AJ(�~�L�m��'Ϫ���!VUC�����$�@*FD?����U��8	u0�8�HN���Vx��X�[�R�8�˧*cD�s ��L,�0mE��z����� #Oc��,�i`��T�l����7��J�!�?�!Ӧ�B�����s_Su	�d=F�a��r�;�j�'��"N�`�.5�#�=x�@�jP�����	�p�bI�)���>��O>�N5#9���O������y�VjѨ����2Q=���o9�+�܄�6�T)�:�` �p���kQe"[?�UX ���w�0�h'd��
��s)����,+�R	�3`_!�U%*k����t���*���,�e.p�����D��o��S,�s<0����U�K%jYU�*�*L�¥���q�O��Q�[��1˳��W�$����+i��PBB�]I!�^�jĨY0�OѪq��X r*�*KH���y���F���%wOB��&+�9��=:�8�wsE)��\q�i(����x8h�F��v�Z�9�I���Q[�����@BVTV�[ilV�$G�g�Q�D&$.���ӣ�������/�Ϸ:{���ŏ>�ȭ���5mq���B�����y�;ȫ�h����O�ö�͢�f�H ���a0 ��R�����X9���\HY��G��+x�_��j��X���N��r,5'��j��"�����RS�g���ٽJ��)+xG[0X�D3B�K���B�jX�T�9[��K�/�-�es��(EI���&�ǲf>�>8tI�����_?�͗o��oM޽ww���$������-w:-��_�������������Hcy���p����u������ӧ/�p�bZ�VU=�Z,�j~�,L���j��a9~��8T�Z��������e(s��M�	��K����4�1	�zƘY�x��6���*+T:[D5��є�ZE�kf�X::��M���؅X��'����^"XӢM���k�9��m�|�d��αUn�,�=>5ԑ7E��k��$���n���jf��l� &�v���(�
	��c�J�ȷ<�PX�8��@�	ZT�wGx�J/,�v���A@֒̒ɺ�1��G���v����U�ةב����5a=h���	sN����c����D�>�%����
rq���:5�S�&��5=���F���K��$�/P��~-�oM�1��ҳD��'c�昉���ܲk{��ً����f�r�e1,:T*��������CZ�&�UQcQ�/�ۡO� i�bUF���^ sR ���/�4������)���e"YU�U*~���E�!h9�������H3��)�"a�S4e��ҡ�J������&�`��rݣ�����$UeB�a,����8T��4D#bW�]6HЌ�{������<XY;y���>9��z�_4A�����p���B���'g��n�]t����]f��+�����1�n�1PȄ+N
�C?���S8�����J��l��W�i0����
L7`�"tX�{���Sc�do
t��	"*���Ly	�d�Q1\]$�8W�* �٭O�r�	���N۱Y/��yu�-Kl���<kFg>J��*��'I�Կ�N���ٞ]�����8H��`ԧ���!�H��ȍ0�3�KT�
���4j۴FH� yP��F��̑�!��s :
�7�z�1=�2e˽=��jXh?>�G��/��˹�����0��n6C��WT��l��'YxgډNF8��$H���c�5gJ���sh�>�&�<TB-�����n
0p�(�r7ݤ>v0#��~^�����Ë�����M3^�����#�������>|�,�>!��L��a!V��Br���꥛���7�>`N��`�G�Y|C?
�$�*�Bu4~���|���?����
r���E�>1�c�:�XRz7
TM��K���R�n��}�N$�"��`;l��n2^�
��I,���m+���V��&ɐWx��L �?��E����<������qmO��/�/7��u���\_��m��S�(+fM�D޵ڄX�d�^ԫ-P]b�O�o�����ķ������5����W�)+�B�L�o���g������4B&��$[������p���$l��I� `�d�`gH��w�2 Խ�jeg�$����љ�)}�xlsa�	�59    IDAT�F3k,f%!w����%���*ZE�����dI�Ux�:�ݰ�� $S��-�1�^SW�*�������S�$`��'WC��*EB!��_c`G���4���s��1wa;��L:���)�q#��ZA��1�:�$�8��7*�\���K_b��5�:���&�E���j`mU�����>��!8|�2��q��W�;O���룵�ǓK�@,j�-k��s��͵����>$p�'�S�)<Y�H���V��Q�eru�lj��5!��4)M�ė��U�2�g�ܤ73;���م����G�2���r/���&�4��Xܽ�M@���8���fI2�$Ʀ�:F�OiN�c����J��;�We��ё
D��$`u��y�c!�a�~�ID������b�����Q�����I��׿���}���w�󇭝mdC�C@���G?��S
�b*�8L�6�'��K_f�,���]�jR�S!��s�-�=���\�?ㄓG.�G�q�\n��\�n��(�Y�QR��N��ي�A/2߹G���5�Mۯ�7 ъ̌gӮj`��k���̀��A1Q0.9@��X�iRs4�v�����r�P�T�ߘ"0��s"�Ve�Dc�L��;�"7���D�"s�����cw�s뫕��ν��O�Ώ���5f����}������������ˬq~�T:ep��g�>y�׿����p5�#��0�,����7��V��K�[u�B3oX4����; Ӈ�ygf\��"��Ii�O�z��Ad�"1�^3��E�%���,�{���w� J��H�g��r'po�a8��,�p��>4�Z��/��/DG��Fn�Rf�F-��0�/u��n�.�=�z�ѳ�g�;n�Xp���Nc$��g�F�h���l�֒��6��Zʵ���~k�PM���Idz ���K �h����� Z����ߜ��ZG_��#A� ��Nv]h�G�\�8w�!S3�V	0�fXw��ͩ�1�Mk��m�HF�Xˍ�T��ÕN��$��ݺ���,���e�9~59�b	/�XI~��q3����[�W���5ӓ���;裥��������κh	���9]72�IR`PM�12?7kWT!*�2?�j֝���T@H��\EU �������Ƽ�����:�	*���6Ho�7A�{"��}UV7e��C�MVJ��@(�k��?a�qW���Y����v�V�R��G�s|v2��G�b����iw��#���h��Z����ˋ��K�͡M��]�of|b�B�Z�]��ty3yv����������sי��ʋ5Ko�B�{��7T�v_d�'�&�9<�+�.�� �by8����jŕ��� x Bp�
�DO�S�@0����1�s��,���Y7��<UZ���"7��9����eiϥ�uG�v{E8�^�K���/�W^l�=�Z[�Y���x���b�����+;�/V�-�nl-??X_��N�v"]�hvɗ��`d���|%Zf^2�n�.���7}�JXĈ�\�gB�A�5�L��쵔�1�B*��V�[?}�*���	�TH+Pr�r�^"\l���U���l�{��E�Y!�
��Xeq�
�:K%�OM��X_��,0?�O�Vnj�3�UJ��%��áu+}e������Lr�,�:T�*�o��T���1��MT�|� ��|� �a��9Q6���*D}x���
�$�:?�ʡ�b����W�p�~� �ȵ�-���}��Ǣ�>���|_	E�k0p�Ajee��r��j5��J����J� �
�'�p_+JB]��������qL�5�0���<�L�c��'��_JB��+�~Hn��,����
&BG1i�`���\� �k6~�!�����rB UcGfR����u���2��<y H��'�@#�,2�ӧb	�NdʼN�����x�QK(IW��z��0P{(_�*B&���%�D���&�.X~�*���S��j����r�m����WB���Y�����[n��
��Х Hȩ��C]�H.�W�r�,D�8i�[_��
�rEU���Y4� i��)*V0�(���U.�py�˭"|���$W ��P*�𡇿��q2D�R�e%o�"pe.y
�~�|��[I�L�o�#\e
�z���ȁT��
�)<�TTL}8Ł.��VH�lϬ�:��cYM��F<=H��rX��v;�f]�F�{6�ŀ2)ۙ�x�b�y�DAsh���L�d�0a��bIqn�IR��Z�99�
_;m�%�eZ���ln�//o>Y=x�u�u�ډ�{����;Q@g�Cv<5���%�?��w=���wޱ[Xsb^�t��|a��˗���jw��P��fb���髺.�GH9=����A���ba{��<��v�w�҉��ŷ����%�Dr'8m��1�^C��MKQ]�������(ia.�G�}f2�j�A���n��eU r��f����A��k���d*�mO4�z�F#�Y��wv�v�^����o_~�r�{32�M�-�Ff�C.޲�߭!����_��O��G�;o早�b�WQ���w�����G�����o����0!��U�3i[�:(%��1��u6xa�Y�0m(�q��yID�S�_~"{���{�W�-)�E�+�O�d���&m�s�\��UϺ]�Ȁ�C��*֊��?zE�D��*h��SՃ�Zp�Ÿњ�����v!oo���X=|�����������y�4'n�$�Sa,R�'ɷ�nb����Y�1VH��\�Ա��ה�Ө��Э|
	<\q�
/�Z�̯�X[�`Wg��dȜ��:�iTkaR+c��@�^�3�t����
��`����)����ft`�36��kws�"w�}�c�g�;v����	uY~��u�ڀN���[��υ��8I�����u�2oʺ�q7:\����m����lm�o���wӯ�g]�c�Ђ
46���_��s�+!�q<�pk�E������,�-��?�m#6Q-�k]��!W ifc�R�@�d�[0B�� �0r���ʭ_��Pȍ^�+]�s?��p�s:K��@t�v|�Qv䁺�b�KP�S�|�M�������HڗY@�~��y������}�lw}w�=��Z����[S3k��Z�p���e��0g��r�΢���qr�4SŹ�聶��n *������k�T���F0�\@!��?0_xK=�ȍa�y	W���H(��3Fb(֜��g'�����S����K����!��#�-8�ä¸���dc��':�Y{���3;m��Je��p����Dl�e�ϥ��\�([A�$L2-�F�6����ΨIL�+�T5�W���~IS $'RD�H������_�]���K/4&#� ["8��{^1V��Й����qv��C%����,m8Pr����<��i�>�;����<0;w'O5�Ș��I�PV[�������������L�2Q&�B˨�,&�~^zU�2��6Tq���1^���͊���z����������~qp}��w��b�Wv7�<��v���seǋ=��;Q��=W�P���������gh,�>S�6�y80!�Ǝ|�iI�|eX�W��$�@)U�p,������L]�Ntm�gAI����&�C&\>�b���i���6��9=��ht�!|�0�̭|�?t�����+Xg������c�� �Dh1]:��
#G��d��Ywp���xy��/w������_�u�k9gd*�1�F��>81�-�ss���.��Pc��*6�s~0PTX�T=Ӏ7D.� �Hk�pPJ����V0_A�\A*T1y��*�����$Es�#��[��mf�d���2�g7d��(��3wA:^�����a?38���>X<������q�FwY�[ېq	�Y6Lg�#��q����_��_/^��.�-T�#���B�ZAW�'  l�HX���C>�~y��o&M?� 
,��М�Ma{��8�C�@~��$GFQ�w�nd��-��=�T��_�8��Q�n��=�n�SCF��f:�SmS`�r�<�t��s~�-��3,�j�fl�,;%h���9��΀6�ʬ���i"5�	���N��uv������f�|������ C!�Haؒdb��ld�6bKt�g=�� ��<@�u2�ap�-���f�C)�1�Ǯ�<R�"�<��=c*�F�DG��n�PH���������ƈcQ$ZLQ~�Nè��L�-f	��-����;�	t�d��`C��Ëg� *H&����9��9+ �6��3�Q*c/�L1�р�aD�do�F�=��m���)u�~w�`ss��omln@W)��Yx���N�����կ>��SQ
�^d�ˡ4䍶��h�ȁ�ݢ��i{J�W}���<�y������N�N>�u��L#���D����oy����dp�Q%[���:w^ڛJ�9#���[�SD(4GI��]��֟�m��oٍugֳL�`�4��}�C�_	�>�]�}�<K��:�ID��	��~����22������	��æ�V�[G���Ñe�5���3�e:;�"M޾������~�÷�/��`^f����"F�7%u:G�Ϟ��4oЋ�ⴭ�v	7Wl�O0�\���U7	/���q��}[�|Qj��k	1ir�tF}a��_�d���a�X�&�B�?�����!��B�؈4z�Z#�/Ӧ��E�� �����>���Aqh�/i��s�e��̓�_�<[�X�;��so��}�uwv��9l������|.��
����5 ���PQm/�@K
m���BQ��S_���ሦzKI�F��9�g�>g�A3gHo<{1Cf[k\8�iV��Y��*�"�k�&g�*"`<[��(}�ZH�t�,����nBpj4�Q!�����`��?�g1�6i�l�g��\(N7����|��*�P3��&�~6����Ӯ�t����`y�d�x��0,��\rBw^���~j�n�)�P���]C�Q"MU�*P�hXQ�A)l��c}�˼���)��C��\BC�1���Н�����0�'g�v��fK�����̜˫�tp�z�-�T���xu�'�ʵL=�������{��^=�"��w@P�CC�ވu����]m`���m��A��[erq(�7r��(c�)MG��.�=������5���'e].//?_v����=,��V�b�X�3�-v���p|{�#%Lr��䩯�Z���UC�G)B�,H)��J"�q�p�,2,0��m�8�^�7�"W��:Cy�!4/�O��My2�y�fCTd��+M��	LS�9�G�O�n�w���^��\��ߜM���֛�$�e;V�;Nڒ(T�;:��/� "@ݿ3yM�]��D��P���WW�m��dI!2j���X"A��@MV�b���n�I`Ѷ�
3yJn᯴<��G��r��P���b+J�r�*��+7��s+������,�䢄ȐG���mH��e.�L`��WZ�Լr���+ɰU��l����S���&p�.E�a�Jl�,J��3W�$�X�S�I��)Q^��瑪��-�*�b%��f��!� .����L
r藉��r+	O�V�و_l%�)C%r,:<x�_ͬ� h6h��� |���fp ��Vlr�Qm9��O�=����hTD�y-� H�'����S>~��vW PsҸ/�d�O�QE�ydk�%�<{�Lѕ�/�Khir4`��	�Ѩ�J�p���ag�9�B��dP�_���СfpG�b�U,��S�B�ƀt+�M�P-��D)�P��&������������������^WFPuS.���G�����t!��G��RI�ܸ���v��&U�W�:Wr�U!0&!'J7ȼ��.-Xy�� ۪�(��'���!��)g��n�-'P%�U��d���9�U%�`d�	�xD�O��P`�T8�#\�*��-R)zA{���t�2䯟��3�L�e[d 8��氯p��X�(��y�j�W�@�<�@5Q���[��!
�eR������+-�XI�V	UϨ�Y]YI�&	�ʹ�ˡZ�g�ed6m�VY	�)>�pH�2f���O=oy��F�Οesx�S��A�c��f#���2Zq�+Į�T]_tHќJ�?�鳛���rﰻ�������y����:��yn���{�	�M�E)Щӭ0�.�~�������N��>��	�Ѯ�[��[T
L�ܴZ3�$�T+X�)��(HebXFne%Vxᓸ+�����i9�i�B6��q�u{���L�}�-0�<��pe�a(�m�]�=��\/������3�Z'Q0U��A��mGH��r�k�Em��l����ȈǇ��Qgww�K3[;k;G{���9�.���̹$�9Y�^ܜ�!��bn������G|p{�E$YR{A~cw������r���������y�g���"�N2�o~r�\����)�ſ���| @5N�;���,�F�!��K%W�L߽����N�r`g	���1'�H%�j�F�ũ-�.�`ct��M?�S��?�����h�Α����<;C�����
���U��ż�՗{Ϟn�x���/w������]W3�Qi��Ń($��32��3���y0��И�7��wz[���s�����B���d!����px0h�H]�n�"i{���	���"'K�l�EQ�[�ќ�{ad���݅�oM�M�9��¨co4nФ9�o�{1����>���Q}[�����[mI%�����!�:��nN�:�oO�8�Bu��ΔO�e�NGz��r��|�����+��w�s_[�]���+������9'5�ӟ���?�YX8��*�q~B�� 4����~���\0������m>/���L.<b�����䯯��pB:�D*�5����9��5$Ҕ���@0f���o�*�:��a>Y-�؟�	d������ñѣmԇⲦ��>V)*���
�L���N���g�����������᜽��tr���)Y����O��u�9lz&�¨{��F������L���T$���"K�E~�o��)	�ba���O�"?aX�R`�/4A8:��Ƅ1���F6͎�6�@>#o��ݰ�:��tp�YN��9\��^{��4�t�m�;)/�^=/�r�P�e<����<R%��⋧��5yvm��䥋"G�Y����h<�Rf�FZJ�2��<�<yBP&��AL�&#���9$�@a���c�f�\Ik�XkW4�0��Wn��W�IU���p�l�)�R`�Y��P�`������LgiW?<AA�x��)xOý��Y�p�˛)��ل���eF1�f�?\�d7�g�s���f6���n6���߮Exv�
���X�FE�d�ߦ��n��L�6l�;�P�����'kT�_=���n߽3�0��!7^q� ��C������;w��v�����-CP#\�-�IX�UHH�]JU25��S���T�)�9	���@���>B�����ϴ���;횫\1����A�옣S��L>ج�EӒ)�]�����i�L9�����c� T+�]�z�� ��k�I����P��g]��B�E�� �-�6=;�z�����˗����￬<^۹���\`�Zr�<2���'�i��
�h����ȿ�k8�sfuƣfT%s�1�C?�r0É����+���(7��ha�U���_.��Y�0�*�xѣ��q�^0m>uP*rc?�B�B�G,Zl�Ѥ_`$��M�5T�V��Y�G�)�rL��*^*ڙ���,bkQ$�$��-[�������e�tbj��J�Q�ƪ��	6�l�F`BPTs<H�tc>�� 7?E�)��\��ɮ�#�+OA��S��J��2T�L�W)�(k��tf��[ӓ��''��;^�{��w��G?2�=�Ě
��뽻<Dy��e�)�u���^�6���@�
��'�e�d>�J��4��!-\������[��3���Ŏۿ;O�n�鋕��xupvyﭥ��i/m�"8GgF=|�6bpYؽ��}7I�6�T�602�    IDAT�u"�a)pXL�O`�*i\Cf(V�U�N1�p�Q��v���n���s�aM�9 s� �00DfY��텹F��#޺�Y\���w�r������v�jd��N�*ږi�Þk`�-?��s�D��>�����(�M��.�#�E7�����x��y2*�! ��!�1ذȑH��1;2>��S�G��q����������'�����ҽ�[c�țl��0OiU�!J1�J�6~�2�-��7^�={��?��xi����j����E�==j żHɍ�]��2>���g���߹믗�cڄ�pZCL������-�{�h�w��A�;�D�ǻGg����S�w��f,�D�N���;��,l\�ܦ�l�B�l^v0�1������Es��?;(�0c
�}Măv_nvÅ3�������#�z=K��W.��>z��t�p�{�����٨�� F�޺���O~���߽��{U����Ҋf��%��i�6_aJ\�±��|���jDF!������*Ȋ·�W�Vr�ia�C�	'��Id{�A?��SN�"�>��־�Ѝ)�DK����mV� 1�Q��$m��X���;�Aq��Ro�S�a2E�#����.j���=�B� !�#�sxd=��_���f�әZZ$�b���d�m{Y��fÖ�W�)�| ��/�����=�R5�n�맲����`a)�n�RP��;���m&�x ����à�G6g���Ђ��-��t��g�>:<ɜ>1�w[��0�HRFٕ���&�q�+8j��l�Q<&>���E
$�b4�,v"a"��.niFk\1d�ۆ�A���C ��u4$��ҡNtv/�����������ɳ�'����;�5D�C-o�-u|l�](��6�&#.G;��!
����������ϋb�*���[w��D��q�lp1
nYV��:�9�=��d|��۷gft:��WRI�T�cф��p6k\��Ze����_L��/��T`�c6O`��,�Ɇ��1fV��wvz�{�VŲ�I�<@��b�ʦY%NF�9���"�X�k�Ú.������������8$8dvK��ttV.0		5~1vK!��C�5~	��@ �i�
^�OYU�6r�|��p���p���Fx�����9-̆"�^��RDk��?���w2�ВLC|�pXon �X\9}�3���+tѦ9�.;
-^~�ul��`4�ϸ���P�-�󬽷�o,le�`�'��-���vRK��GQ@,��7�^�4K�����8�S�=�����b�P�'T�a[��_��by�`�~r���J^����$��_%㑪r��S���
T�TB�\�P0AtKU`9!\�Seշ�!��	Vx$�#[Nx9~�j[�*���jB��W�j�S_ ծa)�'�!� V:���y �V?���U���d�r�˼`�#PTՄ��Q?F�<����+������P
�UO���}�Su����U��ge�l�Y��H�!�,�Y"�T�p��u0A��  E&��ZZ�����V[��,J)������'�`7�)�9�XB\����ZYY!T��U[Y�e���&��?,�}���
5/HYɧ��'�79������r)A��@��D���rb��r�X�R��WX�b*\-5����DB�<Ū�e�劀w�к���:*V'�UZZ��T*��p�\#��n���p@���9ia���Wh��q�G���
WI~���d��҅��(W��E�������$��L�� ��"����\�@�%�E���a���"'z]���H[�T�@�����(Dn~J(Jɶ~V89��W(O���)P�H+����Q�
�F��ON����Tcl����,��)U�L�\�J�-U��$ ��pEU`����I�����&���L����s9��f�����Q��OZ
�-��nk�}m����%�E�udP嬟�|�H��#^٣�o앦��n�K4�zg��ݭ���W�Ս�����;�;�ݣ.۴��o��t���$c�F�9����h�I��(g�:�ф��ga�pX�"���W8<p�?Q�Z��q�#bqI���5�(hT`~_�E,�C�"!��#jy��_p\l��|������M���[����)�@�0kgɛ[�H�v��ӼB�N��E�x�e$�щ)2"��䄵�D��3���f��tg�p�s��Y_����:�>vq̒�ʝ������=A�)��٩O?������?��O>|��<ə���� �b��	�V��kZ����Ɵ���g�V����(�5,z������%�EkDꂮ6�x�:4��[.�
�G�^( ��~����W�WL�JV<�+ȷ}a"e��Ĉ3�:ލ�+A��ƥE��¢ۓ4&�c�K�,�<�J��*R}ՠcm�S�gl��g��'{������_����g/wv���w��[o{�h�.�	{A��ۨɢ/\��K19?=63��ĥ���=t4���9���կ��&��B��Æ�r�FQ�d>��V� N?��`8Y}��ːm"�7v��=��3�
Q�S�LO�Ȉbe1�/O��Πr�4�m�͈3�p�I��ͺ��.c� ����ϰ?�z��I��ޭ[N�`$.C��1��NJԏ%9��*6kb�]Y�\�:ŝڥ�7�������x�s�q@sus���������3~�����i7uS}
w�=���i06�+�=�����ΨI�XS$H� E���O9�r�
�������) E��p?%R]#� |Q�T2U`�s+G@���W����3,L��
G��ɖ����d�I`���?uxͯдQ��n�MG�+zM����(��� �}����ӽ�������[���Z���=������<�:5MQ �X�	�u��,�6k�L����"6���''$ ����S��Qta��7g�����p��u�ˣQp^��.�� |�m�m8�VH��h9�7]$cƅ\G���R*�!ʞ��N� {f��{�?,��ʳ
e�0l(\p	L�Aؾt*EV#3b&}P�e�9yzi�w�;������!���k�㈑��Yy�Ԉ��0�3�� �� (T��?��r��Fr$iŽ6�/�ª� ��W}*g���jy"UEAZ�u�BW�^h�׽�.�2�S�$�W̂N��c��y�������'#�I6fK+,�A���pjG�:����}J��&�F)HS@Y��f�BH�!��9�-h��=�^`Q��l҂�>���z������?\��7˫;�'��s6�O�ήl4	5�J�>�k���(����wHV��{��!,�B�Ѫ��s����z$�r���	N�a��: ��X�R�)!�na��\!O ��'��}���������Y�t(_���3 p���U�nC���@S+Tn�:i"�)"ˋvg~}�"b��]�
���6ͱzQ�/��"9:��������٫����Y��_�~�|�����MCd���F=o�u�6[�s3M�-o����ǹ+T]{L�e��Wr`���Z-t�-�pᰒ@W9`¥i,ԏ�Y��x�,�S*0a���aV׬J��ݓ��ݽ��VH�s�>�ٗHn��eU�lP�c~�`3&}�����y�~r,�E_aP�;e8��g]���KY�v�i��(���"��
r������ӧOmC6���e&��8L5ٗ�{�-�KF�ؑV��9���(�O�
o+�F�હJ;)Ou��~�P_�0\ٚ�x�i*��6RИo�:9qs���^�3�!�����a��PWRl�)#�\b�E�\��i�����&�܆�Rg�`Ҕ�B��BlLѸ��^�&�i+�� y��Wv>\��ߟ=��qw���rc�'�e��K��J�H�ٌ������-����m�/W��5�,\�-j!�5a�F�\��Lcĺ������������rƳ3PƸ��&+D�B�q�DЦ�����U���{����q��77��8p�݈C�Ӯ�%��R�������X�2J�u�0	��.�(±�E��(�^Ն���LǶ;�wrI�vi��+Ȃ�v7Ҥ�<gW������W_}���������:٢m��V�_��|��Xᅨ�����xB����'r`�@���$*Bfʤ���@�"B+l�#�C��H߅�S��ő���[����U��dB�E�w�f������33�Ѕ��HB=7��R��l i\�א��@p�N��ɮ��<ϑ�y�����}���T�vNȢ�0;�U��Q!U";f\j왈,\5g08�EG���kk{O��=|����w:z9E��~�Q�s��U� ������w>��{��s$մ����"�1d�d���?}��ʝ�N���A���g�,�@(���V�I��iLI8�d4ۿ@,H*9 ���`8�Q?}78�~ק~�F��e�P֥W�m+W7��D��g���O0?�md:;W~�QF��*CDΌ���"��?�5�_g����/��r����΋�ͯ��=��ܠp{q�B~j�Mf$l�7ibb�����aZ��*~|L�2�f����BE*�f��p_�װ6�! �OD&B ��Q��cY����A��%̃��'0B,�����"�Վ�:��0�7lqdH04*#�2
�vYTd�̗mmH.��YX��散��vUxI�&`��T�%�4��e���i������v�X٥�P��������Jos�d����Qg���;�*�/�W,uu��<0�Ә�@H�{V"Ll�!� �E~�]�|�8/QimS�"T��Oh�+-d,_]�gjBz5�rb`��٬a��V��&��j߻�875}�qt�9�m����n#�"XB�|\�Mj�� fJa��ԃ�l>H׃b,��P@�7ܑt��Ǧ���H�v��X��Ɉ�����I�3ky�i�dH���6�{D���վ���*�%��~��ʰ�
�B�$<��iD�r~��|%�LyEm��	�� \V�j?���L��'`0z��_��AM��fLV<�H�k�0�,�XJ4�nj�h_0ݝBfr&�٪�-�`�I�w��%����[O����o�Hɖ���6wп�̑�p�\u�aaD��������˗/횅��Ņ�)��3*�pAV��n{1L,?<���rCx?a	r �����Flʤ����� @��@�ʿr(ė+x��*���V ~
���Ua?�%5,W��ڦ~�S�򭬄䗪�Z��p�[EU���
��<����_���C������> ���Y-[��*V��|;-x?}��j��_�[� �	~V��B�I��X��맯$�����p#>!!_~ɋd�'!Ҫ��9�.FA�$��bD����?{����BË��OMx���d@e![&9��_�J�{�u�A�s��ԇ�X!~k�Ձ!�?��?<b�-�8pe���~ʜ��,���t|BC����E��2a`k��	c����)��Cۨ&A�+[����({��i�UM��ժ.V���B4C�� -AJ�p'+�$�8�Y���b�X!Z�" +Nr(�̈́�"���ZC*}mm�R	r��W,xi�/���,�%+3�* Q*���9��$?������{`P�BD͉M�� �Y��)F_��}�U`�짜$�[��p |�(+_0���Ax�
@e�\� �򀯂Z�Q5�^~h@,��_I�R`«?�Q%dX�B8� P��K�R����d^i��mYu������(�Iِ)������ ����VP�WV~�ĖG&�s~>��	�\x��;�CUɗ�V)�E���m"3p`/Ƙ�u%Qc*x�|�a��CۄO��;<��v�7�G#ݞ[�<V���	Ŷ�,�g.ѷ	k�ld��l�?zxr�߹�?��:8]��-s��/_��o`Fc��fgo߿����Y/��UVϷ�y���>u6��裏y��49�Wm���W����Y-//�YȁN����Ш�~V*�T��rJ(�L�'U^9�h�V��X�Je�g�0.��`�B��	�D���5M@���er�<<�B�6D���:�-���ʿq���Io j�B�Pr}2��%Ѥ����44\']`,.6�o��W׏�7�����{��ޫ��a��9sr�酥ə<��+;R/������~�?��_~�Ͽ���:Y���-�VQ�ik�즄{�������/��zw�0�[���WH=!�8���|y`�<��ɿBrp3�#<��&��LH���X}� �k�͎3��эb�Y<���t��7�q�A�W9"ړ�&��斖��Fp������&�g-��_L�L:w�{&���[����g�^~��gW�\�2=6��\��ߛ��k{|o][��TIm�U9� �/�!�{�.���@�Џ�,exc[��'�V{���0S8�YI/��v�,^^��!���v������xj��hw[���&g���tgo�'nEH����Q8uN��uSJ�o_D�QȚ��U3ף�����p���c� 9���9�3�$�,H��U�	?F ;*��l?�a����q�,�Ó흣͝��5�4�z]�Z�#|�뵚���AZt�*�07��?|L�0�a
���AԙpF�_�����K$ ������\Yrhe��Tn������t}�9`�x*9WW"fNH9pR��=��0�$[.�����AQ2�Şc�s�.�i���Xo�[�t��(�S�"+k�ƬT�����ލ4焻��ng����v��|�ً헛�۝n��a�;y���|����IY҄ŕw����B�*lr��l섵�;��6Ƹ�-7��R����&ͤ1ʠ��T!����_�����
v�T��h��S�zÖ#�f���h�b��Fwt��������RsK�� %g�����=�F��h�.n|��E�TgWdK�Ԭ�{����e�����L>����u�ʽ@���WVS~�ki�v�S!V�ʓ��{i�I������B������! ��O(#�59�ߒ�����ʡ�)䇝��8�G�����~F�
O�ʚ#b.w�M"�~�b<���.�r}l+J?�23����\u����������R�YML�\�n�)��m���f��d;���Sc�*SӨ]�cpOPr�<�S�Oz<�١8�sr�������~�������OV����Q��y��[|_u� #���KT��i]6v�َ;�����$$�	i�A��	���G�/�VG � YV��+������)�WG+]9�\���Q4�����>.�38u!�C�zpn���,�U���J�x���oc���T$1��	R.�	��y��k�_�FF�v	��GW�G�(k�mw��|��X=|�x�/y���=z�{<:����K���-aHNt��������<�^�f�Ǣ��!�9���F2�@�U�/0n�^��)�_/��>=�(��ҕ �ܰw�W��&�����5�j�ΫW����.�'�٬s�8�:�y�\}d�^:��LDm7��v~�}�d22MhJ��y���NjN�%���Dt�-��Mz�C��%�N��C[�Ï=2��M�[�g�~B�G��r4BK��0�����-aD�vyTa���
���|9�S4�+
p�}�)��'H?���U�T�vb��E�fTȀL9������-������y�#�L�c��+N����ѹS%���ª.��y`y��S�u��g0Rr�f�LO���崇q����#F���|��;�|�⫯W�X�1ƺ�&h���֭���AbqY�<��o|����d{{��q�u�>�>Z]�������菙��vok�����F�7����'�nۣa,9���HѠ'ۆ��k
ٱ�ŻK�o�uq�q�����o�]�/s��۳|�^d�e�/��ihRc1vFvm�"��Mp"���@�2�қ�a`_l�uƪcq���&KY��F�<U@\;��������#����Y4I�O�,?z��H����M���Q#�^U��M�ͅ��(�x8�6c/����`��H#�9jo$
 �U`m�$���j�    IDAT��:�l�X��H�����E6��煄tL�g�o�8(1��������y&I3t��}��nϼxn���):���(n	�n=�"UƎ �LQ��ڐʖ�<	"S�9t,p�ݒ�_��\9I��[5˪�Q3�'.:�Ύ:��>���ȡQ;�\J6?�o�]�yqcz�u����|����wߛs�޴K�����R���2��]y�������J����7����|���b�'��(���A`%�J���Ƒp�`dL ���[)��H%�b*^��`30��utj��̎����d��ɘ3���Z����ڐ��#���ؽu�d����+ޭk0��u�jw�x����+_?^�>:�V�o���!��Ŕlr�u&a�#��B��lX
��n�$)[�A^s`x+<�3���� �~
�ip��=�sPz�+xp2�����Y��	�W&3MΈ }� G��x�UI���'�y��Pfw�t�_������y�;�@ep䧤�ld`_�{�����l2˾7k��/D�#��K+57��x�=�L@�`�c��a�,�49L�lytp�j������Gkk���'����-���"�8��L'�d��֛�cV8�F��� �2���డ���ߢ���Ox��#Ou���݆h�F!�3b�
ĳ�k�{061�B3�2��J�K��9�*��w{p�z��-��VA��ٷ�p�S��p�tB��s�o4;y�D=��W�sD�����܉i%L;�Int�N�ܖq:�5I�&J�g4�w�H)��[[;v��X�v����CE)	Q0n�f�p�c���I�H+��r�	ʹFA�)-O��9�!�r��vri�&�8I�5��h�q'�������U�E�ﬂ�Ȅ�C�	F�|�P}�ov�=�p��[�
��̖�Kp8ю� V��L���zl�Xx��s��=v�P�hS�M�_?z�vX3|*�x�<#C-�����&?x� �M�:����j�VC�/T�VZ�� %+��7̽�`���9~!V=��0	� �(x����%��q�tt�/Q5d��O��p��I�\����A}�NH��U�(_�˧�$VC�p0��T����5�T���R������O�Vie[9W=�\�!��U����`����2{V?�	T"W`U\A
�X_x6e��"
�^�䄈)�����WZ`\�A���JVr #���[m���Y�����*���*I ^*���`�SN�}�yceE�f|0�(	A�+�)ͳPj�"Ai���n5d�����$�U7	�� ����(gu�(UR���X,kL�j���~�#�AHP������*i������NKj�G�V���TV
���U-��X�	G�R9y*W��*&D� a��j��0��2����ZK�p����O��lH�Yu��S0�U4H�~��
TȰ���MrN*��j���+9�TO�L�B�S��rV����d"!�
DR˕�� ���篂��-!�|UC8l�	l�u ��W>��՜a���n��Z�2�(9�,�"9 ��U�_)U������X0<�+�/'�Xi����$�3�|�
lT*Q����W�B$"M� �JZ�j]A¤�����5 S�7l}�|$^X�F�2+l4*�ax�+���~tu{{[{GvؙQ���l�t�!���q�q�l��|g�l��Ù�e�iveu��̵���"]YH�@ܞ�szaazvaq���Tޘ��F���vW�?���q�ʻ��Kj��]op��
<�A������5aCԐ�� �*����R�B�p r ��x8�FK �S���r+? ���.�5z��i7u�l�'~`��GqT����i`���P����r;�Ҫ���I�.�IW�vO���o?�����յ���O�n<]~���}�.���d?�S�N�/�yg���I[�F=�Ce�z�m�w�}�����~�>��'��zgn:>Q� >c̟�,Q�lk���L�N�}��W��Dk��tY����k�n�2�A�H���I5W�[x��p.��l�"+_�,���/%����Yx��M4v�h�o��G]I�@sx2�yDm��D�qY���ˑ��J/Ǻg����n��������ǫ��l�\��X�]ݠ�]�������{L���P#���Y�@.��IE�������j�]ʉm�8��P��C����~j>HC�W�H�t�!���QFz�^��!:J���i�A�<w������g�,OJ'�����vn�=;�cPw�(��"����٩�����xxҡ�pdv�Ug���{��7c�dn-�^tR��eGny�����������=�_�H�{#�sأ��98��tg�+� ��ab��1�E!D렵$u[��O>��8B6�Oj�iLQL������������! ����M^ С�kʖ���T��y|E����)y�
S�į��qJ��p`@ʾe���zr�5��K^y͵��!
�ϱ�D[�S�!
8ӈ���L�X��.6�IZ��G�����{�?\��o+�܁�<[=oM��ߝ���CM׈���:�h�K�g�ċn( �Ƙ`��J�I�~�s<8�j�YΑ�1jjz�6�G{Y;IZ�#4W���
PWpX�#DT��:�~
/̇��"fP��d�~��Ģ���XΧ%!�@>�\R���ϩrϽ�y>N�:1��L�tx�vp=z�����	�T�f<�<����f6�/\ʬ��rm��z��I��%����ʳg�x̵���A���2\����r�+~��M����j�|�R�Ԯ����,����O���d�[(��CSb6��3��,a���c(ٸ�6`m�r�%I&�&+R
8mCͯ,���͘���>?<�����s���{|��P	!A�1G\��&��QXΨ(@p2�%�Pٷr(���bg�pzr:ڼ�{1�j����V�@�����_>{�͊�\��>.9�}۫}��؉�0�3tr$�M�i)$�5}��.�����^�C�-*M��b��}�+`]3�a��FH]Q�@%�Q�|���rE�_[ߥ�r��8�-mQ�%I�Ģ:F/������#�c�,�wN�nQ�ǚu�G�ѪE;]z��ǖ�/��U{^ �i"����\Fs�H7��\�N��O����;jϾ^^y��y15}��[��c��^���]�GC��C%��u1w�ԄpD^����O���YC�~��z d�W�T>`0���ʣ8�r�V�`[*Q ��J�8�I
���kwQ�z�Y�������	Ξ�p6m���*���Th��j�p�8�M�I���"t�,�z���
�*vԎF_��;�{�����8�RU2y�"��܁E �"����0��i/����9�[�+l@;$B�ʖ��'����r<Σ\���+D+�YTek�0[O�\8��I�24Q;���F[�
�{���L=�"DG�\��X:����K?�5;�2pf���N����{ZH�����?����t;�W[���o?~����˛['��Ż����}�rg���iF3ux�4Ԩ�,׷!2��0m?t��設]����B`!��2���j����p���OHl�B÷3����ͳ�.5�v۔�Zi�O�3�8�����,G��]7��:��g�9[�����5����d�mM,*�
pi2��K	0
����"bf���g��]�b�E����?!y��AZ�9���W^�̕������;�tz/�6��V^�,j��ZZ�˻EBp]�V%"~h��
�\����������&P���R�����}3�12D��ج�)���F��n�i�t~�],K�C]͚#a���&�5ie�\�g����}��{��p�U�'�����OYX����20{N�1��.��g�k��>v~���0��X�� GF�W3�uL?��,2���.��"�13��U���&Oz{[��϶����7O_�����N/޹#[df�����ب%�՝�����೏�w`͹���\FM�>�889y��Ϋ��YTq��6�@~��|c,�<Z��TWVOepKy2LF��8~�<�(+=�K�<\��X�j��I�pӁBLgA�؜Ѵ�1$:[7aݾ�`�A����A�y���H<�ik��>Z!��$��x�S/l�b�����m��}�x��z�x�U��l�s^p����u�Z�$g��4yU-4';ų��m[���`��g�KQ�6ß5"�x(�� ��;"4x4��Yq�^5�}��/�ڑɩY�QaZ����B����-l.�h��ir�R��q+���ʓc�l�NL���2����R��t�0�\�Z���ȩ�zac)�4ʭ�J­i���u�����G	���n�m埛���k�'��ݣ��������/^-ol��-o~�;���A�m;�pξ<-�"G����\7���k�}B��p����C<�dB,��O��p�WH������|͡�ȣ1�E]��g`�����D{��w��j�Yev�1qл��=��?�׈��3 �H��B,�-+GJP��-�J��p�("���}�^�<uL&�;�t&v��=������7��;�?�D|�$�����=g��J�����Hƃ%m�3�H�As"va��Y�$���9�4��g�}9!��G
��R$��YH��k�9	� �����`)뚜�&
&�mh�&!��6O�.݌͡�o��J�`짌G�9���̜�>�k:�5�@Vv vRD�ssUTIcӶ����fl���!�щ0�<Ӄ��>!,-+���Ҿ���swwύ<%��6ۄ(�Ac�	<N8� F�DA_�1�J8t�%���F���e(�`��`T�&+��_y��T��w�����%R���$>���*�`|9!5�T�R��}�P,W�r���S %W�@�y�PQ<rR bS�oј�-�O}�[9���*炔�_��+�*����	��l+���*�2R��SU[.`i9��G��__���
�U%r��p�r�b��Dw	QGl󭲆��䀹��}�c<z􈒤��i#7D/��Q�5��"Ʌ���r������$b�w(��R}d΄����� ZIY�aV+++���B��
�\�1�JW����M ��] ��(Z�J�ji-v��' +4��W3b�[�T�o0X��������¬¤� ��RxQ ��+��P4���#r.�ʰ��@ %��7��r?��w�}������P��Y�}���2�����[�	��@ p�'?@Y�_!2��U�Tr_E�Al�%�ky��]Q2���\�2��D�A��0/�A�������)0��(-3x�[P�<e�t�J[�����  @߿���#7�(�*�R��Uq����@��au.0?�_0r��U)�O0B���J���g��('�*�z� d�U��)��5L/�|���HBq�B�(��շТH[Q9�h���ht[<�޽�w�j0�T��e~~qrx���<���Ý�iW�~s�p�݈X�7T���k���`J��."q]3�M�[䒥���O�Zp^[s�BKU[5
��ʣ�«��/[����_|��,�a�+�.H��V�U��
��SrI������e�cL)��
���8 ��g�k�S���&�J�:KZ8�d	���4�O��P��JZ��V�]6R�
�KY�h�<�a��$$Tb�;�w����Z��Y�d�Jn��%H��vb����>���������B+��B�1�Q�a�,��U�ld����t���UWQ�:+�Z]IT<���t�F0� +L�{�
�d%�SX*����W&�2�! �_Y�z�e����c\W�{�}��'K̕����Y�p��y��أ	g��Էl�(���X����s|�)/�b3�5SKw�ϳ���
kYpyf\8��\�',�CP�����h���עI������S�j��k��~rj΁Q��Z��Bl��q!�8�.�ƊB������������gw�x�̬g}�R+���$���u5��}w�������N���z6����l��t&�I�Yn�í�}��[k�4dPO�N"x�������8���O���6�+�g&����q�#�4o���9���ic�hN�~�J�&����d��9S����o���}9C#�XYYq��
E�%�& u�]UnJ�R���*UV5��@B_�@��pE�Pl���?�����z�:�{�w:}��΁A$�a�H����k�ۀ_�����q��x�F#R�&�l�s:�����7�.Q�k�Z�V�]����ׇ�Q�Խ~BI�GD ����nO��\et0�;��{{�i}:�MB���V����]����ѣ���sK��j����2���)_���J��v��v4���`G�Mfh@��D�r]�L��!ӅʵOrJd�8��O�%����u�%��T���G�$тXU��ꔲ�Fu��:G%������-.�˓�)6j������5�����ɓ��ť�n||�L���~}��Ղc�v�㣃�vTȈ�w|j>�V}��j	��&A25��"�(h5���O�){Z%�B`����sF���C��q,⏎����WF0��	oTp#�H '1d�����Ɨ�t���~�f{�!8ƭJLb\�bj�����.�f�)G�=��'$P����۷�?~���A�,g��p�1��~跙�+��#�X���>9���w�:Wu��������~ޟ~��ׯ��L���&L�9�bnљ *���G;#�H庝��*+·�s8J�!$�K�vދ"S�Q1�9���]�1q������뮪 fd�t	Q�Wo���.9lS�h����&!>���#�D.�w~�z�+�g���<W�=/=3:�?�MW;q]5Ds����ۥ9DS�g��܋pv�H�x�����<{��kǅ����[s{f��Nγ��4=���m��٬ܵY42�f]�r�mY�A��xt�`d��%.Em�# � ��� �=>��(&�	�1�G]
2�Fzbfi�����{1i�+��8��
_�6����Ç�u��Eq���3���Z�ЛۃR����V�2�i�Q��uڬ6��"��9����މ* ����#oȣ��&bx 	z'u�o�$;� ��Q���E�Q ��XR\!���s1LG�T�)Ɠ���
za�l1��b�$��l������o�b�5�n�bS'��73QǶ}�p�J�E�i�x��8��5/Y��*� n7+Y��j���+��Ӏf{�#g4/N�w϶^�x�zskǸ��r�so�-���a���l�W��k����<��i'C/mN��wN�7 ��\�{i:��1H6��X�Q��x/�wጙ&v��������՛:^���8߷���Lb�/�Z�*��L��8���?4�▟��v�6�������?{�5S�>	y�}�v�?�����X����h��D��E�ԗ��K�u=�C�����p��V��ā�"�e��S��Ɏp�Z�Q��3#�©�m�����ͻ7ﶕ����
S�iq�>p�8A[{��f7�	<�pib>�+A7n�����}�.��\�u eD��nV�z���>�\��4����k���z߯�]�Y�ː|[{Q����&�|�t���z3.L�X4�[��q�{io�5�PM\8�������/���?X��:���������|�t�]�������/Z��:�\}i�%٠c!�����D�2Xys��@5��Y
��'��=�c_��pyvy}tp���o^�s�m�Q��Їb�����:>W'���m~M���Ώ��?���Oz��-�թe�f��9�E��]��.W+�WL
4�V�$���R�s�C!���@�,h����<
��J�f�2��^�|�o1�h2=}w8W�.Ef�nAU�]UT�?�v�]ZV�l����v=�|j��~�+�'F�*�!��KĴ�����m�T%�K��[��}����Gd�n��<^�-,�tصV��܎��S/>K�FO��ZAu[������    IDAT.j��`�&_q�T>G9I�zo��j���׾�P-�WNk��(b�g�Z���&l�!:��_5�^"��� ���jt�u|p���[k�+�^v����h�ǒ��]��}\���w�x�-_'\�	j|�,�:��a}�֗��.&.|�Z���Z�PU������������+�����;�~����o�OG��i�؅�j�2�J�u��Ö�j4m�U���9\���x[�:y�~�|[yoޔF�мW��� ^Ł�H�i'>�-�Z�me��M��Ol6����������|�_��;��ꇉ����۫n'\��֋���x�P}}\]��\������Zɷa��3[r쎰7���OH�*��� ���XZ��׻R�Ԟ����6(�2�#̌���ǧ!�'��2�Po�VANy5>D���u̽5D�����\��K�f�FO>	���!��jʅ��p���۩��|(SFR�$o�`Kr��T(3~�_��������8�Сa�70��C�n*�29���i�����N�pk��_�U���i�z'��ʩk���jK�m�\�8��z�I�Ӟ�U���m�!�K���L�48��m�)d Vq�yL�d���8�EƦ�f�9���V��x�����!��l��$  ���b�J�d�"$�$�$5�$��c��x����$�B��F����1\�Z��S��K�A���&�(x�x #���M	Ffr$	i�x�2�������L�8�р����
�	��hK8Ǌ����%	C i�i�I&2�%�>���ĒĈ%�Kڔ���O�����w�}�� ʰ�0i�Wc�*yt��2-4Y� V�'� �7��J"�L�$�="#S�@�ܢQ0غ^n�՛�<�f]����ϟ?G@��eb.5�6�(�=�� ˤ1�2HR��d ����>B����rف]�J���x�zqb���bn�I~���O��#
�Xx���X�����F������]j !\INl�D�����/��:�Ј#!�yD�����I�AF8LdXh	N 1�G,�/ɟ�EC#� �`�
� �$@�4�e i�IE�A�b	�4" �T!�X�Eor$)����T��3����d1<ɐ��>��=$ ��H�++D��!�A~<|�Q(cu�D�#c,Cr$3�����`�H��Q�G�Z�0Z���N��Qm������v6jw����S�a����ή6���L[a����@FLB��W��J�';8�)�Ld�ܿm$#�=J���9-�!��d!@2��#��\�������Z7�LI3Ufe<1!��Vo��G�<���w�	d�p�F�r:��'O��Ð�b���*��hQS��6� �
r�B��\�*��$����'�h�xYb� ��t��:����@�UZ�.���ʝ���f^l��߯����������V6n��a�k�B�!���pV�1�t�R�o�qk�>�g�:��F�S�18�'*�T*#�D 0?��#8�IM�O��#9B���4� �^��.5�#$��S�(�C1?�KLD	j�K�o��߻�|z�޻Ӽ��;^�b\)�ˁ녫�������	�n'W��[b�B��␑�ޮ�j:���/���\�֊SWXjwLl1�l�-8��eJQh5q�G@wsH��[��z�?�1p\�jxX�i4��cl��[�����צ ����X��/,SD�Il��wkyb��ey�j����7����ف�)���F���'���]d2ױ�ttd���Ω�1ի����;��8�b��rYYY�,�n�G[�!{�:�W��4m=O���g�
@��d wR��@����q[I?�]����1��[���dt����k����f2�X8�(�0B���PF��	�F�F Y��#��XFC)�U0���442-�ҽp���K�7�g��9s���~O����3W�����Z�
�6�V
�is�m�.��~�n����٥�3�ӳ��I�������bOU�Zwˈµi��t[\L먛�>&�ݨ.�g��q(3!�`�Ԭ�R�^ٻ�f�e\'�X�W@����"M�\�]X����ק0�'!�rKE�V�� #���5��jF�U�6qc��t�������M��\�~��g�[XjU�K�u-���䥭�N*�_��)�@�,U��d�P�W��b��S���be!��L��Ne�sX�@ / �: w��X{�A�>���.@��T`A#�o�2q�Y~CC�Q�H�.jvn�z������f��ܜ�^/8��6>�-��ht�dR�49&ۄ맸�P�zU=�#�Ui?	xI���Pʗ�B�?TTy�Ÿk���Z���q�3��'�{�t�#����-_�����Vd��[�?��|d�M����;'%���C�X�Uv^��!��-l&��x;%_�cA#��#2q #GK��=vbH�b՛m*;1��:1Lb�^D�;R߾���׿Z�_�-�Ǐ���`�ۖ��ً�z#M;�fW�E݈�>��XJ�����瀏������;���<�;v���{�ު�S���*v}��O��=��Va��x�ʅ�*e!����Z�*S
]N���g��T=��>0��dAr*k �09d�`���v�C eR�$n8G;$� �"�H��X�@*�	�FO����ֻ_��kU�ރ����-��X���9>��;s��ʮ�&�
N����>m�w����m��ؗᎼ:�
V�[R'i$��Ɩ,�3t��'0��q2��~��Rv��*0.&%N~�XH��K���,.�R�pyd8ĺGZt��d�|�B�2�2� ����P�� :�6*�j{[Aԗ��u۳�o��X�T8Vg�#9��d��|��[��1�s���̟�Ƈ�[o߿5�q���sp�cd�������Z�s �/&+Ǿz�����"�My/eX[3�nCi�49�(>�t�+I	���w>/L �ʛ����Nɋ��[���Ѳ;]�)��wW�%5w�^\<�?�EC�Y>��<x�rt8x�����݋}紆��SS.!�]������uduo���>?߹��KЋޡu&�ҁ=;d��zC�W3u�Nh���e�e�~Y�F��{N�g�u����k?���z�f���kCt�qZe�4���
W������d����{0	\�X �p�덬�D��$�Z^��)�Vsn޹a$���`������E�I���I��n]}��ϬΌ�nߞy�>�}9�2�W�Dm谌�e������89�^|�h�p{�����٭��Ȳ�������`4s5:�ݵ�`�����ks/�����>��vv�u��������O����=�u����Î�:\k[Z�Z�J���ӊ���x���*��'>����7_lo��P?<�@�-�qh=�(�k��U?�i�9���������/��JΙ��V����=Ɨ���l����T���ZBk��X�N�  ��ZQֶ$�B���O8�Ѓat!фXS�=�_��=2R,D�p�����������woo����օ��y_:�Q�r��w�./D� �j:�*݆���v�O�D��L�[��p�+*0�n����b�~������{�q=��ӑ���[˳�3�6���H�@��\-�R�W��_o�I�Gm��o�؍�V#de��T�xC,�2�p_��������c�x1����V��.	t����Z�<>�4�a!pa��=9�G��i�v����VjVc`u�$[�|�]���~�w����X_�[��F>S�i#Ij,9svQ�Uǡϵ��Ƨ3��wL�V�63�S���W?�*&
�%�$�Ob<sz~}������l��ѫ�^l�r�[���~c�o�����i�u�j�1�ۄ`�PTڄ�i��/h����S*��y���k�S褹q�,C
�X�ֱ{5��oƥ��f^�5~y�=*����LԸ�&�C�.7ZK^X^������G�� O]�LX0�m^��P-��x���U�F#�����0@V�3�*���ZxUOo�kXn��}B����f���{/{A��2n<������C�ȘNRߎ�V,�-����0F"cS`�#VeY+G1bq��X��֌�����!F�R@�^l�\��OOon:��~}��W_~a9ë���'�g��Ѱ;#�t��xj�6U�JE��	�ѵe�Wi�V�Sd��Mqʳ�u�"q�Zm��c� ��C�ʅ, �A���E
�u&��T�ȉRE���ˏ�-�!9;���R� ��z�%H�`q�J��qN�i���@��y(;���:�|j�,{��q6pZ��i�
&=�"��/N� M���O��Lub�Q��c�G�
�X�	�����a d� 0����L�d�� R	�+�?�9����U9�čjH��dv�dPHe` 4j�	.U/b�����!��1�ȇ$�^ -F�~��yL����|�#�YT���K���EN)��`W��m��$��1\�E2�~h���7xǪG�yDIk��[]�@\̒I0�T�Ȳ�#c?���eX�����j]�ǿ,Ò�a�Tx�'9ĭ� ��Y��,��G(	t���T1�������zH���gϞa7yJ�_Yx� �a9������#��R=��R�jA� Uvd=F�B�>�����,�H@^��#$b�x��$SQ؀L�2pT��G�(�4qX���1�G�"�9+��Pb6��G  %E{��ş �<J�w�bË2,��1�?c$�w�B���18N�R��_,&�R������������G�=��7\`�$�i��XB㨈�mK&��c2��o5І��O�hr�HUu��j�6!=wz�����_��Wci�س;�� ������h]W���޻6v�Z$��.>T��[����Eh���XNJp��9D'�-������oGK�Qj�)k �%
^ �G2�!�+R��B�121cBO'cDPyl��X%z��"�b4�	T�$��;3U���yz'2c2�r�>����5�{��em�������3oP?���T_W�θԕYZ�ѣ�m*�s������ںO%Ԯ??K�~]�=urWY0��j����|s���_c������U!����*N�:d� #���c2���x�°!�0t�1���Ǵ�Ў�\���(�4d��x�򯓲(��U�W������塏|�/]�R��ȝK�n�P����ի8��_�p�hR�������̘q~5I+Aֈ��ȊTm3%�lO��s��-��R�f�N�~�$���m0!&�U�#�̖�$�9'�Lv��1F��xLH.�j͌�����f�.̰j�ǫ�H�_���O���h�$-k��O��¬��ƃ�̼R�߫�����ɫ�)7R]N����zq��v�U���j#������Ti˺6��ⴐ��0��T?Z���+|vl�&��*��&2+`�x���9���W_yɪ�q{H�(]cԁX�����/og�^�� �AL]�97[1!AH����z{0���B9z V��ńH�Tf�e!�4bM��TU�4qP2�D�P�C��B�H�L��<<�^Eu��p�c����̌G5G�&������W5�x==�³�RZ�Τ��Wg5ک�)Ӛ:P���I�u*�hܪ�F��W6�H���Y���ou_Z�q�h��$���R�W�x�`�y���� ^KD@L��4q�����=�(fF������s܌��E���9�v���y���/^���7k�i\����S.,�.�Y�d_'����fLʰTi*R�l+2����PH�*�0�f|E���o�,��`IL�Z	c�w)��F���8���H�2"�������9q��&�3&6��p�x�U������^|�1X�*J�i���mR�&?E��-��K�k�Y���=�۞��ut��4��\}猹c�Õ�\�I�Р�ds����j�gb'3�S&1�"!uI��Q�ᵞW9��vx��/��� Ib&�u�I�ǽ�� � H�`�b���®p��	� ����5A��]��aː���9���ZYY_���y���>1��V5t�4Q[]�>֓c�'N��r1�������u��ZJM���Z�}�?�;qaނ����t������##��E^�MV�M��,�^.?��
R��bI��54|(��#�IJ��� �B|	&��梌{y/Eb�,%	Ȱ��U0����ȗ �Q�mm��z�:��UUza�g����Z�|7M�1 ��7�l�����v���[ŖY��RmK"����b'`�8��,����ŘԜ��������$��A��#&<r��B��q�!��Db KH�D@	 ����ֲ4m����~�X�N#Q̓� ����ߛJ0�adiɸϒ��������|`'�IE%p�¤x���uj�mgW5��ȫ��������w'ǻ#����?<w�����`��^Z��&O�ӫ����s��|������ű�t݊eE�Κ*ei]��v~ɅR�/H9:πe0��;4 ,5^�D`{��u�����l�j��7''wvލ�o�߾;�4xr����������qO�0�jh�u�5��������/���O�����L��N��4�V�>�����yx���_���j-�fn�rs�)���L�����1e�
����g�]�磳n�Sÿ��޸��mYy��������:����z�Iɗz�M�΋*?�Z��!R�,�n7 k\��S!�0��·���=/_��$����y�A\.��(��e[zk�Y�`E{���ts�?]�^�;�u����}���n�����9Sٖ\�X箩�]6�n}>��ۻ�������Ѝ��W*�Eo��:�W'G�Ϟ����݇�=}��o�{�Z}�@��i�VK|���D�XAW�گ�ꈬB�*S>W�~����U����X\��{��2{ǚ�֫�o6_��:�d�m4�nӾ��î���׵����ASek�O���<�����ӱ�1ά@��L���W[?~��9�2���Zӷ�� ��%�������r���꒐�^���;FY葐�K� 0ʔBR��{4��	��x�j���۷�޹����[Z�U�q�ib+n�{W#�����b��5 �pj"�Iڰ7����h�ٳ�����Y/A�>uG����dO��j[opw�`}e��Q���2���Y�l�%��}^.u,"�L�MASUu���]��!ɚG���2| ��m���hH�� n�5X�Xڭ�R�ɴ��d<;7�1���	7�S���P27���j:z��[5 �.C�Ã�ý�7�^>x�������������̠7��/�/{$�A7UZ��]���MͲ�H���j�O�ԝC|��.��������mޗ���?�������7����v�%7n�u��~����\���qM��3���T�)!uO��u��oq`:>I F&�H~s���0!��)�a���o���q�xY�4�`^��$K���_is���)���{��n�+fqa��Ν�7��N��|!urђ�C��^�u�~p�_��o�\����7�Z_X�-��g.J� w�9�����6�+XЁFˆ(Fqj���-X�	s#d�L|���<"���O�8���i���� �2�9�%
=< %��,N��h<*2�$=��<3` Ni��vwv�?.�>�Ŭ.�q?C��P�9����s=B3����j�Pw�1�
�t.~W�@�I� .���>��IƳ���y�)��d!u�<ʎXHv�D	l#Gy�`,�"�]aыLjxq��^.�<@ ���I�0A�H�	`�Q����BT�d$(FC��c`\�cؑ%U��ť%�<�0�PR�`!IdF5#&I0Ab�8��Ab��8xB�⿙,$�2I�$�`��ML�^j0.��Mpك�bH��RY�&�!=F  B�0Zz�=F,d͊���h[pZy�~Z=3H�R�v�希-)MMP��.&�=����ߧ��X��#Ы��&V��6��BC���:�N�x���i;Fd�s�    IDAT,$PG;�&����؏L����9{����od
e��E5E��{&?~L5�)�F������O�Z�1H��I7�嗸�T�� �
�.=Jvӊ8.f-��Y���Ѵ�6s�%�ƾtU�X��칌(ޤ�aD)I��O�<�g�a�������>���g%�Gn���3�G�:yaF���6� C#ɱY� 200�G �H ^���
HZ��HyA{�?��|K&���h��c!�ȏ��xHpt��Y��1 �
ɂG\��N G��Ғ�	`�$H�	 �1ZXȆ$�%1,���B�OJ��̠��IL�=�Р'б��ϓY1Lʈ�H\)�Ћ!�+G�.�ɏuu�ѣG��g��0�z1^03�T0Lj�:�*�ު���Q�z�~�vKB�C�"�e������ 1p%�)�㽦��.yQ�5���f�g'S5m��S�1֊�]5�Ui�?��O-EPJ.Ĵ  ��d|��8�ї����������#x'ߣ,�ٟ��^�%W�=	�#�\�j���«ٯ���+�鯰��/ȁ��f��`��A'�����3S�����3��o�w�
1�x���O�~v�����K�4iuO��D#��w�ռ��63�_��_��WR��x�!=-Cϟ�ٲ,n��u�Z2X�8!I���L]�r���@.���TH}fz���h�#�G09d"L�yԩH�j�^\]����Q}`�J7��DZ�}�������;[-�A���Zu��_;�5o�җi+w���:�J��ژ^��R]Q�lC #�+���Uu�-�p	d�xz�`9h$)#1!���2���9��Ӹs׻�ޏ�co(��I���+��]�2�tU�)��G~˞�Μ�{��h�������h��������K_�5-跲�0���DK/Q~��J���8�f���t�����Zse*��l��SNٟ�z8-�ӈ�~���/�0������x$�{ԙ���{�s�TI�q��Hc'>�%R,�ءOjj/<v4��`�x�Jʴn+���dM
�̈�A��ȑ�-��24Qf  R�Z��ӭ�p��k�hIV(lux�O�i��L��jx�`��jjtv�(���h�sK��z��t�H���y]<�㑖�̤�zK��^�r!w��`���^�۠V� �	F�H����N����-x��i��C�ې|�Xj�5��G�Tdb�'X�m�U'P���[��m >cUw빉��]�KXW<m��ݾ%�-zN�L�$���δ/Hd�!��<0^�$�*�ؙ���7�(a��a���.������ `�p���H{\	�Y��F9M��u��GM�jo(bC/&G�a"�=��(�ӓ#4bIh�4�+�C�0���id	2\bAը~��4z��ҫ���=4��f ��JP���3$$#�h���J"P����6���!hZnz�`H�1xd�	�� ��FRv]u����h�����'F����L&LlFPoX��5����N�V�)A?a�z�a�ؼ4��(C��[ʰY�ݟ�e�'���~����_լ-���U+��ź����ZW��4�D�֎��uf�<bO��6d$��+��u\RU19^��TH�x	��Gd;�#]�؏�o��/E#	��?���F��1K	ͥf�ka�.Q���@mD�Ð����*����X\d�лb7����Kȶ(J�0"��ɗ���T�t%w�I8����*@�8�M,�+ؐ����#�,���0 �c�$\0B�C#/�!VF�N@b@��G���4x�$�ۢ�	�6Wk���s����i���Ѯ(9u߀��* �u<���>����oN>����$�>��~W��.{��K��[�?�{��FtV71�O���|�� HNm��J9j�X�fjx�
����l\�0�8���!1�A0`@�j��Ǝ� ˵+f�K����'�o��/�����{�-̮�ս�\�&X�P��ͫQ��/��G;o������_�~���d��A��H�����q��:J{<sq��ը���;���E������py�yq_t�,���.F)��ߓ.��ݞ��ݩ�O��vv}��ǆ|Z���R�@ָ�{�K�`R�"���aM�8�8u)C�^� ��Ɓ�����z$V@ �E'{�ኦ��T]�U)V�ǜ~]���>eеp1��_����ғ�?����=Z�������x8�Ǻ�Bwj��R�%��󝫃�g;o����继�m����4f�-�8|f���<<=��/��W�W�|xnuc�Y�A�񧹁�q�W�jk�M���@ߨ�������V~����!�n�����{���-^�;Z���:\X���_���g"�b���̫꭯	6K���o�x��~�6k�NpUV�#-�o)�S��啉��x��_�ҏ�8���<V�x�#d��C��<�Z�Ǯ ���[)T�R�A�-&F����c�H�}�9�ض�TT!�����,�n2X�=��4t6�vA����umJԂ��QՅ���?�/�N��*�-�}w������λͭ�7oOl�:9�Rf�5�	�.�}h�2{�{|�������Y}h�Bo����i��\ǫ2��*/RZ}N,�R�Lq�X��=���[�鑸_�
$���6���On{�i��.�Ԛ��,YF��o
�ZϦb�|Փz'ֶ?C���[+�ˋ��V�1]^pQ�EU��Q��Y�Q���?r�s�ڧ�l���!��*@Ǣ�P�q�#��S>�n�����z��<�/gr�Loa~Etӻ��3�'���������&bx=�L��Z�p�8�=!H�8<�*�Í�9Y`n �J*!`��9!)@�3,U��F5��L��ʹ�d��V��&���
��]����أ�C��f5쥥u�����>\����Ywx����+���S�X�.qo�I[�U=?,H��z|c����U�'ƾ7j� �x��E�RqU��ƢM��o޴��� '�l؉��p8wat��!YKǒ 	/!]�'�p���
 q�ZE ��&H�ғ�G|�ӕ;��(֢	�7�9�|���������BZ+b`��
ꚜj�.����R�ZM��; ����D�b���f��p���e��b*�X(�H�l��	I�T@.�G	��b�R@��+U�JFx�Q!@��XI� ���vHI<IT�I#$���Ⱥ�H�!FF�����@�z	��1$9�|������{��'�{`��\,��j,���cQ=�Ë1��:���(J���>6�`Ixŝ�	�82�&0@�Ԇ�^��Θ�K�!��۔F��IQj�:)�Z,��IFflFb�$~ �]���6ۊ�D}�K�a n$$����D�D���L4�����Pfc4����!�����T,/�(��@��H��o���ӧd��������������ki!Mc���*��TY�l���
�R�y�����ϭsXw�C�%L���5�1�)~vc���''ɪ����&�Lɯh��b�^�ҥ2(�$P�{�'S�F_�3��_�xA<#�
V1�I5S�(id*KhdJ�%�b�b����4��9�ŴЈR�X@)HorJ�GNT�%E����DI d��C��hG��.Hq��(5vJ�"6#;���c���l�daG)&Vi`�8��N��@��hG�G6��ȗ<�4c�E��aT ^1b\�GB�a��r<J���$����<ihRp<21bI�ӊ$i�۲8�$��"_j'6��Q��R�9Z��:��/_Zऋv��n}��q`�@��c�À[�N��C&Z�r�A���xU�(]��.�������gz�%@~�EHJ*?hS�;z�2�UN�)�X��~NF����^�lF��XĄ� �*�����t�]�X�f ��G) �v�H�S�3�>!0ztZ2�a������L�b�J��~�x��Ƚ��>7Iá�|��/�<y�c*kl���mѭ!�j�^
�f3��3�p��.�-L�7l�Ğ�eeiv�3�MA�	���6Q9v\$�	H���2�5�	�X�G@`dz�d��H,!��!)�А-_0L��EM��#�f�V��j����vD���n���v�֔�{�����7��0�@߈_7g�֭N�"M
����J�
���^����얩;���/�6�I�W1���i;x�#-��͛�S�L4R�JQj�`b�ݢOU<:tA}�l���]������_��-�;���f�Õ�����g�Gk�^�~����&��M����w�
�����C�{w���ppsۉ*ӟ�u�"GecM�p�߯��3����75_�ш`�q�y��ɟ����W��.����'�븜���w�Y��1�<�0��(�Jm����F�^��%5����'~�0!����2���>�$�##b��n�;μ��Ͷ�}�>�m{��P��ZMu 6�����3�fۦ&חS�S���ﴗ�a�6w��i�E"��y��]��f�أ	�z��(�i,)��T)7�Sd�<ّ��2Eu</`��<!�1�7\� �X���H�R�D&C�d��fNġ��鲶�?ݪ��9�0�hX�?-���u�n�cмܿ\����;զ��j�k��$R�f���`&1CUT<R�&&�6~�0�,G�NA���X^$��#idrTR=�I��%�Pl�f��y�Y^�=�/�Ȃ�CFJ�1�O o�0��$vJqK"J+F$�C�U΁>cu�D.b9M��">Z��v�r�
oB�T\�r�ap�!C���<�����i.Iɒ�c�^4�$#����q@�Ɛ��TQ��f 	��!I��@����#6I�O����7��i��]�֟s
b�%�q�T�eޏ\W>2�G��X����y�k������?���l��s:�q�ȡG&�&]��W�>c�䠣���:(v!`�r�Z����38�8��B��B,��$_�y�Cibc�H@�N��F�eMRU3��v�U�?6@#J�%r�C*�B�rb��3�$��#I�6�7�����SuI��@f��W�=���}m�B����:�/�)���"�o�E�Q4W#����J���n�=^�BbdU�HƄ&U���G.1�1L��fg��d4�W��F�����c�+#���?u���>x�H�E X�Jr�S�5����E���I}�^��Fѫ�O#�-.ܹ����:�[ �-�<�3��Q�����+��Y�/��F`Q�{Q�����8����Q��R�r!#�\�L�����L-�c� {hB ���9�W��>9��ƙ���s�JO�ͺb�G_<4J���G�g,X:�J���SV.%��]z��z��7׿}��w��;�n"�_N����^�����i@��!O^�9ۻ�����Xv�ܬ�j�k�˾x�/m��Y�� .@ѿ����:�\f;~l�`��W��¢�0j��4G�^���2�&LX0����#�z���>$�C�C�[㺢�ٳg��o�&�F�GP�k���E�ۤvB�_-����
L�A:/�����|�brol����S�˃��;�&�����0a��]�q�O�V�7�3���χk�
h���w��>�z�o����*��6�#w3'3��g�ۯ��o����5aumqaq�~u)��١����\�S��g��Y7�^���h��k�;G�)����q�vU�n:�Mί.[
�����B�:���ڣh{��Q���9���ί߽������,�9d���[K#T�Q^+*^��Wz�W�/~��o|��:~Vd܋�{����ԥ�� ��0I�.-�8�#I���q�����G�TpʴS��P��t�*��$u���Y�7o6w���ϑ����:��8��^�ٟ�9����b��[zno�:}lFq��ד��{;G;��{;�ۮw���������~�Ϛ^��s�v�م0qٟ8�q���p�z�:�[p�\��V�9W�l��un�g��rqE������9�-�t 7Ɓ�B���Q�KŐ����Hn���{N� }�ź��ɥE���\�`T\_
4i�V�Rv�S%*��~e�K��to���h`�°�O0�/~��_�s������:�N��������!�[���y+AG�>�25v3��c��s�~�޹Zcg���o�$n��(�k���rvP�v�^�U�vصݢ��������Ud`�$N���@� ��R��ę �cI�qH!���n�~%5\]j'����l�t�ބ�*�B�NL����y#�:�}=;^M�}/��t��x�ݶ�m'�+�>[�3�2,��բK]l�R�.�ϼ�S� V�GU3����#WI�2Fn��s�x;��_�D񃱊v�6���]��ɚF-��K�L9�`Đ��QW�1J�丑= ����C��.��$A&/�$fӛ$1�1#��Ulpk��~����� ϼ����{���ޥ�����ABơ��u����l-��]�~[�|�ym1�S�����PH�Sh��$�"C)1<�<z_t�
 �TI%����Mr����+12����X�*���n%ÄH��$@g�$E	/� �B�D�� �v�'4��^Pj���R�"����0 d !��(	,	qR���\GB`2I`z3 1�GBB�ωB��#�A�FH*�d �� �ў��'�0�Ј`H1uXN��Q�%(a�aIB�~`H�I&��K�$%��d�^ o�	i:3{D�yZKo�m�g؀E@�Э&(_��Jn�ø�HM�Z�fƥud���h�m`�K$`DC/ 5��V.�D/���Ȉ�L�1��c��͗/_�,aQ�h�}����9���?�S9��h"�(&���ϟ?�+6=}�4�rk�?�������� 8Hf���'?����k�JߣG���~]G'A�^�S$q�5b�)B1-!�Xz�$��P��p�w���B~�}���!)<1�b���:0 �R��d� u�^�=ʹ�-f��#��`��
�@*�B���R��bpx� �.�1�F2�6,�	�r	{�(�>��F�$�N�#9Q��(��0=	�f���b#��P"ƅ7x0@�"IH�]2B��L�;�xᑡ�"w�����K��E$ V��&�+[��Q�&�:dxIH�͑�X٭c�4�TZ�G�(�>�a�`������YK\sZ�S�(UZ#K�&]#=*n�@���RB��Z~=
lC;�/b������\Iɪ�B�0vrp	�(���@@f�$��"I��02@�T���>�D�{tu�9��g�bR$S]��L�_�Lj�p8o��#_z�b$��!��0�ƣ�/�]՛uey�aO�������E-.(�:f��cs'\f�Ss��d�"����ӟ�tss�ШN����R"X�f`k%!������d� ����������+m0�< �8R!�=�����;y�%$K����gk9����9����@��e+�_<�dy���y�Қ��\���$�����E5�b��"��I'-��	���ϋc*i�)e>"�b��P
I8F�H� �I�,�$˝RP{-�.�d]�؍mZ��%U.�W�ؓ˱��yM�X���/���J���r�����}������wv�G�S����9��|���c�G4'�n���TBj���W�A5ۼ����u�:���k�(�q@�������������Mfi;�&���U��9�0;��dn�(�`��XR���B!
#)}zT*�˚;z��i�"@v9�1���C�>��A�F����(�fj���������1�v������8�_�%���t���a�̪�8�>�����R�/��N���Xt�8*���I��������T���S�Q�T�FF�T@�]���K2�+���$t�2���0$u\��I�W�7�k�e�o�f�9�����-���f��T	z�W3U,/%�h�h�/.���7ɵ�/�J^Є@/�#Vd�����f�T�B�E�$5�aC
h`(�|��J�Lȑ�%2* ��U��*=X���F��a������"Hë���-��+���F pv��    IDAT�Bd�����kg��r_b��Z���`�b��W|�Ji��F/.��8�a��2	��^���S�%S`���8��?�B$ӈ#c ����J
�&	����$��`�L ARDa\�Z�6$8��3�@�mA�T���>G]UX5ǥ·Q����-����`�_�b����D�a�����c�;�[���z�!n�p0 �xC�r���6�2Wn$}X �9	��	>�RqE�����gd�3�G�(!r��=pl�`�C ��FQs�ME2�CLʄ���&@ �^Q�>�G�2rPB�Tp�Kb�l�J%"@zL ��
2�"�W������UD��#J����%���
��4
!���?(���K,xċ>ڃ	)�<ƽ4��ZOu��J�N�Qwr�B�5��1��;>$�DT��N?�)IdC�QY]\�X�.N�S��C���q+�I�X���[@�Nڵu������#�A��EQί����C��W^<���xZ��iރ���G�^�qZ��c�b,~���wJi��ç���G�?���ݥ�۾�7S�Hp�C�SK`��w��)���������o�_={��n�t�߮.-��w,���c�fЫSS8���Nm��d��m��V5�v��VMk}�J�H���U-g�+�ͨYT�Z%�I�*��"uX�B�ڼn��������<b<#�'.1X��ƴ-�������k��K�q���� a$^��х���-�X9107m���Io�.�]��>|r�˯�=���k�g�{��S�5��A�Mf�xg��z���O�����;߿�����}���N��uBˇ3܋r3_D@*������ޢF2;�sH����P�4�F���9 wzb�L^t�
�
�I3ӵ����ܠ
����{����7�:?\�l����6�ݻ}������sk���c�=�tc4�jU�J�۷���/m%T�\�r�6��ə�+I k qr0���(��)���FA�U6-dą��d�L�Aթ�(�IF���IrתC�{+}5��+��f�直���L�z����f����Pl�O}:�?�	I�&��`aѴe���v�+�:�{�z�6kk�WC^��!_�!���/yo ��r��7�%�5�)f{A�S"��"gb\�6����a(�118>&΄	���M�ڻx��s{ԁ�Kb1Fĝ�G~��"�X����}�M��W��}5`yumimEe���j��ÚdZ%	N�z=��%z+���X����=��%3���	Iߕ�����{�U4V5ZګϒYCnW�6���k]~�l����Hv�#>�o���z���<���|�}$�����!(%u~KN��D~�tF�Y�ڤ>��C����5���2W�U����.��y�`�r��??\.f���ƆWE�N����3�_	l�y@�J'?�G���Ξ)z-W��jNP�d�U3eSF � �b��Hj������ñU����h�.@XPj�� '���c/M� �3>BPb�L�  	��lH���	���	A�1�b .I�����5Y$�w�kh��9[S��#EIE��
� �%��'����sHqfkb� c(d�@,�G���P)�;�� C a�U4J��2>1��z$�cD!�#CCT��q4��*F�]	!��v�/�TZdY�I��w,0b^�h\� �E�JobI2�1�t� $Ǽ$��� �DQG���L�x������`��f��$� AǈW�C#գ����	���h��6^�y�H0`@`�ܩ?B�Ke�uh�0$�b�$!/\zy�Uf�_�xa%|B8J�@��хKocmBl�:&��"g0޻w�r����fFI�0�j��#}��DL�@�H���Y�������p��~�-b�I��6ը�pcQ��=�dj�y������'O�xv���(�d�~]k���(��?mw��3A��M��7�A�2�bt�C�G�_��_��_����?�����i�:�ly�s�"I��I��(IK��C��@ix���'�5��	%�Lʪ��$0ቒD/z�.B�0U�Z�A,���8�#]��`�԰@�����B/;��'� !r��(xҒ�Q`6I B��/ ��L�p�Did��:��)U�"Q�� %2�P��A�>d���x��TX�R'�Մ��(&Y �f1�e�&�!��� !f�Q�KҐIxdg)hՏ��`l�R�X�OM�X~�̴-�o<UWt�� 0v��&� xm�+�|��0�|��p2��,d̤&�F����ۚ��� ��3����N3����1�c�&��L �� �%������	�(��8&>�#��b!m�"�)%YPCBO�@�8ƤĄk�z7N�x-�~��W �Or�#ix;��1#�13(�j�(%Y%��8Y�9q�W�C��p%�r�yw�՛�˂U�S�E
ba8O�Ç�#*�k�b�,����	�7X�Ȫ?��j�a�۲X6m<��o��e��U����|��dT�f��G�&�(@v�h4)�x�F�%��*� &�\Q���R�F��h������"0�(�M����4�/c�wj�~��ׁW|�d����X?���I�	7�Z�Q�fj�d����l�h����ô=�evU'���~3��ArX�o��$6���tʎ���^�T��r<%x$A�Hǽx�˥��%���DWa��Mp��w�Q�Q+oά�,>�X��{��L����k�2wOv��s��-��|������W����og�N���<'#n����E���W�E�ޠ�v������J�aNYi�4�����\]+!��d*�\�d3^HI�x ,�j��f,�'1 �Lm*�	{ "�h��[~kP��`BFEB��N��$
/�HPX�J���X��Q��M'JIIS��Qy5��Ĕ���)u�I��-���_��-��ɶ��S�5���h�Q�Ij#��ے���L郱�]�ո�T8�ejB?Q3��Z�>�S#Ȓ6���Q-:� U��%y�5�<㑐�O�̶������@&HM�ro�%��K�X $���E��?^B,�X��sr2-�,.7r��?5�`O?��D�IXUZ�/R�<�1��h#FI��l��3Iy���)\�xI��1P��- �T�R�]Ս��d�I�.	A��
�%����)ŅR�ML�W���j��j���ԥ7EX����� A�2�5��h!!Kh!=� ج-P��u�g�WgPjB!6��-���ϧ�.�R��ga�$G�G� �#d" &p1�$H�$G,@���SG� ��!�0�F]x�XYC��B�ʐ7uы�
�	��PR
c8�u3��������צrLUK��?��*K#&��qYY)���鐚�ۦ��B�~���;�Qq�@�:]������fvr����y)Y]Q�'Ա���ZQ�h#,]6a�	��T0<FT�U>�����a0�/H�Cf'�jB��,O<�Z�5��*v� ���ZG��X�H�c��:���̩��d�>�7�I��H%G@ϙ�`� �C���#�Z<�=Ff�	�^��jŒ�JE��G���	�c��!`y�^����LS��@Wߘ2�J�l;u��Su-����:s�|Q�s����lg��)_ɯ�ǳSs���lq0�0p���������ج���?��P?�;;�:=>;���0qf���:��V���I�Im�k���)�Z�如�:K�B �eF��^��(�X�ƣ �S ���Y_Rt&�o����tonb��Ŀ}�k��Ks��yf�S������)A7��n���]�M����-��^�v�Ûo����8��m?,�x>*?R�+k}���s��rUbY���+�^�����icG���(3�[�XoY��_z�y�{���(�uyA��g2��ذ����v���c�$��OR9��|K��%6����|��70q'KBϒ�,`R-a�%�`db���_�sZW��rY�$n�<���(eu"�[������xgc�veԟ���Q�����d��@Ǩ/��	��١���Y��w��ͬ�r��˭͓�����p�eQ]t�B���[��K2&�T���9����T1Y�Aê����� F%��X�3��q!�!u�N�R/:D��q^��f�sS�~�ٽG?�������jnaЛm_��]]z2�ê��#�J���_o��������j�c�3���b�'���{�"�m���S
i���7`0;�@!���$�^%b!����B0hR�X�iZn���aږN?����0�����5.�u��G��|1sv��דZ��}� t��R?�}���-�+�����'�Y�Xzs�E�j zvfx������j����ڲ�N��d�Z��Zw��[3X���:�vkB��>梪��"nY�F��� ��A�,���H: ��&&{e�f�G��^���y�z�)�/�uN�!5)a(䳣�g��ރ��+K�N}��-v�N�D��׳oF>o��1��K��m����Ԥub��Gs9�+_á��#B���_Yvd͍V=k���
p��3��Gj�z0Sk�I�K�iP㧑�fr���[y�E:T� ��7����k��^�xI�	-�
>�R�	�;E�#���EP/���הƭ_�Suv�S�|X_�Y c���ꫬ��ۛ��|I�.�����\\��\O~��de�S�뷵�Rm��3�퇌6��kw�` ��I�A�ݻ,I�H벏2y���(�8R�FO#2��v~F�v�����c�4xLx=��@p'A<\�m6�Dȧ��!�,7�j	 ��(��.!���~���{��.�2����71i<���ݨ�J9��`�d�޽{���7BC�(6c���%%G�N��$K� Y`�4qfG ��Tqq	����_e9rШi��4x J1<9�K)hIR��$ ���r��#d���q(�c?OҮ�Y%)q�F �c$^ĐR�������d����z�!�j>I��GB��(|�#�h�Qhr�} BH���D�L�A�E�@R^b�c�_%"ЋR	�kP�q� |�z{Ɉn�N��6���ڈ�@fD8;�� ��
O��@��AG��cz$c��	p�NL�H��(�d>b����eh�f�X�!)�Y�4Yʙ��pQM��<}�����«W��_d,�"	9����܄��gB�y��Ƀ��B�t/ov�)N������v���ng��?~�/��/�}��Y���%q��#Ϟ=>����-�)<y��,d�$��F)Ń2��H>K�GzS�r������&m�S,kt�9+������L2i�ĕ �@��T��a���i��N �M��a	��D |�zd^�@�<
���D��т���/���TV%5�`H��1'��'_�#K�+Є�ˎT�����62�	��G;J4��p��8�h���N�TFz���<�!1F^�}b\��x턧�x@�h!�y5S�V'����� &!z��E�GI/!,L���iq�t��qE`1޸q">N�()E��� ~�Z���f�1�"9Z�ƪ�I�����Q`s��=j�R#��R^�;Q���u��un��GݴTr�z�DE$�:��� �b�kw�GEFx�I  �
��b0�+0BJB��`b �Y[��/z��O��/_��b]��|lÛ� )�+Y�h	%8��gO�?Ww���Q�{�S{���Ipl'q;$��~!\ �07H\!@\�B:�xLBF'����T}�+-JVi�Z�zְk�w�����J�`�#��ສ�*bR*�����'�4f������	�O��Q��3�@*ͽ�&��mo��Ϗ��IpQ��Ta��EH(1)t,����x��K&``���aY-�8�	��h��Sx2��ȗ`�4�+���rQ{	��˅k�+��#�m�*̆4p�i������ߞ��j8Z1�H��o��?��*�"J���.g@K�����+�h��ؐF���``WQ�F�y�i��+�����o!{��)��]O�#��Ŭ)UG���"#���pTeE�Fy�����(�#\$��*ČG�3L�̥D�*L{!=#�/~J�a��<w$L�(�o�*%kˌ;>/.�j���rd2t�q' ������9�=̪c]� T�U`%�-/�dK��08�X
���8�Jg0��)ł'� �(d&%�/���n-�TBG��$K��fA�S�ai�T,���$�ॖs��j���1�QV�E�/�ҳ\Y	G���r536<��`,�!�|uҙ+Ou�E��a�G�Uu����_��0&�����4��9ZK�T1`6,��Lҫc4��VD�ҥ�/!H9���iL�q��Y���A�����g�/T��ǔ/p�-�0�p��99w��1�}$:~��X>�Ҭ� ��΁玓�lv���+&Ch0u���i�Q�1˟U,r��#���YΖx�(~���4FHI&0�a2�����/b$��גK�r H���}��vTLG3N��\h�8�8d$��R�(C3Y�څ���D��Y���f',�`[�𵤔<%$�'MU�,O��%�/l�
�H���F&p1�5c��-��&@���R��6��RV���-=�0��|6�L?W��)�D�(#��R�����W�v}���Z�uU��{;��n�}�s���/��V�l����#���-̚$��ƱqԐ;jby]��&�2Ҩ'9Ϭ�)�j�:��{�����!	L-Y ��^e�I�[A�����_|��[��������ɩ��u�'�f���]=�������������7w|����࣍On�����|��.|���ر�z�G����&���Kl����j��"�K�J�o�h���3e,�_����Ҧ��]ጻv���o�ݍ+�6�I�������3��2n�|,����{�n- ��;���oْ��2����0�嚐�2���bOy����Ϛ�Q�󯟻����~������l�tҏu�/��T�#�����90�;^��L��ѣ/���{���޸q�o?��W_>z��c_����a�+���_G�1Ƕ�T�3�Y�������}u͙u����_[�����8l�N��
R������JW�z���+W6�}��'Ξ?6�\��an�g��Z���������V��Ւ�R0r}#w�.�x$�L�7÷,5�p�
z��Gs��bU��#
��G�"���������_Ƶ+�8GC�h;�?�`Mv?�3.��	C��r�v��ǃ4yg���mG����Ǧ븶��M�흽l�JF���+�4�L�CfzI�gNo��Uj�weK�9�%ɑ�	3���D#�I6��2r$dJ.ahP�-_K<i�H�\ :� �LH ]B��� ����0�]3kOe���_����Κ����q��l�"B�:�	߰�=泥�0E1�����*�r3�p6���K&ծj�e�D3�FL4�p��hȓro�Ϛ 0s��e%�*��8y��\\`#p�rG�f\R�/��ja&�q�αl�q���Ҳ�ėm�b�-	�d�����l�6[V<�f�؄h	#z����I�F��5	% 	�,�ȼڥ�,�!#17 �i��X�-Ifz2�QQ��=$%�Ґ�J �F��:.^�\�d�@�3
�7$����*P;�{!|b�,��B`�SBٮ��TE.�� �Yļ̨d�@n��{�0`	����R�ZT8V�B��$�&Q,��4PL���!�~"�4^:��6�X��!� ��8LY!)��36��P\荖	�|�+� b!�����1535�`���� 3}� i���x%УZ�FY�9Fbv�y1E+U���^Q���6X{�%�hc[�Ն�@�YJ݆yRx����"�s�p ��qqQr��K�L�O��"�pXɆ�
G,=1������U&m�x�TlK&�Gr���*���I�nt�����{(J���~�#�z��ە��P�"��x�s���2C����M|�Ɇ�2ʳkjQ-E"\�t��T���    IDAT?�9w�I� ���+"A���'���+��O��'(���8��T�F��JW��C&U� ��|%�ʥ�2)�RwpRv���� 4r�
C�n3/<�f�d���Q�?_���4L���r�rfB(
�4h��DS��D���Q����+
@9�	 V��Ă�(���Q�_0��a%Of5���גCi𥉓�4�A��Ysl�0��i�[�5�2)H�x:4a(qQ z�S(����e%��&r`��(F�`*�al<[��h{ku2�`�b�Z��� @).�����az��2�	f��Tz��^02�9<�p�fVC�jq������ۤx�����ƃz<+���.������=�����2������샷4 ]L{:ª]\��{\�	��:�ݠ/O3�� ��z0.��X.�|��Xe	=e �y`�zNh�lmmy���k/�d2�Zi��dQb��� U!���`���"R�@�T%&B��'��L��@(��*�!�����+e�8�K�4�a8�p�! 9�sm�%�ѓ�Q0���dY&	��r&?0��"���И9Z��@��42G�a����Ku�F�3P�?km�����\s�wKA��mi���'��d0s+�R����%����_�|�My�a_T�GM��_p�	M�k���:��J#�`0j1Z��d0�9��L4����K��~(��]�]*��J5�.�H��bI/J�/Gxr�Q�L��*��L�	H �f�L�Ҁ�ӛ+�1jodͅ*&AƏ'_�r����`�8���_���Бsq�1H�̥���J��_�Z�[`�8�ג�>l�NX�+g��@x��U�xJ��Ҡf����o
��J#� ���9��%+���g�m%P˅�)�%���
C	��Z"��n��b�|U����a�ϥ�I�@�͐CiK/Z�(-�1 ҫT�h}�뀎ї!=C�Z�1�a/��2�i�1�����d�@�gҮ���-�d�^9: �:`&6#�=Z3�*�-c.��R"�ޞ� ��jN�\9������C�7`*[G��*���	���@��&Y����$w�	L�Q*3_��S,�0dVW����DɄh	Hb�I�ި"&`���d���`I�#�q��[��Ϋ��y�R�5��2r�p��9/3��*V&T�Yi�Q�����Q4����^�@�Áˁ��͋@o�$��PV+^��y�,����r)Vz3<S����!Z�K 0h �j�Xr�ӈ߻}��������EhPVe 6?/��,�Z�Tʜ�{2�A=3wR��1���R˂
�J#��;"u���Հ�� %����8�����=��=��a7���'	<�9���������g_|��ݛ����x���O�G���1�D_��!�o�xZ��nN�p�$�:�b�$"�V;��hd+��+-�l���F�@�x��0jg�����~{����}��g��?}�`��)�j�;=�+&F�SD���'��gGN>y�ϑ;���Wm��8پ���ώ>����|�������Ȏ'7���<��1�����X=����������@�e�D�eMV;�F���Y7X5��,f�������޶�v|!9ց8�Li���������sM/j.} dV?͵Q���oh)c���Dci�E��-ǁ���Ϥ���'��=����N=;���ǟ>{��3'�}�C������z��0�9��֟ٷ�Nl��8��ƅ��x��W�|��'_޹��׏v���GO��a	{��G'Μ:vt�g�N�9�x'��g����/�oxjy�3�yqp��l�U@_�w�#��8���n=zk�k�\�x���O�za��u�p�,�a�)�_�pgo�7��ӛP�75���D�1g�4������(�e%tEe�LǗ�������G+�����C��8�k{���;�e	��ѹ ��=cc�ꘚǁ��H�`6��Q�_�jrt���_���p#�7;��;sNQ_?�J{bG�E��9�<~�`������,��d���Z�Q`)A�Z-�� _!�H�KV�L!�/�A����`ZJRmd-Qh`�L�KiDϊā�/�'��d	�;zb�³/"��_X�H��Rϕ�)6.�#(�|�:\<ڢN��q���0�j�H�$OɴH(W�����Y)��,�%N楄�U��ŖP�q���dғ�iY8&�v/Q��ޠ���@�ޤ�r�2�!G Kg�⡱�DA�S�U�#+�B�Lɋ���d-g �H��\�|ɐ(h�L�1]��a��v�
C�$P���@�&$_K�D1�0�h����eϓ��>��(��*G����E��LX�*rgB�i �c� B�/�-:�Ώ��G��L&Y�|sW%r~�L�3�[2a��O���; 3�9�<y�����LcYӪy��([�y�r�7h,�%��\��,hq���,C ���0G��,�]\�*8���Hof2���e�$����4Xya iJ��b������IJ�|���X����	)P�Xl46^�$+�\����Y9-�:TD�
!�Z��CJ��M�M�n��ܹ�S�u��Z�@B�7�"S�(�Η[��^�|9����̔e¥�����_�t�g�F���I���n��厢g���H��D9pQ� �S�R��@8�@ J��pT�,���u�˕�����?h�q��ǯޕ}��G�o��"=���RDG�f��ի�1����/�J3�_��W?K�\l���h�u�	F��Go��D=�����*}i��Yxd+��C�M�4�#�)�^�_<�fɯ���g�4����BFkᆒ���aYQ��Z(-��B h�ծ^KV�h,���;X̔L)Y���LC�� �4��sGY�Lj�IJ`��@YxM�aÑҠ�IV������-Q� �Ê�l)
=l�z�A_̐4S �|��V�4� W %~�|!20TL`�&�l0���aW�~�д�&�/|���в�R\2�e&� �z��8��Ϛ�<�K)y��1K���g�
�^��;�c^���It^�-�C�AQ�eq�,Ed�����d�H&3�@��&!���D�	�: �1�JLD��7��-)�e��Lf��-72���aʍ��T�r�䃳���բ�[[[��Hb���Y�J�$K��қ�	�p�[s�U+�V1s|K�#k��y0gKi�?G����RZV~J���!�јY%�{3���+3�V�HX���$y,E��da�wE�&�%��u"�`}h�9�qK[4����4��!�v�M���dii_�x�0$�1��}��i�7(�d��'{�g/j�(��j��vAV�5X z����K�?�-)K0^�+洎3(a�w��DާT8��Hi�Ԡ�CI�Iυ��b�Ֆ^R?�������mu`��w�!UD���+��`�?�loĉ_OD��#�ٱ (�E���2}�`�4d˅R 3$�|�)(!YCҐad��"��&�*If�$�Y��F�a&�=-�s@�TJ`l$��n��1�����U��e�4T���v���`1���Z�YB�z��&��!P�xu�R��Z�8c+��*MJ3���L��������ɬL!?�\�^�`��U8&3����l��4!�$;��i��i&g�E���Θi0L�wV�ܑ�6S����
	��ɮ*�H�%3M��u!�
���x�<A�[�%���PtJe�
1�5;���f�P�m�L\J ^�eHI�*���D��#CEF%S��`�D%���<�4L�0���e����@ʡ���qa-���o�4�@4������.J�R*�|�r��l)\����Ab^���Eғ๗96�|��螺 �st�h�%�J,B%�Cbf�\��!�*�;J0�eƒ;+AL�L�c+(/,`�,E���J ��,� �f�R2,͖�� (:�4��7Sbp���
�#��!�B�<	�|Q0�K �Е@t�7�bP�a�Зd�R�Li�� �h,�4X�P0L�4	`Qѐ��o�U��z�J���([3<�0�J@b�����@��h~'��gs<�ٻۤ�~�����+�G��ʤ�⇧���#G�-6��E����j=9�W�J�^ЛI;: ���6�tK�:�C3����&Cm9��%A�	���9����0:����W��i����{_�t����ܽp����<<���_���w.H���џ�7����~�����num����/\��͗_=x��/�y�x�>�^�89���{��z�b�D����W:��G����k�C_�Җ�Ci�������^§7�	\j�>�����v�@��}�HO�YCJḓu	S�d$ LтY�����c&�8��h���������=����'�|���'_��ի/�x�Km;�˟���)W[Y<��ʹq��Ƴ#'Ϝe�£�_�����s��������>?5~������ٰ�6�v�s�cz�~���_(��J���Xc���Y�"�����8�t�=]� l�7޼���޹r��W.��wS��[~ԦO��ock��=���y�Ԋ{_}}��M�Gַ�p$th�k�����5_1`�^3�����z�T�s�o8x�ゟW��1*�p� 3�P�f�K��%@�%B~�����ߏ;��.)N_�v��|����ޫ~����c7�c�x�Է��e���??0늢���NO��8;�^���$T9�+�lȧ=Vb`�7�Y�O0�nt	�܅0�ǡ�CHKT0"�����o�`@^��_K�_"�ƋL	fHR���&:r�,�tX!�9qҥw��NN��b�!�a�l�Ή�G��N�'S�j3���>ڈ��ι0i`��D[u�\2�K���T�j^�|�)aH�0Eȷ%��^�ȳ���$1`�"��s��E).�V�G�\v�ʼM.
+�'� �lY;�f�1�
gvЁ+�e<��4 a��4�RͅL0�k�ѹ\[0�QE���0������H�#�e��yY$o6�i�0�@�� 7��cC��V�b�o4��������"�z9;�*�-ĝ*�8�d^4zbH�/0��z�ob�#�ڹ`&�F`����-�M,���li0ғ��L��iJÜ��i�4��j�L���j��,9�_�	H$��́-UGF��Ʋs6	�&Ф�iT5�dȥ*�Q�45�#�&��wJ�zE`*n5����
�Ţ�a�΀#"r1wp�Υ(����NmJؠ'���W�(K�qc��~+qc�aTfoE����\$�����݆������ %ٞ��H�sD,$�/_��͛7��r�}��G(V��J%��������|Ж0N�d��o��^�O�1�Ii����_��>&uoy���x�K���u=g4��?���/�qu�+�����\ىk�7+3��#{d���v].�I�*dtm�k���Y�U������7��<���q�1�-'/��j����7#8�����8){���ow�vR����c�̤ݤ��Y����ĐG�&�	�l�c�	�����ە=�y]^=�R2�}[����r��r�Ѽ�w��,��B*�V<�v�9=�[&� w��=�ۺ��p7s����V�,i����f�?����ߛ��d�[����X#��\
�)�YFϙ:AC�@GDjdSn�x0�=D�{,�Қd���H�T����r��	�{ۋOr�G1F�G��l���ͣ*2s��-�D��>����*P�������1�Ԅ�(�/.f>���#�IZ�cI_2k��A
��\������uv��@&���]��>VV,���]x\���h��\���?10��Y���ᬇ8yq��+%P�\��YZ���sY&���E�V������j1�R�f�-��=�y�oz���<!�2��/��cx$"F��c����Xa�a�(��jZ�����칑��|������&��D-Vy��)p����)�#U�ӹ�hqF5oC�
-�.T�Vʹ��oF����<d��2�1"��!<Ї����}����
\��P�sZ �k�4�N��VmX��c����z:�Gi�=�g��ʨ ��e���Ũ���^�D�:�t!��x��&��n��g�C��2� �9���QFM��6�޷C���7j��eV�	&ޜ~o2�=u������m�[,�A��x����?��Mj���=f�{��40�Du��M �$)���k="d��Ψ��q+'0��0]f^4�@߽ZvL��S�S���/���|����`�^g��8�zlSX���57���g�;f�=�%y�8�6��i	-�^�e�5A2R�.��Z�D�����5�tkl��~i�c<Ǵ�z35�� L�F�k]&��Y�U) �1�7�1N[��ml�è�2�ߪ+�jV8�gHU*,���*�>�Z<��|zr2����GZ-?����WP�E}p��ʴ�*�<���>�	��q���.��GH���xҍ>$<��b�|2KUG0:�ّ8�JF�ʦ*�!�e96�eĤB������_���@8��&�un�=�����"5(���-��|U3)�0���.h �k���� <P^װۦA2bw��n�S�i�b`D���e"u�O���)p�����yE���krYz��ņ����@�I� 6�",aa�OӀ�)��Mpf������'ܸ+F%�Z�䷹��R��s�e�p���46��W;�B�X���-X�e6H�� ,�	��هFe��5�z�#^w�|�%�����mn�F����jo�k(i��4
�p���W�OF�-����9�T��az���p��j6��������w�N�C�Z?q��b�6�K��(�tG�W�w���Y�/
�J(��t~���t�w�4Fӣk@��(汫���Kr��>8�k��G'I�ބ������C��ˣ^�W�3��p+��6��5�v�;�}��"�ڇ��������d��C�D��/��������6\eO��\nȳp�+b����OO��}�>��Y���������w�
�[B������>vN��J.�v.׊*��w䚽��N�W�#B�TUNF�Q��p�Z��?�� �Y��j.|=�����"���A�͢e�g?n�d�t�}Z���8vŋ�jC��d���Q�e�ю{W��{b�sw휌d]u�)�m�I��zޭ�w�<�Wp�8��!n[S���e��]U��Y'���"�_��$������3���Y�O����~aS�������,�:�:�t*����W��ѦB�*	���:y�����rA�b5bc8�mJ��N�������9/�Zލ(��F��g�X���~��j�)p��1+��o�nz�cx���q2�^�U�sWh��l�쾰��#!��4�*����it�&��+��V�2o��J���_?y�e�wW��#���E	�+���W,���k~oy��e��z�����o͢��j�J��n`&����f�L��Lͮѳ�T:���ƚW�>⼡_$mԈ��Lܿ�6�R�[:�ez���T[�h�$�eeS;���j[jB֨|�[�U���m1�=�+���!��I9F�5��$v�#\>��K�Y�������N
t� �'��D�!���Y��!���Ѷ�ڪ�D]�������#	�`Jf�.�6KOPjQ�$0��>e�-�uA� ��1�}�۳rH��`��:A��r+�2�� �NL_U���cH���a~D�%=&w؛- x[E��0u�(BPL��_l}pjJ��Z[��7�@~|Ǚ���-�f�>�A� . 9���e�ӭ�`I�\\2��~!X�ij8(�E��.&x-�3*v!��f�rA�i$��L�!U�+g��A�H�}b�!���aْ���*o�vRs�������hUII)2#��{����*�6 !�Wb����$"��P����bE�L����'�x��5K�M!&6��x(�rWM����.En8ҸIZ��t�}�I���C�ѻ0 ܊G�#�-(��R���*Qký�{@X�!�kXNRe`���G��4f��;{�`�լ�w"8�7�j��w��p��7~F�����'8�6�L�O(BW���� ��� �������
��6$�~~l�M�����:�$�%��3>z�K�d����ǝR��Y���;��lK�Y���G{�
��.��zYW��{����-������N��(�[]���O��?>�6>o1�� gr�,b�����>�\�4gk琗�ך�R��C֬ո6D��ɯ�ը�d6�����e������p��x���2���X�6#�����<o�K.���wa�s�қn�����%<)|K��A%�j[8@�Ώ@���b*ZL=��&#r�,'[��5F@8���*}~=����_��$�H�,���6ޒ3���y�=�)�W��E�2@�0�V����d�@"��?<�43��@:�$�tQ��>���������]my��UdoT`^�y@W��̔紾���*@^��|V��"��<Gg}�����n���Cl�nk~�V�j/C{��wտ������kIvDŵ~�Q������_��o�wkO�s�W�<r Ƞ~ǚ��+��1bē`��N�1�w�G>��25h�$oL�$�a�����zv�S�Ƕ�0&+��j�^�٤d����f��S�\��ٙ�����$uO����xz������P*�9&	Y�''ԱDZ�^�g`��;��;�|Y�R�:$�|�g�c�;�o�R��r!����Az���R�4/'5G�r�l�Zv1�P��Ud�χ�������4e�O��S��V��&t�4�>��VK�	�%V'��䕆�Q�H#�2��G����Q!��xf	sm���:�>��Y�S������}vh*�C^/�e�%�H����[���"�Ȇ�2��%�j��%�d;���!.��Ha2[>��=��O�&��\��}����	͚������Ɏ���M\t�ʈS�;IDF!�):�Ɨ�5&�r��3��vᲸm��7̉�٫Q�)�MzL��H��I(#s�r*B{,E�o��< �&��][����z��n6�.Nv�\k��>��-޸_�(e�֣HRs��g�8�ڤ��4�αjh����/��5c7��K��r&��lq^x�a�Z^qg?�\�CX�9V��[��'d��Lc�I�	}ǁ%/�N0�J߱����d7��-��>>*&u�� `Է�E�]��`;��FfNI�Q��j����n�t7u�	0B� �TbY%���h�kL��q�#7PS�辡a�"���r~B �(�?_sc�V~�&�p��%�h�$N��?2'��z���㳍�P�ő<E��O�3�CZ#D��N�-)�*X�g��;b"�x.5������{�s��`��՟㱹�N	��ci�.�ГZ"�9����dA�m��i�-�D���j��'H�aΧ };���~6�i�@���  ;WG]�D�&�����`r�G���c���{��?n���;��`��OQ碛S����:H��m����*{�e�u�%�!�T���;\�a8�\X�CgF��(R��%���Q1"T2\�k$�@���_�]���\���|wI�����ͱ_�Hm��e�Y���Ż�M�[����ηR
۪���,�0w�{-�w��u�R���%�_@壆�Jj����%}׹�����jէAULYP?V��'��v�A	�c�vf�x/�u���s��?ߟ���=�5J;_9�6M�rl����DƘ���K�\��@��ab�����W��5Ǟ����],��bM}�w����{�*g�I��h��^�0��:����u}��K?;tS6,Q�?3��گ]�����z�!qv�j�'��)D-����l��=��Ӂ������\��Bc�O��~'�[��x��r���%�}fv�����gn��I�j�c\�VS��Af�W{�K��Ǽ6������e�W&+x�~hKV�	��fh����d��v�i!%��ȷP�A�؁UJ"�NJ��z�$;t��we�i��6�w�s,�]������;��	�<���3>}Ӣs`�y&Wb�Y��ݍRU�%�q��'[}'kVm�FJQ��R��wX-���e>E�'�r)�+իe��?�k��A{�g�X��^k�S�ڹ6��ˀ���f=��e��"�\��"O���}"�E��[�ٜ�l�ky.`����)�-�g��:���j8�$*���"�K�?�~RY����t�3���q�?nkOrJ���5����?
�c�T=�n�0Ce��~Ot�UC�a5{6��I��70�/�?��.�-ģ�4���l����cG+r��d�����-��7-;1�)-+���w3�8�?��g�l1G���4���t�o#�>{����m,.iY�|�j�B`]J�9�č���.r�I1�(�zC��}ͩp�]�̦?�`���/c8>��r����Y�5l�.7S�vD��u��ˇ5��W\)(�<�_�rՒ����mxw�֮�l{U�n@��y����K�FzIRv���q�Rr���ˑ���`���$��[�z\��eq=_����"e�!t.��^���X�V���{�ɘ+���Ѿ���C� f�S3)cq2ȶvi��)�x���y�x��<A�ނX����o�Ϊ�P����K�@Ur�p�pQ�A��Q4����Q����Mo�Y�9��{�Gޜ"w��}�y��:����֫I7��J�Yt�k���O����7�_�p?�=ȅ7�w0���h�#W���_�W�c����������ؐ"�
����M%���i>�h覝)
�?�
^~ip�| 
��>
��9djC����@X"T��f[�L2=�Ó���?S���ϗ�|t�,�g4ѣ1��j���P�Uk}�I�� ���ܣN��U9�eoS�XO �� <q� d�q*1^���̍�L�TeC�Kܽ�j���:�l�����N=�YrH4����m*K���S�x:5~�^��o�9,���M�z�X��ضvN�����Y?�e�ip����\{,�ષ�l��|r"oA}�rW������U�*XyGr\
"9�0�=9�o��ٗ�9���-��z� \J�����T��8�˼��Ðn<�u��d�4C�r_���9/ah��ma�U�]VF�Vk>�2��M fސ��FLQdr�h��W�\4N��Du���f�u�h��B�p'ieb͋�7An]���]6(]��W�a A&�Cވ1g]TŶEG�Hg����-��(�M�(���g��ϲ.�*���K��k~%�К�W��˵ ��,������$NoFƆAO±�a	�+�2uh�
@�����,�~���*ۉق�u�9�+^ow�|���"�P������������3���XWM��lƴ=��_���-X n.L��cp#s��-En�a#�9xE�A6�hx ����~�~����=�VG��C�h�C&ܯ���I0�B^�nh�m[�4T�f��;��jT����ǑB�X��BD��y1_�S�\ |�n���ş�o��s��`P��9���P&{"/��W�0 T(.��	"��p�����e�Ш��\�����l��
zY��>�7��P;-GN��s`y�y���޶����mXjE)8ŷ�"I�kۮ���f�ʵ���7X�,�$�݇|2y-��X������(1>�2Q'�Ը��Ͼ(����'���%dF���?�>W�. ��_�H������b '����4͌u�sY*�A���^���c���๱YR��eZP��:��ř��+	 &[v"��19�֭�٤����ժ�Q5�:�|o�dv�0
Q����F�L(��QQ�H�h��YY�3���X��e��qNp]�9�mc�P�:ރ���EJ��2�U�&�R��ǧ���������$f5�K�v�:�er��ᨛ ��R*�?�&�!�iJ�	h�xi�q�A��m��-�\ ��$�B慧��ɩO{C���n����M�,s�d6�:���C/��%"7�G�)gu�ᡎ``3c~U!��Ƽh���q!Z`e�G�s�_����/C�7D����'s��X����	PE.���1r.&�r�+T�i��?y�A��h/�z��{*��"ܰ�;��K>�'vUwN��G�hǿ0yӰ87*6 �'���B:d��a��lN`;�t����a;��2���R��S����0����ka�}=R�z{�r��w�հ=�:�;yӁE�Ȅ���vN�`�{Ŋv�T�'	
:<��=+8�W9��u�H����0iz旅~��$i�x�2��mt��#��F]���������U)F�E�sV����w���t	ێ5[�xԎ�/J{�F+�L��v[�Q� 3�h�PH�ƞ$��> (r^^���zO�<����g�}�{�Q����#7��Ʒq�ص
M�I�?��6���-��&Blތ��ܞ����E;��á��o#�ƅ���.?S^QOc_��.X���!|�BWx�x�#j��G�{m���q�~���=)0�:�8�*G	����*�+�N� �8R�O-�樤.}�H넚:��Vd���I�l�kz��:ϋ2�D�HCTû�[]w����$|�
�2�y���^�%2\���𛩟��N�ũk�k����7H���̉�w�_��%�1VNs'O�c���⠢v�@#	���XЕ3�Ę����(��a,�Br�"�l�����)��f͜I�@��XN��
����`�$�i�wA��:����(�7��h\A��T���p�޿lT�b�5A���ލ��4�I��l�#XX7��aN�+��n��`�{�>��5��ٖ#R�����ۨ!���O����#�w�giw1��m��P�";�8��@���R�w
 � �9c���t�0�-���`�x�M�A宮;q����C}��VX����-�eک���}����$a �n}�E��r0I{#S7��<���V��3�;�#Y�Iڒ,yEPv���m6ndRf�T��c�(��7T��;��̹3�>�]qx��Wfj�!��b韭�q���Q%K�v�Io�X1����> I��:� \�E��4ݐ��fn��9Q1���%iۭ�y��8b�Dt�f��X4�Y��nx3�����"$�>k��0��.�/�Z5��O��B2���V����{$�A����yr����*��5�[���n�`�[�
�X.ˠP���~ť;g��!��KL�)���	wӜ$���1�_�������G����-j���LU���Q��'�5���F-\��mB���K�;@����G;��U��.�.D7+}�i��������Ǧ�q���P݇�T[��[�+�4��_v���ȟ�l+��-t�r���~�WK��١`dr94�5�!,�|5N��=c'm��v(�
������yV� �#�[�P��-��*�G/v1ڭ�'^33_�T^U��,��� �TLMa])Z��f���"	I��ހo�'��>zCz*��;\R5�#��H^G�p@Y�Z�b�@Ш�TڔܡR��5�b�0\*���m}�Cn�L�O�
Nj�x�S�R��''c`RpL8�����]����yʑޜ�l)���L(n���GW�`A���c RJ��aF����v��,/5C����l(W~X?�&(�]⁣���΂LN��}��!�p~8��]��)�;�"$�d�ዢ�y���i���@�7��Y�:��C�A�g���~Or��oR���R<�L�+���]3�\��ԑ��I������[	��΍��P=�dka�B?�MJ1��1	�#����:'.�� 2k��d�-�I2�'k효fǾ佅d��֭�_����u�m�&���E`�k+���%�^��>�}D��Pw���Rc�Ю��C� >:�`�.E��(툾іG���Y�H&�<�%��+��������1[�1[�M��F.WA}9\RL����am�ڲr�N���C��	"��It�/��t���9��.)�q}�2�v�9S�7%� �@��<R��Si���̗J;k��`������x�!W�5�ld6;�o�R/�h���	�i��Mٹ�~�r��u�ɬ�q H��}6�����aLK�62?����ZV{bJ	�c��D�/��X�� �Es7J%?���W�)���5x�qo����o�Vu9��U���)�6�q
�*S�!3�&3L,&�@��A
Z�K�q6�W��M��/:/,@�X2涓���|��e,@5�l�ȼ6l�^N}3���GV��tr,MK�?��A�D���M Y�0�za�1�vqZ�J+[Wɱ��PJ�e3�^������JE����������u��a�.��z8k����X�J�$���=���,��.73�vą�.�"%&�0s����8��h���J4�tX��[�/�H/��V��6==�DW=�ѿ?��/��__����{ ���K��֓\��#&�������?��Z|����&6�̞iH�����u8}��V��"sP�ݬw�Ќ�ʵ���A3ǔ����m�?AZ8�!�5I�������1N"����JkL~*!3�e�r�*��Yn̄�e�X���s��d��x^�b��s2��4{ID}�P�?��Ew��2ќ��%�s�c�g�"����~�9��þe��֊MjG�{����+���ϩ�Z��Q&��ȀJ�ǜ,�-����\���p*^�x6�i��9|�HN�E�\W��Ņ�F,m���{��i��$!�o��p��+K,*O&^�S�J�������¾�rN�y��i*[�f/��ܸ��{�	{T����]�D�*ӽ�P���0uL��Sﴙ3�H"�8��k���d�%�~?_�j5�}���T
���s���h0��,�SvGG��[��W�0�P�)kWD]��ܣx�4�g^�������O���?�0��Ƣ?���uc��8c�����#��)Tl�X�S��8��Ѐ�-��Z��b�>�?|]\TPN��m�=�VPJ8�AM[���P�"�����n�էƢ��Jז��Z��_+�p�&�8&��B�n��V������"7GOd/�Ǝ�p�(`�����|.�	�`TR�4?���!��=�C�$���I��d�i������:F�=�fEr����z 7H��}�k�,�s�/�x\ҍ�o?����(L*<����S�LĖ��;��� ��/��{4�����=��L�z�\�w�Y�~��پ$�qJewѴSiDڍo=>�,bS�ĭx}Mj�Bi��Ч�<�[=�2Ly�H5wם:O^�L��3�~�Ll�IA�̆O���?$NJI8.��^s�3�y0�\L�(�.Kc�1�)?,�=F�H1�Y��oMH���)@��}8�,j����cMQ'��6g,�
߄>�"ʈс�\��T銩�:wU�`P��5��P�wO���3�����b�e��|��Osw��+��wH�#�v6�&��m��a@4-�[���c.p^����N8�B9��%V9��Q(_���LO���iy�HR���CerФY��(������k��ڀf0�`�g�5FJ'����3a0�?3��B�����a�^Cm oŉ溗�~s-�1G���E��M��P�T��1oIۮ[+nND7ҿU�q�{t��/�/ ��\[p�1�!�R�'JӉ)>���72��7������Y�Y#5f�G��>��/��&���nDp��(�]Ѻ�tǰ�E�|H�8�Bq��.=,��Ò��6gFA��a� `�#G�K 8>/��>�.f:*����9�%���x���D[�8ma�Wl�
�����?;�������b��O�`-g{�0m���<)�"�H��=H���Y�)���T��/&��!��fXI�{1��+���r=��m)�Y�o��7�v��k��Mal�+�]s-�j�,�����Te�Cs䓭��Z��N$��8���Z�z�20+�x�&`/ �ؐ3��tKe*,��6��r�Pc6���59�Gc]Y�%�����T�o0]	@%�f��a��5q�D�J�W�Q#�z�^q��Z�ݭ@�z�1�9Nw�VA����_��'i�t���g�d��o�Z�j�.�4��p}���<DH��88����6S�"٥���%�I�@X_gRmy���0�I*)U��Y��e�_����mU�oY׆�}٤��4����Q�&��b�3���>59��R��E��X�P��������,m�����&���d5�]�7)D�Tש�7G�ic��D��l٨�t. ul���Μ��H*4�m9dG	 ���(:/�d�9W������\^)���VV�K*�H��r|
xj���18 *��tH3K���h��/z�yX93��l���z�M�F�q����?��m���Y���0wX�+��LT�t���Ӈ�T_X����{jy��(�,��=�Y�����m�ΐ���~�!#lq����|(��Ħ�����vr�,�b˱X�%���!2K70iN+d��5��c��1�/�Aԏ�)�|/����``Ѯ̞uH�E�_b횱'��}_i~X��V��wJ�4�N��@�9�����t!w5_���ey8ɑZ� ���������0H���#GG=@��z�G
�>?�qEb�nf�Z�����6|�]3"�������,/�Y�R�I��gPj>TT^+,mU�A/��,��(��u�Ϫ,n���b�;Ǳ���c8�K���~̍޻�¬f��U΀X�-��!1Hd�k��s�$����o3)���D��~������z#�M� j�^I0O��8����U��%L��~$����EE��>\	3��R	rfB*�y���2Q�����j[��j�ol����
tQ&������rq2�����eP8�K�#Z=y�Cv������$�6�y���mշ[5��ד!�xX�-喘>h���o�V�������x�Sc���j^9�Q˘���0+�=&Zm`�+t202@�	O`��*/���mK:�5���<.KNgK���̩n��
6hZ����!����<�

שk���r���.��~/Y��������1�m��ι9��·�e|X��I�s//�J^}�+�T������>.]y8ެ�8�y�3e��HM��i��i�D�$#�iΏP�  1��ΌtI!Kv�nK��d�M�u�s�@˫�fYZ2Cׇ�ʌ�".�άe���>�G_@'|�8�����Dȴ�tlW�AdtY���������?���s�q�
/ۿ��Co���:8�bVC #T���b�����K㳿Xy��YM\r3��M��Q����w�Q��x84�����M��-iSf	��O�-�����@-�L+�c����&߷�'��)�˾���Y�X�!&�5sYg0dM��'�������k3�Ǉ}ӻ�d�Mw"8^�ܙH@�Ol��E�j-��Ø�E��(�;T�\W\w��ԇ���L��!��3�P�۫MҊQ���u���w�6B���i}��iY��ğ;�~�P�J߳�SIsx1�7�S6�k3��������� ��K��c�l���3����#�n��i�So�����9����$E�;��������or����ȫy�ד.� \���#S6f��VG2ܺ��d������}�4�ßn;Q
���M]�%5�G�	3�U���Úk�ԥ�ZD���DY��f�����pހ����Q�������7��n2O,�$9���)��lUN��S�����J::�m��GL,}gv!PjX ��)�p��8qVx����G��|MA&����(�?�.��v�IE�M$o�Ƈ%P��/fnx�#�&�2ϙ[�}#s<ΰ�&�h' �	���,��/�2��Kr����kɝ��Ҧ�e��\Q�T'zZ��sN�R|�]�C�s8?\=��+}}㋞����X��~��Z��~�ή���OFF
�1Q�#*������=�W��j��%��&��Ti��8�q������~� �f4�G���s�쎚e�n�%ߌn_D&���puIy��yW"�����#��3�L�>��Ȅ[��DX!3gw� �,X�z~����*Yg���h��z��t�G��i��hv��ܶ/��9:�W���g+�"�ٹ�eb7�V�$��h��xhT�!o���z]���QZ*�S�W'V%�oޢ�Vū lh�Iv�mL4���%�N�����5-0�F�՚}i����>��۷옊zl�0`��ݣF|�$�=2��.�"��]��lL<�BB<�挢������V䰳)y@tT�	��ED�*�A��^��Z��Uh�8[x�f�،@sB��@Bڛ�Bi�Im�����M���7���Ź��5�����
��Z�?���5��:��k\}Z�A��8b'�C�+-2��	�0��`���o\&G�*�Ǡ��(�e��D��"C��!�]������=o,4��)�m7Xw8�:Yu|���.Ugr��X�"b9l�!?Jޛ�E��=$`eg����4�M�`*F�1��6O<lT���s���s�#gk�ǈ���'��/�D�T�Uw� �Y��O`��%J�d�d���V4��rG��⁄m�HT����ے۞Q�:f���e�)��}S�0)����?y�Z�@����sFĥ�i�R�K���5�5��g�Ǻѩ9YѴ�.�oG桏,�*�.�Aa�5��6n&n���.�S3�tu��+<�V���:�lx&��ݩ�0���
����|�4�j�,���R�*"k���3�s�U��O�	_��_�>�3M���4q�8h�-���k���]�Y�@U�]�p�f��0��ߕ��x�?#�i�Wz�N�ܕ1:��.6�a�x�"�:�R!��[��{�{B�Q\{$n�n4ޛ��QuT΋�o&cS�@��Z���[����'8�An����I��0w*���,m������mu)
��2���P�&��	���O\�nnd�Z���(e��&�(�á��1���IBͰ����������E���`�y����+c��I�}p-U�����	�̾�=�}��GF>�	>I���$�c'X���=���&� S����Di�u]x$��i�6ѓ*;���>{���FV��#������by`+�Շ �12s�uM���e���	���A۬Rw���YH�~L??/4|Q��H-D�z��@q�g��-���CT�mHSqr���2zs��>d�����L5�H�Q�^<|ڮ�5.mM/�AK���xj-��-*����t8�G�����֙��d��r�:*��'�v}
O
7U6⏽
.AL�H�����qs	6�{̬��?Z�7{�ut�@��ȕֻk�ZT�9E8(7!������BM�n�0��S�ŀ1�ס�	������"C�	��	B��uf���$��*�uhԼV4��eg��$�k��ewՋ�1�P!�_�/�e�'�E���!>TK��DH����k����5VY
`�(o�C)��sU|�A��2$-i r�b�M>kD���e��^֨�go,e�Fyl{]������(/��u�k��c��5��O�o� 5Ni[P��e.��|"=�Bjz�;e[� �y䧅���	��0�*I[8�
5E� �Q&��Ypq�ɸ�*��l'~�ﵗA����"鍳�����ٺp��m����ۑU�/�����Xq�Q�J.^7�cBгQk\&3��+Л����� �PMu%�hn�
��A���"�	f�!�,*H�=Qh�!�����O����Rd�m&��71�r�T8��8(F�a_<S�^���ސgG.B�@�p��(�7��n�(��*���a�FvEP䶬�K\&��%�b%����W�@\ߠ��b�Q�bo���UUR��T��}@p�y�ϑ��9qC���ƪT�֗ �#��%���?�}a�Nȸ.ٻ�8�	S��zaok˾pg\B/�F���� 2����P�@��8��`�r�7�r��.f��(=����2�t�z/�kE���[�����&��?��܊\l݈7������o�����>�����c�eA�=o���Ĝ�O��ݘ)�{
��v/����xW)�n�5ч]��j0�+c�X/�f0d�c�uK�o���5�~���O���U"q֝�d���ͧ:��W�F�����'Qr�R��NbB�+�=�]���>�F�>��(�z+y�v�<����/���I}����*8��>�в�Sk�^���=���f���ލ|3�~����<W;�P���߃)��.X@�ì���F���h��܇�����W��47�S��v�͈\���^Fjޖ��j��k��#�eԖXp�޸o�P����xY�Nb�����Uch�P��
���F�qߟ|n�K�Y�Wc��{�� �R�x�k $��XSw��Fz�Z��������ڍ\���5Zj{yw���q!1�r��~��q�h(�;��iͿ0RQfQ ��Uom�̧K����g\�ȏQ�y^z�����h�\��7W��EG���bp���G��`��%bN)��u&�?R&�"��P�;��B���Wq(u0�s��."����.^����*8���=�qS�S>��4�a� ���6PJP��Q�O�
Uj���{�zM<zw& �L1��xڲ�����ր�N������u���L�Yz����[��sm�P��-K�3 +�"#	ʫ$�H���RpQ��/�o�Z|�r�q���`=�v�n6��-x!RY%<�Hs����3��ͻ��HY�@�=��8J̓����t�x+4i\�B��.�i����څ��Z�wj�ĵ�.h�R��X9��e��L
�4R��/�D�K�Z¶٤��)�0��P��o{��vK|O�B�|F6�Ap�(ݎ�m�}I��X7v�`�+�s�s��_򽽽g>_^Z�Њ��t7Z�)_P�=�&&�{O�7e0���5��mt���V�i�4��M���=˥j#�
�)ܽ�#AQO�ǓD?�k�ږ�m��������_kϿ�����H�<��1��V���g�@H�G�cG׫4�������v�=�/V߫4X�����ztj�Rĵ�$zy~�ΓG%�uZ�����L.����GsNp�Y��'z��Y���%_O|�����3�a�ib�}�Rۑ�5�&�W(�1�u����������AN�M� J��Φ���m��$��z)'���#��t	)!�gV�1'�d|dۦ
ޏ��X�뷻%5�C�P�(��@���� ��_V(������ob��
o���h�1����v���yu�b��I����r�G�C@��ii���1F%�����-T`��I���>"��W
?j��npFv�y6l�k�.�����ח`��Q�ի_�Hfh9Rm��{Y$!c�jX�Wj�ۭ\�q��
��&�\Y��.���I�I5� �S�G�*��Y i;\�܋�o=_=���2��u����h�W�b������,�c�#W��cؐ2����{n���-ռ��������>[�3~���C)	�_�f�τ��ͱ���B�Ms�j}��jr䌶a�F�,T��Z17�r�(��	17�"w_��J������<���y���܃5����:��"�n�~\ڞ���I�N����[k:�6�Ę��.��R������c��}H�l`��kc��eiv

V�z�'2�!��Z��;Ĕ�Cx��ka���k��qMHk�{q��r蓟����lh�Pv�"�
NoN�Qf$.��W�w~�ц0�n厔�����QQ�Z���K��H�FŎ5D�^�;�$�qTD�)-��t,�,+-���kmom����?�Ne�1%��S4j�j���4���^8o)���t�ʰK9��Ո�1Q>.�����K|�	;��d�1\^@�bhǧ�:v}V弔D|��꺍��Yޣ�����n��"�Z�G��s�>ߢ��4�+�ݲ���L�/{c�58`@��
cu�^���Y<�Qy�I X��N�}��)�!���}<yM6<ʬ9l��9��
g����Su���ؔ��?�Qb��{ ���TN� �K~��D㛚��>���^��	���ɸ�� �2�і>�E�~�y�-�}@I�|�LBು迪'��o
:,���} uc9o�Ҕ$�`w�ڶ�����w������R���s����r`9��=�O��6��X�x~X$�������n�S��騜�A������Ӕ`����O�4�#�'fv -WG8�e���Q��|�>�����	y]Ц�dm����ٙ�䕎+vI�/<� ���ƍP>f�$�㆏��{�v=4`����/+6o��,�Hz�)-�#���F�j�ƨx?��-�:ٮB�Db!�����Be�R[P��0� ����C�� ��\_�jR ��RӤ�[Xc���j�j����Z��<���I���ȑ$�4͋DYjy�ԐF�١��f�{Z����	7�HuiO����Ȍ#�d����F�:ezCxSfd������{¬B���vS32-�������XU��vɿ�s���0N� y��[]����
e���5ӊ*d �ۓ?c9�옢b-31R]$���)\U�ƫ@8~C��4&�����l���tU��w��:��|p�)��v�9���w45l&�v���A�F$�5�4y�����,��7T֑�����J���&Ui+���r(�msRK!���Z�,\j�f�n֍�Eb 55]N�g�g�H�V[����>���ꮋ���G���c��
����bw���)�d��l7!��˩�����O�"1��E7�yÑ��/K�c�VC�Z9�=��b%����{������	>�"6����2�O���CBgW�Ϳ�M�"$>G+E�P�ӾT����W_�\�Ы(�)a|+9I�ĤԸ���^�u�� ٜ����U�IU�3�۳�/|�F�Lj+�l�4�(�����E8C��AZw����/���Bc�G�l�ظL�[;�k�q�s�7_�3mId@N$�@����Y�����Wmb�kŀ׍f�l�a����2������~�z�H??H�l�(ڶɕ:�;��֧2���28�����{�?�b�����@�XL�n�Y������y�x�Ӛ���+("�a�
�X&w�,SkS��������.Q��BmT����=�`/���3�DN��a�C��L��+>���)|/U3 �L/!*����M��K����"�bl�^0����	�5���|����\7��a M�w-��(��;��7� ߢ��#�`���?5�H�;Z����I2�"T������� o�ǖ�1xj�>��n�j�6l����Q�ۺ�e�;��qf���:�u�X[
6+��%�2���O��r�_m����&y�>WXg��@$���PR���T_Gyo���wտ�;m������-��٪�����I�K�{U+i䈞��b�/�c��/ے2C���]x<�v�+��S�/��������2��C�ʔ�)����\�����ue���o�)2W�smk�J���;z$� �7��UeQUjwc��G����%�Dŵn���3�v��-�?�e�w�����j}wվoϽ�ß��$���(��)��ty;�� ���C�*P��cԞ_(�u%F��#"%rW�����^1~�b��NA"] ��h����	;1��3@ (	����8AiRG�����֘�9r�`.XT�G�ςG�k P1������~�� �{
_O��Z��r:Y�l��+LD˸�ȋ�{7\�y1XU�.�a>�" �n���[c`��,F����� ����Vk�F>��V�{S��d�:�]�bqI�������Ovcը��&o���Ǟ:C"�l����Ε 
�I�,���h}�{�l*ͦ!�3/�ޯߔ~
xl�o��@�����Z�O�[��V�a��:nv���	��v�ځ�mgS/(�����d£9x``��׭��&�E�i�1 ���ܮq�9a�d�����k�y�˕�H�>��i���~[cF���΋M@�6ZQ�"*�:+Fp\WK�qV�V���q
J� L�C�����li*5��)�W��l��>�������ZBzs ���î��ә(����s����'%�g2:��ؗ�Jռ�_(�NS�yX��+�?֮VU�L1��
I�GYT�ț��I��e�-  y��� �p���:\������簼O��s��X���9b� L��++��>�$mB��4"�Ε�^ᾌ�� �YdW���O$Xh���D�L�p�^?n��}:���(�k�_T�T��ЫK�{��T�A:#���a�n�̛�'ʦ ��q��'S)xh�S-Qw��{�����@G����ur1O>_+�q#k�@;�n�����X�.�+o���00�P!N#��+�T�&b��L�^���)rZE��� ?'}U�z���T��S�S��f�M���B�4wҞ''�~e�	�+��r��׷2�-г	�_?���֡�hbb������%z�#��-�P��m��H���T����R�Iu��[��H�da���<���C��O���8����"� �T����Xc��?9�/A�Y�4a��+�u���,�J��=�ņlJcp���q;��>�H�z�'.� �Bv��=Is�L���äU��`�h ��N���l�DC��]
��tWu�>.�4!��覬/b���v\����V�T��0��,ŋ5���c����a��Vh*�b�'}���v��]��x��L����M�1��B[�Y��Q�=��Ff��ȃ�T Ȗ���{�iᄑ�]���[s}@��<��pE/ѼA�7Q���
:��d�����3��Q�xR��_�"��D��V�nǗ>ݮ�R�H�ǣW���ח��@1�7xP��d�'�#H �chW������t;���%T�++�|_�6�:�q�=�~���Gd�'�,�/��G����Sy���T!��20j����<(��(^�������@�9J3���q���k�E Y��T��-�^��	��%���\X���R�Z8+[��qY�0�c�����܉`��\cf����D8_\-r��	C�(��"c`�&��8f��2�/:~��l(U>2�ǾӊM��t�&���rR��ȓP)�R�� �/!�ˤg>^�7l�@ )�:9�0��cl������7��.oj[� ��dl�_%���Y,!�7�)TBE�,��֬�n�&m�:�m�����WӋ�<n/�H?�e>���M�<�s0���(L���)����k���d�����VF�U?��%T=�4P%�t����:�K���+�x(bE �ȸ��P-�J�(�8"��l���dU��������2K�\4�+�0����:9�5�<���.7��X{=���I�íW�}���C��<�����W��(�[|EM8El��D�NOs�Ur�����	zr ����C���(gf�~�*ަoX��g����&3fpP��j�j`ϊ綑%0��t��P�"AQ��x4�8}B���c�1z��C�U��]�A�~�kޝ����_���K{�U�� qP[�J^cKK�U��F1�����,��n��������4�.�O�`	��s!_[İK��.�l~�K9��a���L�f|�.e��(�Lt�bq��|���"��e?�T%И��#�n�����z�v��zm���E��P�rN��x+�&J�YȰ\��r�i�vj�!*$h����t"E6!��l��|-�t�vM������nF>���<!��5�6|��hf�C���-�aR���q�>k�8v����ǉ1�/��3�1E�i�4�����(�%�����'��f����S��p�S(\xy[�2kј��s�?rێ���u�v���C���y���3�W;�'555�������-r�4��\@շ�Џ��5fj/��m��-��'��R�P��g��+jz�(�1UD�N˚��tr`����=M�Z]6/]���ܾo�W�c��o�5��rj6�cv暤|��+w�e�MF||�!��+{�*ٔ^�z�����K&53;;{�FzQa!����a��y�z{��|G�f}I���5���O���^�Fۛa�S6Bo���.HB*���H��h��=�ƆCK�)2v����Z�G��q`z;�I�[�2j��(���Z�`��J������Z�$2i�'�D�x5?�j@����NU���]q��4���+������;��<�x(�	��2J�Re'��ʹp�92­+�Kg�������,�˳��Ӵ1Rɲ��9Ɍ����V��σ;�*��k�����w�i�X�S���y`E�럱��5�n� I6�>�SV��.r)�0hH��-D1��ex�*Up��?��CrZBm_����\HWyH�_��`���*�;�BѪ�8��1��MU��mi@���DH�6=`�;�m"���Ӆ4�y��ں+���n�����_t��B�"	��{h�x�����w�i&�Q ��Dr���2�H:�>n/Us�y��Ϧ[����o/꽞|�Vsb��&�<I]�P���	�ό(�O�+D7'�]��A��@��c$|/S"��ɵy��SfĿ^���X��"��.�H y�\à�.1�����8e�^[A��m�jTYld< p���k��2���
8��,���g�Q�o�� �h\H�h�����Pb�Hָ�?v  b���ttR\=o�ƽ�f~�@���_�F��o�_k��m�1X��B>D��&ODƳ -�o�?R��B����k�v�4�OJ��l)R��\+�{��n骦k�} _a�,�y�Vׁ���m�!��|I1�%Q��l�O�?�-y�!�U��$����X�I
N��X��<ɵ��}�lJ��%�~>��o�Z��`�o�g��H�ʖ'�tce��o.[�ʧ���Z�{���?)Q9v�sA�������E�7�A��sE��?������KB`n�c8ǅLͣD�M�-r3���bH(��i0u�i����I���]��t��=�j$d�	��[x�I��ZZ:N�^~�;t/Vr���ty�>������{2�B�\Ք&�P��:��k~�ޘp����N�Y�Ճ�����b��H`l�tݻ�-C�	M�$j���`�~}�TC��:}��b�\FTy���t��J�"��D��-|l��i���v��b鈟�UZ����o��?z���TQdK47	K�� ��_�7o�t��r$g���tx78�Z��S�A�Z8�c�C��� �mS`lc���p��G�k�Ώ�%A ܚm���pZ窷)�\��z��=b��S�
ɊG/������A��Ю�jó�_'����� eI�\>�����E��-,�𑑿&�����T§������_&����@�+�_�/�=�z���}.s���5�vv�e~�*�F��^�Дda�~�D뿊��V�'6~L=�N�51�yE��^}D������A�5.�/�P�Ԁ�R�]J���Ϊ��d چb��µ���YW"~�֛4	<s��ySM 3�Ѩ�*��Z���`TO�>BU�켛���U���B��D�� C���",A�Ӷ��G�RX���ޭ�I�z	�.�Rq��>�V�Xז9ow-m<�_v�"�&��PP�!AI��$�����������Q��]��ۃu�
�&DL�\�u-k�?�(����),2/w/�ĸ�Qa�޻�S�ی۟�\�v���žQM�<�U[.�g̲s:��O,�>��-U#���.X��]\�bL,=X�i�2Y|3J�nl�D�����۷�Ԋ�h�L��U�����B+/g}p<����M��<׍e1�����HDX&�n��(�!\�%홵�
Ɉ�hlNXTz+�:vXڪ�N�Z�-� �CV�B~F����U��������q!�U������i�3(����v�x5��~*�*<����9R���{�'O��vx`��@�F����$H�%����	R"�X'���}%*��Q?H�I���N��4��k�ce��P ��.�"E~��[[8U�0emw�݊TxCDϲs�m]���L�%���1wP$H-�=XfM��·���lFW'���R֗��'e��˶X�5M~��f�[#�m���C[CD�:����Ċ"��U�Z�B%���{���sV9HHC*O��A�I��)�/)6�-�e�^�
5ǿ����{���T��{Me�8����5<a �c/L��e@(��̢���Y�!�]��:��,��%,R J4��(*tl(���b���q�
�dX�ZE2u*�Z����w%O��R��
 ^�;��Z6/��G�Vƞ@�lP}���U.컮�vI�R����4X|ezk�%��V@� ۥ8�]�<RU_�-�
�9���?��rZ3�SdX�̈�4⯌�'?3cVm-t����N��R蛗�Z�O���s?_-���Dk]L֌�s���0�XB�a�����^ϻ>�}TN�*�L�Mk��X����o�=����!vηć�v(gS���t�A�㏣Kǳ���\�|{o���!q��5w_o��T���(��/�>_����j��S���zڼ���`���~b�號s�b��o̿�ʩqR�=���x0Cw���74�g�+��{�
 `�4�/䛙�`���}T;۷ݍ?<~׫�\h�?����@D�c�r�3�* y��̴�Ys�* �JT9��Ӽ�{�~�K/���Tl5�C�%<������˰���1���N9�m�]�נ3t�:>�Ч�Dv���J������^2(���yň�7/)�Ab��-����m�WO��:�}��GZݞ��;����@�\�wQ����#p��*�-��Uv�l��T��=L$M/�?:' kr\z6L�VBcG��;z���E�G�z�&_0�EqN�PE7�E-����	.�t�@X�Q��f0�oM�踗��v�C[ͣ
�~�;roX`4���(1�+Z[*q�?G����aݰEPG����rzoj�9�S�����8�p/����s�V���m�e!O��"%8fW��e`�j��	�� D��y���pMy���SWwqM�{���Y�����Q�F����x�Jy�6��w���_6��
�X.鹽ub}�t'H��V*pJ�Vj��S�:yЖ?�JK��nV������hDbh��@Ŵ���N����ќt���Ή���ẑ*�7e���p㵄��p`K?_\�+�`#^E��̫n��3@GSDl��B���үY�u��.uH.n��{Q`�4�LL�hO��(�ity6��.��Z��+� 8�,ҟ����ǒòCuۧ��w�L���.���5Z���~��s	��=��DR�c̈́�v�g��� ��f<������@`
L�ku��)�=��ŏ�&��kf�ymW��e���,N ج�R�1��2�&��݋C�_ϟp�7��	�O��e�z'��p3梤���c�u�c��s��T�����>%I���2[�o	|}�rx�~-q�OF�����V�ͪ�t�nn��L�0�;��_8�֋��s'�\[9��J>�%�Sa�+P���eY�o��⠍V�)_�ܡ{��p�_PU��n�y�HmPޯ�x�	�DTi��]Q 6t�����}�������u����OA��S�f���&�#������bk)���W_��H ˨i�dM�Ĵ��ůڐ�V@e�g�K�l:u�����
G�H���OI�[�t*�Ă'�1�h�4���8���`�Ea��ge�׎	P#ͳ�S�bBI��%9{��搴��D�J�pǟ��[��ڐ~�Y�{v6����@B/u|��ư��	@�A�U܈6;C�
������p����\��`#��4�BO�T��>v���-k��kМ>��I��ɇ��ש��N�00���f�Y�ȧm��[&�oo�
(r����5���p{ǈ,*�IP��+�.��^EbV�7�,�gkx��ĺ@QC	�$�g;�[���}wp�Zq�`A��wԺ�����+�X}I�1��SRS\��CB|Z��B9�:=yV΍5O�kz�����XZu����}
j�����v�z|P��� ��%�h������nXl#�$�mH��8�C!�̩��'f��PZgc;�?l�+�󉷟@�tZ�3�C����8?�=M�t�b�ܩ<�W���`�}� H�s��F���~�Nx�F�R��O���>����E�׹oq�h��+��ԗ��Wq e��˯�<zLݍ��n��G�Ƌ���f��>��T ��W�$��eC��볛5����V8��\~� m��Sjb��B��h �@X���]�%��؜�ܘ�DoH�z�ж権jANA�c'D�H���Km�$6���I�R;O��Ble	<�>����n/+�m#�v�d���4�,����F�U�񠮔�3��p��1^�4��d�'����oO
�T	���PMA�ߩ�}��o�7~��������*�����D>cL_�ѓV�t#��kKw�KZb��0<o2�'X |,-���p����� M����WO�4��(������6���C��k�~t)A��Q��<�����%[�Ӳr-�6U���3=���Ų�%�4o	���IUX��}gm_�Y�(�7%��dM~��j1��.)�~H���ŏ<&�:��&8�����
pq�n�J+F���w3�����#�Sb1r�%!����$;���N�iGm"4
�e	���m�e�#(y/J���X6�8�,����`2�Lzȗ���3>�*��`���D��9u��DEj��03�v��;#{e���ˡ���WU_?R��?��-]�����o_��&�p�q1ja3�Ik�靟uwo���
�Z�KN^<g�cF��ڣ�ՄEq�,���N�������J��������ZI��a:Ƌ������H�* '9�����dg���3���PK   T�(Us�7+5J  dK  /   images/6c71542d-16cb-4630-930f-71c4de5e1144.png4�4\�����G%�F���w� zｷ�e�D	QB�����+��=z������]ks������s�Q�*�xؔ� O^NJ��|��` �_Q3?� y)q���m>�Գ�LWm�5��G8�� ��0P�����h(_׎��hx���๓}��2�Y2���e�`e�e���Kw*�/��|b��G��,�\*k���-/X�F��fg��œr�z�cvvJFK�G/�/i�)m�b]��8�X
�LTjYx�*?>��98����O"2����.d+E]r���q��JW���5,�3E�G\w���_����� �Bĺ9���� !A���7�D�L�2`qx�^2b��z�-|�_�Q��o���O���|�w��o2r|u��؁�P,$,��~��v�7�5==�ʕ�����I���1�B'x��G��'�w��*��#N����G�vW�)�S�J�К�V�%�0�=^뽌�S�13�E�j�^Tj�i�xJ,_3��������T��ٞ�Rd#%*1]{<�+KSH�������`)\�}�^�X&.�.C�f"��#Dj@���a!�B��L ����ecŇ�X�\_@買Ox��-�C�����?����dʲ�J�qQ��s�JC�е9���tx,xXb60u	Ȳ�l�Lˢ�:�l
�Ð��ق��}ǿ��Yn�x�t�E^�M��x��-G���M��άG8�jε�:��C��#�,t�H�M�Q~O���Q�)��%#�!���2�cS�!)�����k�l&m��%�� X�)�t�琰X2�_�N��DE��W�������(�]����R��TI��F���Q��A	�
��)�)/L�<�٣�п��yR6��n)R���D'�-�G\
���FF�K�Ă@g0�/"��9�	�M�#'�9H�a�
B�X
w>KF�"	�|s��/iIġA���a>)5�:뿦���[:y"�B"����N���/$5vq!��}�Y$>��X�3�CF1�y��h9�T#���!� h��+����ގ\WggЙ^�E�-����]�ȂrO�Q�����#���:NSA�Q���|Y�,	�����Rj��[�W����vHpc�z/�4g<QZ�v����&�^�Vɭ���a#���(�|�D�<��MQ�KO�Ѝp�/ �l����Ѝ �d+��ྉG�O��Q��{��ڣ��u6\�@B@����0�g���㒒��QF��c��
MHBQO��3�V3�rP�� ����V��J$���fvf�����v�Y{�{~�Ű?�������E>�=d
�=hh����I���Ě��$�/����š�6�:k��D�0�U;��`�e��gV71"�qq���O�,�ظ������;َۖ�E#�3�=乚����ԭ9LZ?�˾nP�6��e=F@$���'�����`B1@���a��C��4	M(���g�1�Kq��t�-_��,����pV��7$��铂��u��)��eɌ����=���m�������II(8=33�Q~�˼F�~�/�g�K�PxPI��y�6n5[���i���X�O����ߑ'���'�à� �����3V �
��F$j�ö}&=�e(!��s��M���&8���(Rjal#Pi�4���O�>%�|�jm��7o�s۶|�-��w�}�7���aގ9��xh�r-�H�L����=<ʪ
@BD�j�C�r޾�5ȱNw�#[�S>Y�b�I��������V��[���|�b�����=_�kX�Á��FpI�����V-��-y��B����D����^L�4-�G*L����pz�1��
U{�^��6)#g_L��B��['�D�Li:�aAU��ɚ�I�I+@����ދ�4��ޑ�-��؎��M��L|A��"�É������ҧ��T���}*�#O֪�x���ٿZYZ�>�$�������~�<lc�w���]��TW�Z^N0�ZZ2�̇ȧ*�p����;Sc***:����hkk��^��?�%T[��;Ș�������k��g2*Q�����I�ʲ�I�H�(�D��mN����7���X�j����M������(���Qn4t��Q�����}���������@�?�̉������;��&�wڷ�����ɰ�I�m$���2*ʠ�:�Zh=�MX���e&���C��X7 �Kz�G���O#����６|���������m/?��l�"�
tIr���$=�е����_��m���C��^Ӷz6��+^���-G ���%�"O���_鱧%��ώ9��r�!����d�; I���|8˗�(���8���EF��׎W{>��Ńl2#֏{��^szdM�FD'1i��	j�V>�*)Y��yq1��8�	��?I�Qz�C$:��h?�􉅲�_vb/�� b?��m	8*�䍳-������@�{��z���ͪdԹ].��;{���X/V��_�*b8OP�(j������̱K�w܌t�Hjz�:�����Ҧ�5�m9���O��Z=,��X��\�����}�W)m�����CKPe�PS"�N��Jq?WgG�v��kt^E�} ̩����$�R�t_2��QRRv���!tZ[G'x�G���| � ����˥֝�ʳ/5���XP��R�/x(&�ݟ� ��xJͣٴ�[?n�|��ܪ������l�bZ���;o(�5tx�b�x3k��I�Q��U��c	GD'���!F"�Є ������}���8��BP����4f9e[w�o��@�l�&��E�1��p�˷�HQA�ֲP��S��P���n�"%R�Q��\ڐ	(��ۘy��3������Ue;�?�u��)�-p1w�s�Dh~�	���:��;J�VF,FR�}�B�.��Z�Q�g�9���O��!Mr5^Х*V�غq�}�g������d~�xA]����H��ː��w�Nf2 c����R��l����m��]���oyےV�:���i5��D9�1@IYy���X{��>ӹ*����D|��w��¾6}k]�5a߾PI>!�(��B�d�jg��/��P�U��\���l�!v-���1�~�{	C�����7�tp��ফ���T�|P��?�DL���QSS��8bBt嶫������~�������*��[�8]�Ă���$���[m'��4�:i��zP�$E�o�/�2&�������Х�'��:E��,�������l��H���g����=�*������3ܹ`J�`�5'���cD�rN�k`��[L�p��& �S�kV�g��� ]��^Xˠ�;�#��G����4;<��ߗ. ���\ 4W�	����2K�n��vd�L.��x�����e1lC�~	vjЦe'A>s�����%��X������	�+�`������S�8q�Ý~�tgc�܎묎�������[��?����OMu`���3�tߑ��v��۷M����}*�3��Z����K��n��9��d1��>6a����\���YZb�Y�閙�%�2��td*���%��p鈈Q/�����R�_j�HQ��%����k�`�Xo'�VͶ�Gn�;:�+kD�<=�̬�`Lj*���&➞~���lUW� ����4��������*�2����m�������vH��"
��UI!e�N�<"ȇوHq�^��UduW+}/	yo�C.A ��ل(AS�
���+���h���J���}�vCF�!ԓ�H�a�ޤ�;����HRS�уC7���rMC��a@F�,��@urzH��Z/�Ns�gK\ۇ˵�.v����/�4 n�pr&&��DP<�<�
�e���5FO���3UТW��U�~�m��� m`*������z�eˣ�g�>�GF�1	w����o���smJ�M��"�?o�u&T��2&�OؘT~_�=�>s�Lo��K)�<��{ӱk�baB ��TC{���o�B@}�ıi���@�FEa��Q V��ؓ��f`�G'&�LMQ�HOO���`���.�é����F͹�F���F)ju_6��4,P�<!A�e�2���m�Ȼq����4e�����%	MM �� �&�Qr�G:�ذژD�K��@G�ϝ�R�u�+@�#�i��b���Kf�f��M��[����=���q.Ȭ��z�y���9tU�d\ò��pi�xAj��-@�'ڟ'f�	������g#m>���J(�P�:��� '�p�bJ��$�9��v���I�(�����ųv�w�^w�77��1�(��Ǉ�������ՋY#r�J^� �����B*cTlB���
����7n����_�?�;oOM�
|8�ո�������BWM'2�bآ�l�C���+Ε���|�����H ؎������X;ݷx�.L���S.@-V{"L��!���+�ao愯i̹(ҋ����F���!T��z���<�l\U��?�� &	����7s�	�'[[[+�(�N���Kآ(9ݣ5n�|�����ݍ�F�o4nXё�̩�JJ�6�pL�I)����-﹠o���ѿ�ҋР�]w���]�oxx���΅b��w�Q��\`��5^�lu;�m�]��nr�������|g#u5���J�|��*7�\^�4	������ Ȳ��_�)��lO$�=�>��3�q$����������9��ZT�Z������^h�?�pV ��uϝc9f�铀IA�#�� �<J"_��"V�L{Է�o��6"t�A'z�#�}}j�Y4�&���,����Ö�Z�rLB�t�;��r�m��� ��4d�����>i ^d�{�}���H��!]E�Y���]�499���x���g�2�����H� t
y�f ������:��Z��3%"
�L�����>i�>�T����������5������I�����������T�Rl�i� �N���W�0 :�jjL [z�&! �Wt<�ӊ��M8�"m$����g}�@�d��N�?�:�	�2��p�~3�=K!�S4?����giee����wfQ޼u�Vi���l�3�Q^'�X�r��PN���F�ÁE՜�z��@h����v\ta�:��RaȐ�V��Ac���*�'��q�l�d���l����2�*�����}���J����(���dA�镑L�F��-u��	OX����,���ud%#�x
��s+b-'�tr7S)�O%V@i��,�3a�;�ĺ�S�����rCRGa�klW���$�5~|wY��o���}}��y8wI���P��e���;��o�,�7K�Z:n��D�UZ�Q�ܾ�|*7��1k ���@z�6 �'I���a�3��ˁ�p�0���56���|��	�G��f|�Ώ�3�;���s��}1*�sZ�䦘����rJ����F%��960|Ռ!�.��� \J�wv	��Gq�=B��ڕ��$i%+��#�����N�dR$
���JJ$��g]�?z����)o�����u�ou(&�u�����t��^(M�:���gֶ#��
dW��Cǃ�b��z&�������l���&i�����dɎ2��MQ��//XT�p�7�2�Ka�Q��4_���hblPmCCC����9e���t7��G ������A���;OЋW���X#ڎi�ǧ�J,��_?�V�<�D|�'�����v�x������/��� ��9����B�Gd��O�C��^���İÓ�k./��M<�8��w��yPp��`.��A;]�������dnY�fk�Z���-�tŭ�߻zX���j0;5;;�ے���vʺ�^��Zߘ�Y�e��b�b[���6���;�u�j||���3pq2h���<7%�Z,����籝����~��R�p��(txyŔ��C�j$j(����Q�t���Na�?�|NM���5_��U*:X��@�c�#7����{	�H5��T��������:i�M�����%{<ʒ\RU�a{�0jj)�,�*�^`�^�b�S�	������W�>�P������n���o�?�;5����G��l_�m�[���2��iii9Jf��])�ÈH{�S|ŵL"^�vtKZ����ﾱ�,?z#��揞�V xŗT�Sm1��r�+E���B��I�E�/�[�����.%���QLw����V��g�{�-�>�k ����=���;��^�cit3Ӽv=:j7�[���q��MVK��Q�I����*ݶU�w ��H�G��4�^K�Y �0�]��8J�z�kɪ)��6j�N�Rl�6�5��y曫Uf׿v�L���x6:4��Q��~������P}����Co��<�6~Jg���ĒF���/�?v����|U(K�����2"bʑ׻���cJ<�0!���fl|�+�I?��\rc��?*Fb��q�i8�iY:������q4ug��c �ɛ��g��PSQ���ճ�j������.1*.:J3���H��.�����%S�[�O��p��i�f�U���l\�������� ��p/p��6tHי�+��!F��9hu����x@G�T��ళw�5�� P(]��0�����6_x��XʞN�\V�:aX��|il��3�<}�ҨOyO�ak(K�`6:l�GZR�G3��(`���'q~�/ϰ,X�����n��Z�m��-�F�Cf'��i	��Q���g�����Z��PYM:������o�
a!���Xt%Ҍ�Y�R|
� � \�����D�_� �8�j�N��jt�迟M(!��S���cn�x��T��Y�V[3�[bƗ��R���^&~~����.���n�.��&���Y��ZM�e�q[�&gb�p_�z���{:��l�K�I�g�x_K�?w���4CÈ9LW�غx]��B-t��ז4�)��g��  T�II�@1sX�?�To���Կ�2���cOլ��$��U�&��e=v�5�K>;7H���~*�j��p᪴,n�o� ���w}:��YD(����J��Ƌu��l�*=�lښ�1q��&"��@B�͋�J�2{A KC w���U9�,9�X�$�����,���!���Ð�ȵ;�]��`O#�$�	\��oJ�	Uy����N��G��.�f�P6�GFy%4=>��_ez������E�m��K�KV�d�MnV������E���Ӎ��
��3�]w�:�g��d�Fv���7�d�+A��OfC�DD�z����ĸ� �`�xj�B��v�����H �O�BAv�zd1J�[�Ĉ�0�]�l�~���3F�0�H1��Ԯ���W{v��d�T�
�V�$#�M,,��d��(����lwƐ�*���Z#��������y�4�rؗg�ۣ~u:�۳�y�m]��2�`�z_��Ȃ��r�ni�����7J�Z�t���}����q���#~�z�:V�ʦ+�����3����
j@�c�t�r�o߾537��� R��'Q�Q��?��dLT
�opJV)rY��t����=�K�;ep4_¢C	rz�\���}e����1=u����V�����x͍�<�0j�:HH�D^�BaHj*�����A�r���7:���߶�$7�g��������=�=Ze�:Sy�j���h�s�(9hΣL�gJ��ͣ�K@��K�i���+���IBUm-0� I�<�Uʟ/�~Y�f���c0+�m}�ݵ��h���r��� �bQ���P�`h����&�72�_�6V�~��J�Z.#L������b!	Ck��?��7���T�Cub��ag���<>����Β�_�ڋ�|j;Q%��Q��lN/q��4S�^��������^ ���Z�^�|�H���䐇����	��@���8�����O�@��\1��_�֏7�q�p{�PH7�'����͍�Y�n�l��LF�����+���3�G6���c���#/�(0[���t���nZՊ.�՞@�Ej�Ɔ9	�5=@� p][+[cY>��B3�]����$!Ќ�h10m�1�T�c�OY�@A}�-1������^{+���|�j	���N��w����Qm��{�M��<��c�w�G�����������yCG��J+1%Xv�L�N�6p�����H�����>j��l��I�2P�_l!�G�zz�9u\��������)�r��`K@֪�+T_�$������#H=H��%C666�����*�ХeP�D	�xW��V�f��� }���ng�Y�Dic�8����� $M�x� ������ɂ�{�?�{�M����t�&'U�c:����JS�q�^�O�,x�#��
���h�������C���%�WX�6���{���s�Y�Θ쌊��:i.�ä������NJ$�HtX����q�*��>�NI�����6VH&1d���PRr�CrT�&��U�?5e��D�~#�|lm_�i݊�Z��x�A4�RU6�L��PLe�=M2Е�6]߀:W%e_5���ȼH�L����V�`+�:h�@�ϙ�vZ8�kk�Gal#��D�������.�?�?���� ��gӟ�����
�t�9��_�%1������9kʐ��ߞ��Bm��B����0P@H2�|�,��i��[�?o/�H���P����:��Th_�E*��H��:Gw��������l�
�fl/�c�����W>��~]�v�ӳ��>ߌ�
{���[q�~l�I�՛p�Շ�k�Bov�JP���4� Bh�;MO����������c�($����{D��������oo>���:�����#�1a��r�����M��G���8��`΁�U~|́�lp��)�q?C�cbf�jm-�r�IR5�����u�ad�1%xU���;���>< ���װ�)x�viG�5�P��ȗ��c�S�q����\�t_�_\���9v�9���$��	�7:��?�,�
ݖɍ;��UJF�Nu�](��-��'7{f�ֈ*�uI���yŤ`�c�/]@d�ԭ��[�h(
�ޖ`��`;�Mz�������xL�>z�ߎЭ0Hh>4��~7�qZ
	F������dx����Bm�ea�j��f�#��)�sU�?諔$u�H���py�b��
�ߧ� H���4R�a7�13$�(s���φ<g�;���Ҝi��@��F�·�'G2�K�Ee�aL�Vԫ��q�� 4���e$��ϴz�s?ap��!�&�ρ{�o%*ɗ�ڭ��qli�? 4�}�*�������[#in�9�D��)���n��li�{{0Zځ��s�֋_z��&�	ӟ�Hݲ�*��F��U���0}'�%%W[�y|��gKf�9G�Ht6P��`��{g�z���&75�8�.�H%e5hn�r�f���f�3i(���E�T�BW��#l����?4^�5��l���B��p��n1H<<����p 4���v�"w#0���4�7{>�1{�j���cs'��I�~��*�F�,m�А�Cԙ��u�Xp�C��
���jʓ����T��6xs�X� g�� О�4����X;oP����u~s���`ݲ����^�Y�c��@�y!���GP^�\rXF��B�+C0Ȝ[�)j�|�q/�ە'�%A o���I�g��Y��VU˴�`�%��%.��0ժl2h��P�R����ro�Qo&n�_+�}������U��G~�,����kzv��ȡL�?Ǡ���7�T�v�N�/�����&��j��p�Y�k/�7{�;�R�T�Y�rA��r�pp�Io:Ͼ2:�w���hm���A�BZͻ��a�Y���^_Ћ<-i��]���s{(س`Jn��P�B��~d�[i�Z��P���˞ж���q1���g�c��*gXQ��X�gϤ�2b� ���8�<B^Zp�iQ���4	N�|�5b�2Ijel�W��P҄����3a�hfP�NL�;��{�n"��f�ΤB-PE��V�ދ
��y�X-Y�l���ڎz�]N�7<���v�n�ta�ڃ�5���M+����&\i^,S� ч��`��C�Op����V�b|��7nXuL_���d���;���������_
�}`#������<OH��0�$�u|��$�Ўc��� <`��h��,�is�5��q�#����?��Gm䊊��F���W:Q�^�:[�`B�J�Vw�f�I�ƛJ̋�<W�ͤ�6e�{����{cƸQ��2��|�G��]����h��síp�DsD���ؾ�nw�՞����NZbؖHZ�v�W7&ڙ;wB˴-Tv�8�m�u���-VL&o�g=�":��+Z�
Y��$Q���cF���`=,�$��:_���(;C��%�6Y��B��%-�k�=z�}���~�%̹F�/6� �Z�d�ɬ\��?)O�����A&>u翃�����~D��>��Aƺu~�����ľ�6��e~���v�qJ�r�L�
҂Q؍�G3��`���ц���iK�|K�����w�����_�-��r�v=4��~Ŕg�1C�\j*�|=ެ���~�aB@�q�:�w�!�p��u�����Z1I�0��|q8T*�y!T�>n"��l���Uѷo.�c=F(�s�-�L�[�x����)L5e*��l"A��j���t�QE��ԑ��,�LQ�Ӆ����풆��w�6pn�_���!#"�.y��i�i���Fe/��,L��)�����Zef�a��M��?��$��.�?�p(p8�ej�=�V�t+��+�f�+ �����"�u�`�yM~�/[{��٢�]�^#��6�{�w����c��0JJ	�������qn��.���@}p�L�AV��O�g��4*�Ǿ*�� )9�G[?S���
c��ޯ1�ӨW&{��Z)�D(gH(1r|�(�^�<�����v*��4��j��i�F���\(����t�5��վj���$#�ԋs���@��&��������ٳ$�`N�%�`.Q
�d�VT������/�*�:��-�vۙ��K�f�X�/Gт���d����	 ��glI���uܯ��t���$�����X���r��,����L�4��u3g�kx���Y���57�{%O���@ӵ�W/&�(~���xv{���5<��PH�ۣ���GWA��C�8Ge�k�\C�̂&��v.��L����r�t�*�9<��3T��L��>{)"r	��$((�V9���~�z�P6�|D��菣��/P�12�Hb��T��s;3
�)�Wy]�G*��ٲz�&V��){^��z��g��t��sI��ή��I��V��-29��HN�6Ûq�(,�A���M��)JJր�Z#�H�9ߜ�}�n�IM��y�wc���[���/mWݯ����I����޴���y�vQqN_(i��Z��Y��]�����ۚ�G�D�\f L?Wv&��ɷ!��浉CEƵlW����/��B�:a\��}��D���|S7��0oO�����������B��7���h����V@�xp�;;�Vnۭ3�,--�	�$��:�ٞ�(�ѣ���~q�@�����~��(7�Ǧ?�T��� L�͎%����&;J�F!+�2%��e���LCs��gf�(�a��t�v�^Vgh�����9�MO�:����Pi£��q�m扖�ǳ�ǡ�����S_7�)��l��&r���"z���͆1��de��'5�2������.k�7~�@~7�t����j+5w�x��ߢ��O�lj��!��:eyڧ�7vN&9�ޛ���R����(`q(����D�M��aTk<uT�@�H��U��N�g'[F{@ª.Y���?��QO�Ƭn��gu��3a��r
Ғz�UVB�@��jo�$�l�����#:q,ܡ��+1IM�T��w��sQ�WY�����"䉖��gϤ���ذ�D@q�)�R��)>x�oK��"7$�tR�g㌽�*9�T�̥�����3�����=Ѣ���%K�__J�Go[ۛ���ѻ����N����;濩��sx��U�q�u����o d�d��֦�گ�M�G}eZiBJ�`v�W�*L�|8��\��⨵�������"==]�|���y������"��V�a��_���<��>~{�z%���]�:��%�����}�R�㝂���G�5�������U˴�v��>}J��s~��q����*����[N8����������G������5�ט�����*��š�����_E6��*S֝��8u~�G���#�3�P�y��p5��Ap�8��?Y���
��������z~�2#�"yE�{S}��2�{K�ǲ�������>U�����C�t�D����-a����Ɍ�-�/_>�=L��X-#�ksg���|T�k;L#�ʶ��`����E+2��tt�DO�����(�o
��a}_~�[M�	]��a~" #(��9�s!lޓN��ܝȲ%η-��a撓g2�@���{A4	JP0��r�d�YTՍ�/�����Wd,�o�v��Vzmc#�
�|�츛]П��:����WÏq�7UTx�K�S��?����S��$�I
��@A��h �\Π�!�����?���t�!�A70j���a�w�� ���=�<5�=ts�%Z�ps�wy����F���Z�N�
�^=?�Ӟ��y��m�����Q�iHA�r�<o�q,���7KsZ7&D`5�#]0չ��X;�_X��>��!�TzЋO#O{���d�{�C<w7�1�{*aK;����
�V2p-GY�s~ε��|�f�5Ϙe���=~���&P�ǜ�?�We6�!,W?/C�T�b]�C�h�%*B����-�O}7(#N�i�։�;=�R�ť��hAƀ�J�8����)���4�J�e;�R>�q��?6��)���ӥU0?���,%���O�e)C�.�fE� 4AD���5%�`0�`�=H��P�4F�jҏW���#<??�g��k��1���n"@3O�\3���TPv�hh�7G�2�.��Y�E�`"W�Ö#�'�װ�I�<� ���#?L��5Y�?r��T���u�җ{{�FPi0O�C4fD���ׯ�֟���2/pE�Zu�	-*'��?�
2�VJ߶3��WDA0�U�K5:����c��\���/>��=�a���P�p�)�o?��Xr8>���"Ab��ƾ�_��k��KɃ����N}��o�lm�o=s�`�,���-����L�Z�`��_���Iy��^z÷|9=f9}���8ս�!���a�Z�E&o�7��T�d�W����I������!+8���u
2��?����< VW�g�)��T	��v�פzm��!@U����o��-/@�+��4by��?%<����r��,��N4��jn������P�����~�oi��OA��{����k�k���g$�6�ms���R�#-�I�UZ��۞��=�Lh�B���m��yO=--�3�9�ޡ�Z�c��v��F�=�Y����K	����KBT�y�Ĭi.	D���0ϖqAǭ�g�2~':R�?���T7-�I��D�g	�	�~����m+�W�"�mmvgA���q�6$�Dr��ZA�lj?fE�<�_.	^���u<������
����z�e�Z@�+�mD��#��!u4��`�⒄L��뷁7���7<�,V&����쾇�[N>����l�~�+�urt���U�{�$t��:�ʒ�%�����ր����Jn��`ϰ�e6��w�~�.��pcm�a(���&�t^�_X�0Q��J2�R,f���+M��a��<b0��6wnp�z!ꈣ$#8�]�S��"���8��R���V��!�\�e;??jѻ㡷��=B��I��g�)L�����lYu�ė�Q����C�/!��ȡ��UHŒ�S�WJe�,����:2|Y�-, ����`����^��̞���c<
,�?
�D���g�^�^���w>��T��Oq�9�A���GK&5�i1����-�)��1���� ?w��� ��O�Yjh�0��#Tbej'�ݡ�'��;�|}�uR�l0����dxӵv,Xeraa9��L_�-V�;��m���jIɛ&w;D�/|��q�0�}����P ���[	�7�"W�F�k�-�7�FyW�ΎA.�Bl��ޚ-9P>����H(<�&spӵ��'�bϖ8s���#O�Ќ��Nq�[��O�hW�V"��]�p�p��N:NBd�5�e8���\t���gS�;ю�i�������Be�\��^����=�
�F?�!�9�ۦ�IھO��x!=����d�����M���k.���/q(l(u�hɊ��:'#a��㫎IOt�M��^|lllX��Y�5����Q:x�I?7�d�&����x�/���ux��U��u���\��҇#���qq8�Ӗ��e���G�k��˥��8'*zR�뇒c��}�/��y{��������&Ϲ;�
��y��.�\"�E��7��Kf�й4����2&+0C/�2~���єPB �H�H3����(g��U�![�c�[��M�d��(Zn��s�®�`��q�.�z�N"��&�v��/#
t�rU+�^K]F�o@b���M$���	Y㬀q�\^�N+���\��S+��_7l��`wWg�)�9�+�\f�I?͢�G�=�t�v�dB$���������\777�6s��>-
" �T�5r��}��m���U�������_O�w�5j�英��*�{��i�q�#t��F����8����Mb�I�Yȧz}��K��ѸNO�@-���j�̓M{+z�҅y�a%��Rd�ɤS"O5��t0Q{>(�d?wy����V�Mi��2�C�Ɋ�������v<��J�w�5,E������`��Sw�IF8<�z����`�(0͇}Χ�sf�ϝ�5V��"F��e���F���J�Σ�UJ�@�� �'�$,���[�����Vx��w�=�9	�[�c���CT~/ũ�1���5�3�0%�P���:J(�w{��&j�"��v�����#�L$0R���u���Ojld.��^�Ε���O��&��TU��z�����'�:ϝ����d�o�|�G%��D bV��*������1SOϴ~N��n�p�������-�,[�Jw�6���a��?֯�ă���ɠHp���+2S�XV<$y������FRD���	s��!�HS�"����Ic��<[��ju_Ҽ�b,�m��l��$�W�gk-��S����p����VT�΅ﳧ��ۣM͓��	׫��<I~�Ӎ�z�������Ht��4;7�Tx�S�Œ��3@��.��i����@a``��������-"Ǐ��$�	XS��S�B�߿,֙�TD����,�xTTT���,߳?���������'@ŧ�|�
g�)ڊ"fn�e>�+U�@����Zt���i�	���
��2�>�Z��,�[c5��~����(/����[�6�kƑ�(��2 �����P�5�{���4�����.�XZp��$�Bb!��&E��y��A�1ɗ����1�s>���y+r=�M����O�c�(�F\�P����5vi)���?W���]:5#�_�������d{��@q�#y��J�N��gg��g�EN[l:M�MF�l��ޠ���g/�l���=3gyJ�П2M��`����1X3��6���d�g~�'�,Z��`D"�O��-��J
�5�3�O-�Y�!~�0%��S*�[��o9��O�9��Z����#OO<u|�S�ɨ^L���P���	d��e��Y'1��������XV���IC�m�\�m$�O���SK�!���=!h����i��;'Ȭ��,�=���A` ]����ܡ�s�+d/fޟ�V8��3T��(Z#A��F2ɕ�}��LP��)���jϾ3y��EA4�ÿ!�I|~��}�rX��V4�=��=1Z�>خ�?|��f�f�.��m������Ӏ@�N�.�M7��xAZH56qJ�e��a��MNid�lw~	u�����`�����T5���л��k�И�������_�6< ��p�)�����N{?\o�p�C����� (�o�ě�)I���Qr?V��d1�)kO�qC�>D򥢽]�:`�^�*Xt\'7�2{4r{I�����_[÷�o�#)�#�Rc��!��sl]�Ti�1��_�҄���P�����)����n�sc�|SU����������ܗ�4�	�t�=��"1���m��)�	���l��Q���F?��Fkw���O��O.��pqN�G[O�gm͔���KҪ���Hvσ����Z�Oϩͧ�p~U��_���{��J�Jq2d��~�6��p��@�*���F7�iQ�`ۭA��8[�� r�#Mg4H��@��XѶ>&��>��(�S�ߣ�!(�ku!|��.��k���?�jQ�(�sE��\�]�ׁH��������c("Z���G�G�:q����C��v�����0'p�3kR�LmQy)�u�&}RU�h��)��;X��;2��� �SQa�p�I��l��x���Ã��k��QMM��k�_嶭���r�J>9@�bs�#����n�8��3�xZ���_�>=�����C��Y@���o�\�Ve�X���w65E���}�g@��� K���^�r�\�ZJC~z�O�� -DϞ5@H��K��D�l��\�zX1���&��CG����ƠT��y�޽����{�{���˘������''���>��f������jW�^E�^��˨V�q���,�l�ZM�y��XZZ���
*�
j���c���ݣ(�ds�ztt4�����7��f7X�B�=��h��]k�eo�M��,K��Ǐ���L�|]��0133�ջZ��̙3سgfff��".��ٳ�/i�F%ۇ9SƵk�2���O��(�3g�qN�N�s�ضoߎ��%,,,�ҥK�w�����T*���֭[�s�N�B�lf����)h�q���4C���ܹ�z��z����E\�x̌������:-�8���(�Y}�"�=�!2ײt���2�og(�� ���Y?~�����_<|��J}��F�W�+�2����f�����>f���oI��i!��9�{���"�ipY���������	���s�d��!8���&�A�)~�3/��h��-�f�N,�P�a^3�܀��̏�N]���o�4�}.K�Y�׳��Տ�U��\��n�u>͠2��777�����>������ݻ�W�7C%$I�Y���H!��I��_��������D�·�p}��#_k�~}&��F^����}������m�=�&02�M/x�e��~ԹW���g~�}�/���o��C��D����+��P*M���{��O���i��1��Z�}���ر����������7�[�g�f�9��zx����^�7�ٸ�|w-�� v�����a����Z�M� 6���޿�9ڊ���1���7l��봙~l��4y_�A��ߑ$�����v��ѭr���)���
?��t���?��?�g�<p������o����A��`@�����GSSS۝��)��3�^��0��g�~1�X,n�i}��$x���c�Q������ǯ������2�ES�ibb��U9�@�ݻ�������(S�����Mp�����H�ػD� &"-"Ph�) �Ҹ J�G2�̬ P��-DQ��0H.����:"��RA=�S։�	@���,B*�[f ���v8�Ի��>�vu�F��o���G��ז1�ވ=  |��NXk�*��
�P�I�:�����6#	H� l"�Oi#%Z燄J 3�Ŧ�[!!2V�b�P��Dƈ� B��rf�B�H$![�u��"Rld)�I����zL*�xJ��k���� ���$Pd{�'�Y$��rb��Ɛ1�����K��r�M��dD�0��T��0�a���lL1SpZ/"!bÜ:�ot:SF�<3�|~�K2ݸ[&+6̅_�7:_��^@m")��(�b���2q��`��Doa@K7�d�D4��N&(0C��@��C)��� h�:M�� TJYf�"�Ř6�z$��Dj���B)Cƒe"%�F: e���5�%	��DZ�\E=P�̖�%
z�w�Ek��~�7zI��0zcPD��zgV�:��ט���F�D�fٲm��S[}|���A׉�E��-=���D��d`ź<�@�!�Y1�LzM�"C"J������Y+L$���T�e�$}�D �DqZj#
 �E� J"���A
�b�2E�$ʊ�$�6&k��E�Jk#�Z�Z��*�tq��Y�~E�;���- DQ�,IL�Y$
�c-u���֚����2i����DDʥ�}"
ED($bf H�a��	��Jqgnn��(������9kmh�i��(��ur B�#;:��8���~%t���8ON�(ȋ�    IEND�B`�PK   T�(U��4�� ̻ /   images/7a4be1c8-201b-41f2-b584-263fc50cb409.png 5@ʿ�PNG

   IHDR   �  �   �6.u    IDATxԽ	��Yu�yߚ�r�}����EBb��@		a-�ݞp8��ɡ����glI���'&R��l-F��Q�#�-4��@�M�U�յt-�������~羛�*��7�{��������{��U���}�{_�ԩ����l���4��T=�z�z�V6�fsPI픪�ڨ[�������aj8��<�%C�WYH3��L�9SMG�Ri���f�ުժ3�zs��g+��\�R��&T��ڨҪ���L�Q��Ҩ1���a�T*�7G�Q��^�Z���n%U:ص+5��Qg0u+�v��ەJ�=�>Vz�٫T��`���y&�Ľ?$�Rܫ��`��m�'��*�ʨګ�NoП��*un�~��6�Z���I����Q���0<��})�>}Gejj�z�ʕ��kk�pd�[��[��"��ߵi��Zo�H���N��hX�u��hTvW��.*k��h4����a�oڍ���^T���zke0Z�k�cm���T�w�	t7R�V�T봎z�Z�J���H\���{j �:	ԁE�{��F�{��FN^�Zu�- Vp�Tj5~�|���i��e%p��>>T� �c@�C�*�A�WG�����bP���j�_��{iX�`���~j����x��F��VG�iuu��߹\o�n7���Lw�Ύ��̵F��Ơ=Gc�i�����Jsz�`�U����������Dk�����&g�;v�15�ЀKכ�j���T�����!\[3��i¦������;���t��5V�&��B�2=��15�NM���O�����Tu�h�R�sWj��s�zcNn^�sÁ��)8��mro�a�Z�Vk�Üis�e2�'A@7������N�3��6 �z��[�s����V�z���\�]�f��>~�� s�w�)���uoЫ�S�s2�Z���_c��;����*�Fs؀C4F�zc�6��k4�!�i8Z�v��n�Ќ6���:�X;;Zi_|��}�����/��������XJ�45��ިV���6�٬�F�S�6��f���J�V�;J�]0��h��''����si�֬��>M��Z 3��p��� 5"H��J��̠ޘ�WG3��`��]��<U�զ)�F�:l�氚�Z�GM��`��f��U�pjĔQ{�@=ti�~��&U���`ځ+p�8�
��az͙FO�4K�WKM䓪eҲaeU >I�`�4��z�FY������3�Ju�?\�W{��G��M�f��X{��\��{��'kS��a3��ҠI�6���u�oZ|e���C�����-X�l/[�/Oķ��]S������
�.%ޛ{��Φ�\eX�g#6�A�ҨUa��ҥ�+ w������B�A}Dk�fm4���0�y�c�E�* u�l�0�Z���@�� RL�)��-��n]k�괓J�E�W��C*��_�$�V�V�aT�����h!�9�$�6�j��v��?��� w���?E���fZ�p-�!{y�p��L<��1lT���R��9����r�M�
ʫ�`�HC4�Z����v�ta����w�oH���kmG�ѩv���Yo�#�]IW6��a����� ���F��N6��c��7���ԧfG�ֹ���9+)�흭�;k��;����1�r�G0!8%�Ym4�*���pVEXE �OQ�C���R�	����+��lTk��<��p�f��:,X+��&�n��"������4�w��ۂ`�$�x�^��ʆ�+u80����hyv�mD��0����E�H��/#x�� ;�7��K`�J��^!���br�0��Z�F2�]��z�D�a���0�&[�j����Y$}�[g�MB�K��A/���ty����W�6��W*��0:�����t���:HD34�3���>��O=�p�Ȯ�S�.Y�/��o�#oj�Sn���ߓ�t��P�5��O��޵�C�����J�Ԫ�Ȁ�^���ht��F6�:��4C��e�V��kC�^���:��5��� v������C�3Ih&�;̵�-�A����3Pl	�dɽ�l��M�#�qv7���,��[p��F���r��M��i9�v�E�66�m�#��6Z[[c�Є[2r�;v��]$�t8x�	��
��{�n��h<0^x>͂��0��0�?�Dk���]���Ӡ�{���)�huuuH�Ku�4��~���_�W����'N�Ξ9��c��d��h���2X�IYIk��N�CSb��t����T�I/q�#z��Cw��������_��h��[����la_��;�w�{ߑ�f�A��H���F���:���BlTj �-D�d����RZԨ�F��Ezպ�u�0?P
���f�������.�F��0?j9�J����O�q��Y_�N����ⱚ�:[�;x`v�_�V����0a�ܪ�
H���"+�wSkz:-..�;�#=�� �3V�NT��Fء��I�
�l���1ۆ��W���󎷱?z-����\�k&�����M9 �i��4�X�t��yԅ�M'�5-��6A�477�P#%M��fg[�����]�y��{������p�����7�'����y����f^��[�\<�䯮�;��~�k�O�c�*�s�����X�ô���ܫ;�0�:��۽����qe���X߻w����u��ý{�,>�ܩ����Sw���tfgg�Tp nzj�t{��
7��y�|V�m��F7R��NK�.�Y*k߾}���<� ,*�
�E�"�2�-��faa!���H�A���#�͇\T?�	��r3�*�,4�4��߈�m����І��v�꣙���ph�(à�h�C���7a�1�MY5��u�2� И�������joТ��p������?���Ni��S��m����4]z�4��/_�۰\�4ݬ��w��;��~�׹��gy�	}�������������g����y2�DI��C(+ree%
.����ݯ���}��}�.��f��l���F+k��s(#F0��z����~��=l�رX������,њ�� Y]^Z��߮=�cCr�$ph���6�/--%�.)��f�޽�g�}�fc9x�`ZƟ�p�����ܹsq|�����ŋ^���#G���gϦ={�G��#�M_@{� ��`�]����?���E�f2�tg����>�9#��"�W��vف�-!@��>����"�!:�4^�9Q!�� `HtY�Akz�7M��puZ��ܵ{7��;}����Ϳ�7G?�����t����.S�Fp9�y���0=������>���?����_Fpg`������O?�K���-�kQ8���۲���;�����kp�����9x��={`���3���,�އ~���t(/�o�!�v
Q�"v�ڕ�}�8�ٝ�h����r����4����4`��.����>Ŕ�v6�1�n�׿>=�����o��?w�y*���g�`�xꩧ��wޖ��Xg �ћnJ�^8i7����G�&���ao��栃�V�p��=�W���m� "~|�{�d񮝽�ϲ 7{�tן�0� �\��]��s���}x�]w���;���ѣG;$Q=q��G}t������8��8�����z�M�"�����{ϮԚk}������G��ۯ{]j�^��t�/#�S���z����>�K�.^��馣�Kt�s��j�B=�ēi߁}�[^�����鏮v��ӳ��gN������ޥK�y�w>��cvu�#�IX��r-�V��-�/�|��b��EZi�� 2[���r�95d�L�Yw9�~��J�cCAU������`�28d�-h�X�i^�
�uX��KD�cںf�e*�����z��nܦU@�[.7j�5���6��6��_���Rb��VQ�[nI;w�L�N���߾���<�dT��T?�هv��Ϭf��ި�"�ow������;����=����w_�=\�e����8����깳ggn>zs�Knm%�$h� ·��=��p������1MG�j/_�����n��w r��4	f�&��Hʝ�V���݊ ��qX1���8���V��Vhe�^��[��_��&�h��n(�#���� �n���̣q	�*
���U@l:��4��~,���hܥ���_��w�w�툳 �{y.`6-�ҿv��(6#?>��2/���������7�����������y��O|p�"�yl���B�sp��'Ϟ��sϜ�@$x�?/��{�{~�g���O������瞋nފ��������������nk���c��_������ߊl��y��(�Ĳ�#єQm�)Ǫ&���-�ӿ����b|֘�@ׯ��X!V��a#�b��%����q�Ƹ��Tc:����l@��0W�q�N�\��დ���|�|�y������2L���ް�_c^L˸
Xԇ��(&�7�X��U��1�n���GI�<�.�����;��������MGoZZ\����|������;���LM�^����g�=�tgj��~y��?~ꋏ�N���z�*���E����ﺵ�z�O����B�þ�� �2�I��-o~c�5�������^������G�������w=��*Gsp%g�V���YQ>[9�ґ9u/``um��0[cX+ɊП�N�[�Ƨ�>s��9M�nV;�^@\*���?5�9�y�bi��׼��%�l��ccN�9���ӫ䭼�?Ǒ�e(�3fp�p�����w�$`�����(so7�-Ƽxƻ�g�q@k٨��~��tӠ ��n�ߌ �K��K_:zӡ��˗�����k���	��M�O�����ӎ�����G��󒧯�Uү%�K����;>��_��=���5?7;���G?�?�rכ���W:��M;w.<���C����� �D�$��%�
 $���z(\�
�Yc%Hl�c�������5�m<��e89� 7��U��)r�፿?�m��<����<x�������U^�b|�1�Gc��5u�ž�u7��ny��Ԇ�)�Uw�1�����g���x�
x�*�x7�H+i�/��}~�������2��t�w�qە�;���_�B4`�c�~�4?3��U0'�.V>��z�f��Wi�a�޿���������O��ϷZ�dVpQ��,`�B��H���������������������'��1�{��A[fg�g"�Y��B}bრ�����ejx����������4Rqأ�Bԁ��l��)@�Ӛ&�G蜩�aW�}�j/��a(J 0b���~�j�:[R��<��`��/s�?&��++�V��#��X��/�*%��HK�xU]G��vbJ�Yr�_��~I�r�O&�`0���^�
X��,}�6���dI��(t⦇{$jY�P�u��������0ݬ#�n��}�ˏU>����I~���5�=�w�����~�S��,.�D<�2� #Y����Uf�����[<���kR��o�y_��5����?����(Rn�r@'D����_��Ks�|��;j�c�����7�8�,uX	��% ��X)@�+���\yY�&C�K�Wg���CN�����Q��y�n��a�2��N4O.��l2�
@а�g�cI7�<�7w��	�MIO�(�ʥ��;ؔ�IBoq�9ά,q�D���C�L�8K��w����4������7;m>i��Þ���}�L�g�o����0����'�no����='�y��Lw>����.��_{��������g�x�׈&s����?� p?����++��w�������'�����y�Ϳ�ꠍ��_����ן>}��N���X�`��@�E�簞y�=j<�#����Xw���\}Ϡ7�Z����O�{ En�'�{���`���lq.����'ee�a�'�2>z�e�ў���vYB=��3��%�|�`h@ή���IK&P�wpB1&�L�E.�q1���0�d��g��W�/q|�=�q�:�YTV�ɞX;ELEAU�6p�D���]Y�����S����<����Q�2�W�c5��ݲk��?�t����ľ��o����w���'��?�!&2��(���w}W���~`��٨l�}Ӈ��}�)�i3���2�fP�d������.mԖB�_86�G�XN���/;���P�A���I�ͺ��B"��Ńn���%�|�4�������O�K6��Hs|�'@56 �~Ez����t�LZ@�=��n�_y/�"jDb��-��%������r�x��U�7�ǶE�.��ږ��
�29J����n���t�������߶�4�n�	6�c�(�م{�6p�ʕ<pח����}�o���~�\^^Zt)�\/b�^�-ߜ���w��Fgu�������_��ĉ�Qߔ+s�����11�`ʰ���O��$0� ���GN' �2��
+Ŕ����U�ygu���A�+�4�!E�٘��`�|�?b�*k�
�W���d�1y��q�x��J�Y�J������8X�����U�s�tuf�ysU�����w���iM��l^��0���6��w{��T!�Ὂџ������(��͙Ji-7������|��e���Ѵ!��K˨�w�޷�o���+��4�w�����С���ǿ��}(���]�>�D����8ל�;1�X?����/���3�Tv�H�n)ڕf}Z�GFEۅ-,̏�.���b�5�Ӡ����.J��ݻ\_�ɻ"��H���ߊr�������&k6�Xz�ہ^,��Y7A�����+�Ҏ���ɘu��t���� �"]� ���}.��v�V�˽���b��b�����/å�����"�嵮�&{e񩩼āY��Gx�Ȼ��{.���o;y��#��Ǫ;�8���Ղ�-_<�w���kZ}]�޿��ٛ����g�y���wJ��Ξ;����w������w��?��oy��O5����d�R� KL��<���h��I|�R3��$Ga��G�E���s��n
�r%d`h�J�M�E�֗�5�|en9���qF�!���6�h\d2dp"@� {^��bS7�'�#�JT�{�I"���1�`����C\���O�1���s�{���|�� ���/�mҮ�+~7A�q�W�"��|��޽"<ޭO�C�}|V�)�ehEty���w�yw����ؘ�����g^���zh^�"��lk��YY�y�7_�׾���������F�y�OY�������Cϝ~�飿��qЁ�3R��<�����Rg=D��st��e[����	B%v���<������>�G(�"j����e���d������g7���䃻`�ar#��E~4���@w��2��JQ� d<g0�-�ρ�/��ǱN��8�چln��R���pԜFx��4�^�I��\�&�9�����HW�޻i��՟���=�����{ｕ���ﺀ]����Y�� tn6�'�X\h!|𶩩�S++�U�k�d�k��>-���ɓ3-�E��D�������z��������/}�ᣮah�X���y��Ƅ��
5�ᓐ�� ��V��4VeT1a�G�t;rǜ?���9����@��(���������E�aۭk���b�Կ~l�=��v"g&M8u����4/��bW�ѳ�+�l�ٕ���:rJ��\6�|݆[��tH�+N�����Xp��"���r/f�k����t�_���!(�e/H�ۻ9��eC׉u�]�|W㰔������ df��=����Աc���_S�?u0�8�o>x��W5��D7l���<��{�a�"9�v�J�����0\9��c���W��ڣ���k7�v�.����]2����\h3�ef�AD�W�#L��o��]��sy7�b���m��e�X��\�l3��Ï���h��ޏ�j��6��d͉�[�R�\b��a�n��Xg��Bf2Y3M�`�x�����^N����`Jy�t<G[ۇ�m?湔���Ky6��>dx�    IDAT����O�O�9�g{݋�ڌ×1j���R̱�l��+^�џ�ٟ�\��$�&�1ק����=w���똼��:�����W�ugs�{#�i���TR�Jܷwwj�����4`E��e�Q�VY�In`u0qiy)Ů�̳6�-�6�☉'A� �LC3I��.�6���~��C�IT�n�aC<b����iw�x}~��cr.{1�bm:|���74h<�Įw�ʺ���/������n#f�����8^8.��z�N�Ӣ��nᪧ��t�t+�%��I�W���,�Q�z/����d���nw�L��/]��L�!q�s�������_��_�x��_�rՠ3���?v�-�^�to&��'�����2�|m{�����-Dk�klXJ�����+��8nip�����T� /�AN/Q���bO��s+���*��ƈ�5��P9�w��9̤=��dw�KT/�-�4�	�{����i�VByqe���p�W�yg��W��{Y�Ȋ76$�̬�(*o
Q%��Μ��7�]YM��N�>�����p:��P��v����ŝ�m�̯9t֞V~_�g�,��4�[�b���~��~f�~|.�x��~�]���2:{��`���`��UR�w���f��;�>y�q������c�f��?���7��9��G�E�<7�����'��X�����o��'�!���*k�i �6��c3QM ����	�D��A|OЍ�F�FL��_؃�,=!/�z��	b0�?f���d��U��\N�;���r�V��_H?��ߛ~�'�}oL��c���z���;̬�7�k�c-Hħƀ�=������ ڣ������}��!�O1x2=�!��ɁhЇ2+��eؽ��$�^�[�z�Aclo����x��ڞ����a}��ƫ�gY]Ӯ��/}	���i�'�|<T�kk����;23?�.����<\����]o֏*7�(�����G�{�P�͝;{nJ���-��#[��V�пkC�ɀ�Z�����G� ��8஀1TS������?�j"B�����B�i)\<89y��D�=s�R�;?�w�;�y���׼P#J�Y�ȅĤ{lx޽�^0s�e�+�9�!�� ����g��w����w��~��>Ė�+�j6����l��W��(�n�4/��!�F�I��<��:�=���%�k�Z��-'Wl{�G�?���c?�c��[oM��ǂ���vгէ�կf���3�v^Y]�ET����l����uZ��ڕ��Ȓ"c��F�u��r@��a(Q�~՝�0�;�t�W�� 0:jE���c<2���8gH#��Dp�<K���A8�$�O����Jٻkw�����t{#�G~$���X^�H+4R1M�⍃C�:K	f)o�%Ͻ�3"�u��"����^��q���tӾ�閃G�/$;�u�?'��^B�xH(�$G�Ř�k�'���k�y1�M�1��{2~�帓F;/M���cq/~��]	�B`��Jw��#I���ߟ~�~ ����+1�T{��T����g������6�iHC��NW�?ɔg3r<Qj��խ��͹ʩv?�yӖ��% h�W#s�1]"��ݳ����,U��W�^���{L�D0DD�=B7q}6G�ʂ{�?�?�~��~*zOv�ݧ�v +�LM�R��@����Js	��"�2�6lv�Μ���"+�s�3gӷ����w���c���
�|N�=݆��5.e�T���z��I0Y�k�O{��)�-���Hw2|<�G�>���/�|�L��Qc&�����Z�݀����/~1@���iP�_`�Zm���5��=!ou&� �W�;v�sG����÷m�3���򣜫�&EZlp��^F+�xg3� ���\B����! �HA��n��wWgi���Nd�96�J%�F,s%=t�6��\�cu"�I?��ޟ~��ޛ��?�����/_f��q�+�zZ\��a���B�O�G�xfc3皱�� 8�"��9!:��Q�NU@�8~2���#���ߖV�	.^^IQ�'ϞN�◝bI�;z�Ln��c�y/d<���=�ԡ�6(��*NbB�����qz"bO�����u`Ᾱ���tB\���w"cP�d��;�U�+��w>Bw�"ꓞ�Cb6����=�G�%�%r�jS��^P|� u���<�ݿ'�20�ڷ� ���$�z���` ��\S���[V���o�;j����ڿH���:�I�R�ܙ]��}+�פ���yw��Jq$.�U;�ڈ
;w��xn֚�s�A�_~�{g��U�6�)I�R�ڳsGZ�t�6��e�2���X��(��UQ������:*�U� �� ��,�an�R�f{˂�m�4���������|:�z�5&�R����r[Ȣrw��L�������	Ĵ%Mt���k�->mi5IG���V�H�Bs�͠��`�r��d\���	46ƥ1L�d4e�=�=��=�Ju�s��&���m�~���PGG���y�Ec��f�v�S
�I 춞3���eoȫM�G�$V�&��zZW��9U�l'�G��V��8 �ҕ����X����t�]w�!.'\z���1���HZ,ɽ�]��}�|ZcAm�6;]��dznW�8B}�͙M1E��M
�9T;fgL���F+����3�G�T������ԌϞ9�����Jg�.�U�p��.���E��Z��^��T��aB=WU҈H6���Y�A�U����M�n�=ד�'S(�W0@j�$�����'�o���GJ�(Ø�n�5|��a}�4iykLt��aG���I�Q�jm�ڵn�y���w��<qb�I�>0�=��9s�|�BX�R��,h,dl�3���E��eL��;�
�L����g�� -&�bU'�._:����7�����I���� �9��tGD�H���u���@�����_XS/�����`F$k�����W�퍛I��`�TnL�s�q�Ip�*�g��K�2х�2��uy��w��">�ܩ�O2=�����w�5�K��w�#��W8����$"4�<�cj!��wa�a��H�B��,�|�n��:-�wK_��R�M����\��/�3�-v�UZ�=D4p�h�Vf.���Vޑ����y���>��K�R~������!���tkz�aW��Pg����=��gb���(�<o~b0�����j�R�%�<��X���D*B���kz�h���5�񹲲�J����p�}1Y�L��ƨ�Ђ �yuWN�J��Ҁ��2;��h:jk�����BL�BC�1�x=��"��R�yP�i�Gn�����?�D:�[ED��Ag���e1�-1�D$ٍ۱W�*��N�G���O=\���Sy�M�u�政PQJ�lț��!�Rli�I �n�+\�pk���1Lwm=:�)��T� ;��~�?��������Z�-�:�;��z�'�2C�G�՞��*`ɉ^����MfGjC���AFs3��啥E�I�:��p�(�8�n��c��[�i1�.s��	���Y�m���]{�&�𨁟�'�8�y���3'�4@�Xe��3�	Q{p�S� ���p���rڀc;Pu�X���Ȼ튬��iT�jGPq�/�_�#}B���A��H��M��80���{<A�u ,�bn@���6��t+{뷥{�}]�(�?{�f7���W�*���X׫�0��b�i|[�վ�Rҭ�W�:��\W����D�J�"�M������K��p�˭����^6��uc����/|�~���[���Y{��z�F7?����}3d�A
Q��N��~&���	Q�0�K\>oAo\�lY���� ���� p���q;vK����u>~6��}�8_h�S�{��kp͓�}9�/�O�����Ѭ4��S,5��0�߿l����"�Q��C�'r���54B�;������!_ I����J#08�>��	����[̊�h;쭧=��|���6�z�p�̗K�?��\&����'�oV֖kKK7c��xs&cis�r��������f��>�V��h�]x��lH9��0d4�g������jL1R�J.$sבu��n���+`s��a�x��~��ʕ��F|pe����& �#�k��HX�( Vރh�W��W�L�+��ь镟����M˖�@<+����-oyK�G?���Y��h0BW>�\�s/q~�n&d�?�h���Ӊ�T'�,��ڼ�m�В�9�ީq�lҩ���
RW�y<G��$.E�S��&NդV��ĭ1S�R����O�?�h|���f9.Ã��hI8c�m�i7~j����sHP4I�u40�� �T��Jm�"����(�zy7/ l�.�:�9�W4�q�e+�\���S��ǖ�]{����)y�.>���������ǉ�����upnN���8g���ݜ�\�6��w٧�n�L[����֮�*;�LI{Av�w"�,��rU��6n������/��ϥ{�]/,q$�M)k<��G�F����s���=��� j����i��5w9��	`��\UY�� 22 gZ+��(|X&]D>_ر��E�@�Z�/rT������6��a�3����~�i�H�k⦶D �)�f}*��*��`2�f6�~������v� �RS�C�y�x�\C�vG#}��u��*���>y�Y���2)�j|πͽ�n��g�Xb❚��d!DF���j���l���zm��޽/����p89����B4S��� �%[���}�p�K*-��׮�+�˰7/�{m7�I�����ݖ��?��t�+_��,���C$oʦ;��,8O<�x:�g��9 �gQ���"(׈���@jED��8���LZ�f)�x�7'��a�e_h@�sH�N���K����N���,	�R>������"+�X�AW^������&J����Pi��/|�ߗd"��R��_��y�nU�t� o�{a�����T"_姸��r��^6�F�g��Y�g����n�\e��:S���1���Tk��Ũ�77̹I4F>N�68T�c����f�hip�b��d��f�6	q�FX���X�r	�sӄ�$����3Ǖ��>7�/?��;����'�����4`���g>��t��ϥ#�ȧ \zp� �8]8��r�=��gʕ��I''@�4S�3i�!�Ѐ�j3<yG�H���x�w��~=f�؁���j��`�\@eAN���~6q-M�M��V���6�r���}u,�������S'��+i`K�]���+!��%<����h�lD�VSh�s�؇�Q,�N�r{����f���
'��	����c6s�����ZҎ7A�r�oݪ��O��i�I��������	�L�=E�F͹p���%�����N`1&�x/�;
[(6�/a����7���W[;���E���ۿN����L�?���S��B.?��G����t�-��>��5��2��2mL% ��Tī�Ь�����9����W���'Ʋv��!��@`��9dcW����s|�δ�N#
]^B� �X�iL��-∹�>@����w���ѵ/�:s�1��-]F��F�~�s�Y/=|�Lڳ{1-!�HJ���1����y��VM�4�7	�C�E�V$�ա��2�<gcrح:,75'��lk�,�|�Dw��k���-Y���͎z����ʿ���d�hV���lo���+�-�o�/��F�c. �Lɸ">?V��3C�iL�#�m@?��M?�C�M�;L��Չ����i�w�s�O����i��*�r����. c�%��D�wbG�yԡ�"�X.��+1o ��/���j���������i���YH�j4�MT���Sس��R�B1��Qp�<1p��Qıspp�z	�3�����T��5*D,�^f�ٻ��c�_����Ef3�\[?g�P�c�1�1C�\��ľ��۲��M�1L~.�.I4�N��l��ڵ1E<5�ůq��G����{`�C؞�tN+���$εK1��K� ��(���k��ߟE\q��#�b6[,��b_�`���Z��7i��~�p�U\z�ь���Mm�N�;HSgܡ�����N����ʙ3�>=Bg�d̀uʳ�q�i	hMɓ���zS�U�,����q�v��k��^͛�tz����QE>�.�.l��ľ�H3`Q�"��*.�Jaa�M��ʙ�
Ո��t�|�5�m��ťt������ߙ�Yܛ�<r�5�q/4Y�I�����?�5��+3�l������L��Y23a�~\�>��\dKT�M#���ڨ����67Ĺ�҉v8� �����n���Y->��(��>s��-Ԥ)n4>�4�� ����0�%���~>�t�p���^���Tn����G�U{?Y���-��3[F��"('W�l?��ט�9���rN���s�1p�B�p��` �<i95�;��B�^j�A����q���!�Uq(��^e]>��i��KT��� Xڅ�S�|��o8v';�6��J��%�|��T6�7��,�VM��\�d�����~� >ק���a\�<WX�Ӵħ�/��m���eE�YcsL�5���������?7���m�Enؽ�~5��8�&" ��J��M.�*2lzɅ��AhʩT�7���F�NNeoFăa�f�n�@�'���P�~:��fn{晧ө��J�3s���I��#���Zѥ"��GT�@�2�������L�Ϧ�Y�vd�M
G^qs�߽��*��U�ˈY�d b�3�ӽŠ�M�tÔ8�y�&\U]e���j�(0vP8B���&~^�� ���ͺL���W��N���/=��	��ӈ6�g{/�Z�����b��t/��=ב�����rz�����l�+zD���
Ӳ�S�]���W���b��;�!c�{>�__k�EEO/W�\U\2kf�e>A8V���2��(ﮃƖ��N����*L�G��7����w����ҿ���v��B��b" �Z����@����'���� ��}�tϤ���d��3rx�o�L�z��f߽L�����=%ki�u�s�u������v���3�P��5�c5~�͌'J�@���%�p)�K>�<b���P�9�P��O���#�D,�4n��Aj��F���M�N ;s<�lV�[�I�?��t.�L�-�l��w�˜��ft�0�
=H��g��!����uFP��ɍ���a�Ϟ%4Y�ųV��?��`Q�GYۺ6�b���qbt"�"T(�.̥%���Oͽi	w���`���;���N��i���S�=Ϻ�`,Pf��:O>�>	t߷9��'*����W/z����7|����A'gg�d3L�4���~�QA~�T5��hE�Z�l�K�fĢ����@� NTI�/F\\:#W�n#[��3��ʠ�"{�wltJ���U���Ï�8�3����U�i
=:/َE�tZ�U ����
����N�O���34�@q�=ߔ�L�����ʈ�#l�� {'��C�S��̩��t6O�6��y�V������.PK�J��ٲ˸���|���.N��=}�u�d��"�<C8��Z��&s-��[\Yq�w�x0{�6<�Z�@�]�f�f��]Fk��
��	]�m�]n�z��1�,w������OR9p*����,�b� o0�|���=�;p�.�dЦ!8�)Q��)6 L���C�|>b�h*��;�B7:�1cRn�������\��o�����E>S:m5/gS��
m��(�zQ��I״����u�������\���KM��Px�
ǐ��S�<�q�ƫ���
�����q��C��;��bV���4v{F��R��5X�jg=�+���."����L��r�}�X�\e���n��]cʸK�]$5@��š��jYu7Y���R�R�r/��%�f�m�>�+W ���=�r���MG�
��	4'J�\��~ .@ѿkܨ�    IDAT���i/����f��mqn	SM'0<Mν0�p��#��=ߛ���J���Ui{Ӳ���XcA7�E��Efo3�ƅ�U�+����_ ~�����ao�r~�rN��ڕI�2@��8��q��q]9]YhTl,�o~�I)z�3�E_d���wߓ承Όh����d<�-딾�6���178���D4r�|�-��U���<b	{�5�nK�N��l޽̓v�b����5+��^�ܨX�]-��a�[e�-	�ƭ��~/*���[�R���{)p���_q+���XKN����^�'���o���1��0�OV>��͌��O=�N��ob���$)���h&_������U�jw��n��hɩ����+�Nm@���3�ɘ��)�A��6VH��^f�+õ]�!'W���$�w�1�֘K#���2�&�!wg.�o�3po��Y�z��'�����xi~��4˦��L�_�1`><��^{���矤�6~~�K���.�BN�L˘��xъ�d� �ԅ��f��8���+������ɺ7��.ǖSkWw�;��6���Ԗ��D��~C��ر���#id#�6�9Y{N�'��{K&M�dz �1�^�5ig/My.�aIr��؁\iW�!�����RbwP��S&����g�MSI~�#��QA��=!��q�������m�#P$N�Lm(������Sl�=�� ���Ɣ;u� �ˠ���U��C�W~ﱟ��������ܝ�e�<�P�-]A Y���"��&�ɷP+���;M!&bG���=�qc?P��2a48^x�D�P�o���txa=jG��a�̆�T���sQ��2`�N�q��y���K�}�2��W��O^�_	��������ۚ��wم������8�?�����(�ҋ�=7_f����R��B������l���}�oy�C��v}���l���O���#S.�f�?�m�e���4�� �%����If�����ʼ��Mk~G�^D�/�ٟ��>�.��\�*�ԔAϔj�n�@�*�#E��T�2wpb9�y֓�+8�j�dE�X.�xY�(�BKa�pC���Zk%��(�Lr:ζ�]�p�=;XW���f�:y���M	���8h\j8�7i/�=f�x�fo��8�sWUɻ&��{�����.#�\۸��4�����)�L��h�֎��Zn�!p�l�'S7
�Ի��:�9v��NrҘQ��/�.s�ܽ��hW�OƱ��mGV�'4�wя��w�}�S]�+ru��C=�?��8B͡�jЭ:(� �xT�~��$�3�. ���qR��1f8�!ו��d4ʣlh�T��+L�;Hko��i8#���j��ĲE%�3�̣?�%� �q�+ ��0į�t��v���� O�K\} ����9�P�^��Vqe'�ܱ�{�|��dH˝E�d҃6���U�d}�z�S�c�N�{�a�W]w�uJ\%�r�wq3�Ԟj��y���/�����ùy����t�����z��*�n�*א�Z�Gf�D�ϚRHߣ°�^�����8TMł|
mcz���S�����T
bXy:��3ibՐU��7���չ��9�6N�i�Z���No�����t��'B���n����y�yF�����}w��	�yf��W�bBrC��(�o6\Z�'�hq����co�p��+󦆈(�D6 O��!�=#���{���m>�t�Y��(���i�<�� NZ�,���A�;�O���[��R��;9n��Wȡv�G�bL��u��8}�2{_�TH�D@�t�*��ue�Pyө�h�X����(N�8����yAQ)LT~T[k�*�gk���q2��O���3������[n��@�XR�Î2�X
y�O?�R.@8��E�-��AbG��C���x���)v��%���W�F�md� ���K�|�
p�B8��8�3i�r��q�J�ҋ���#�4��Q����[����Z�ӈ�x����Mhd��?����+���0�<ɦ�U����(�)���:$��ȏ�Q����u�яW�� ���=�O�(G��+J\���ɸ��H�qVj=�zis]�
~��۴V�YJ�ϨߺbH9>���_MJAlW7���3��~�Ζ�&�.ݾǃjv�)`�~�Lz�G�h�w坲���A��KP� we���ݜvt�7����<��vz򋏲����&q�%�6��sPF�!V�8v��3셸���+��	d��gG��R�B�ɻ���+U��
�bo|qR-���v�� ::ɶ� �Nt��=�$���%ݼ�u�g�2~�C�׏��&M	/(5Qd�1mC�~z%���{�k#�VIbh��p��:f+��x��f�Ih�A8�'�9
2x����������)v����ɰ�LBU��_f�ȑ���E'\ �����I�����,ge1]n�*�Q@T �qHe�D�ͺNd��G�Y��H5MsN�i��C���ś��k�J(rDu�+;Fz�l/�&x�[���?�w��4��,4 E����e{�6M���8{�	T�zu�*�m�r�+jq����|������E�j�L"�@�ٴK}�Qy�*�͌l=�>�g����WBL��^Ϯ����r�R�L�,%�W�o܂
}>E^�.7`?���[\!BI�d�B�����ݏv��a���h��]������7��8�	9��+������	&Ťj75%�H���{A�I�@���7Ϡ]`�b�"�hQņ6�M�R�Fg���@�b�������`	-X�["M$8�)�[`Ƞ7�2��F%�n�c�θQ����A"�� �Ac�}��ZCd��|���сY^��!�A�n� ��]7�� ���36Je�h6����z+�.T
wk_��ʢO��('i��1�s(�)>Ðf]�y=s��~�=;��9	1��X�&�٬�<f�
��@)�ϥ �7�cEL\ž�_�o�n�������@A���'O�8-�t��2�3s�>�E�4M]�i���Y���M�z��SMO>�t�Ϟ>�P�f"��RY���x���&rӍro1��\�F'MN;7� ֍�5ʝ��"Ϥ3�ڦ'���lM�ȹ�(u$��l��=��g��L�jLu�'�vլ��x���I�����{ɧ�r?��8���S�;�u2J���<�q]�7��b�t���H�'�+�fƶ�k&	2��]��-�𺖮��4ۤ�=����Τ�#�xq�;֕o��x�=�-�w����dAg��\�[�qڻ_��G�\.�'=���9��p`��,����w��`����+�W�.Wu@�ϨP<x�X�b��B?�!BO�#��QN�J����G?��~MŸE�Cq��&��D�2��L�g.��g�2׭��ix��q��ٸ�Ճy�e�b&ӑQ���ʻ���&o�,��4��-�]�����s�K&<��%�.I���xŋ�����B���|-w��3y�21z�Ç�~���1 ���c��r3Ƶ_8��L�Å��L�Z`X�r)�LS������t��[�Y��i�W��C�"F�(s �J�y0�B�(�؟v��i��'hS�Z�O2������[���mc�!D1�SS|q�w?N�#Q����3��iq	h/M��~J����h���̻v���8�S���W~j�u��y�Q��_�l��K�����{��vB��$K���Ff\BJ��Ѭ�v����K��5o����X�IfA�0��|��f����"m�n�Ҡ��[�J���p�&�$�Y7=��
ʪ��q�XQA�l��G^%)��>�-v쬥�_z(�X��]:��z�xUM�渂4�p!�#�嬔��6Ċ�A�jZ�4Uo�Y�O�sY6�:rw��=hå!����ʹ����@��>c׃��6�lE��{���:*�
c�a�^�	�9D��ǭ��_�Xb��K��]��3��Lk�x��@{JFLs��}��ֱ�ԛϹ�sc-X�R�/�R��N�?�u+N<��g�&r<�vֹ�mϼlK^�����N�WBc�w�62j�hJ�-���\���G~���}ҭ<O��l�eiL��FQ��4kN8/�]��1�c#�1�/?O��t���i��<j\�R�h2�v'+ *�4K�@U�+ؼ������!�G��4J��g�n�z�q��R��U��v�<>?���+V���9�Uęqן4*�+qz/v�^�,�O�'�M>?��G��%.�Q�CQ�Q��/�3�/�z�t�}�;uO9�6�ġ<%�ϓD(�*�(�X���(�fl���e}�\�V�����g%�� ��p6.�C�W���
�\H{�:6���MԂb���v���"�U�g��B
7�3����@�d�GZH !y����R�Є8�2���3%�!�O�9->��`�N��<�Xā��YW����yv�	�0׵�W)W�Ǧ=R�Z�-��{�W�y/n>;�_�.�O���ne$rx&�#/�!=��I#J�fs��4�Z�&:mz�8*p�E=��@�%��^�}�c������]����ɾ��5����D�I, ��#8 T�[��\2�C��U#P �Z�k/ZR40eU��h��2ĄqE(�X���E<%�F_��x�x�L�d�Ы���d�S��]���n�vW�C��(��9zzo��~Eg�����2n����~�5�=�~J~���v֭��g�d�ʵ��Թ�'*m2��g9��lj��Y�s�(5�?���E��yL�YcQS
��@P��F,�o�9��x�	�C9�D`XeȲVqAbL�.�<P���]�'D��j���,� ��͑����R]d
~N�8qt�o�T�m��z�9�oEY���%��(�"å⧔�<���W�6�I��T���\�Phf�qEx~�mO�/h.s	�t�Q�{��'Aܹ��Uc�d��uoyʏƭ[��0���I�4��F����e�kv�<����S�7�ڼRn,C��	�~KW:�S{dC(��t"%�T��&ʜ�qb_�Ѹ�LF�+���h�o� �#2f����rq3���+��	ϓ�RI�ʗn�s;Si�jI���q��(�nu�+��X"1'�c�]��EOd��7��A��`l��Y������]��w��E��2/�[�?y��ڦ�ơ�v��1"�q�tӽ�*<��n"N�1;E-�{�߲K75.�r�jQ?����f6B\RtAl1я�c4a��U)��%���տQV%\�7o�\��f�����c3�R�=3��Ʋ��2fHp���)�'��䙕XfH���R���R
:i��/�p�$������6�-Q)V�1&�D�'��g��j>W��K��	���p\p�yw٨������o�ek�vW�ɉ��+���p�r9�x4K^�Lp+�N��`΍"�&�"�d�uW����ރ��1��z�HO����!��qk�	c�^I�k�盎Jw�~�xL�'�[��l���0�r/>�~��-��>J|宨��l����E�my�#g�q,_B���͡�zy&q.^�Wa���5qN��۵#y2�y(��n�BD�����$����s&^8dhS�Icr_-����0���?z0*P��&�<��6tYk|�����qؕ:�r��KC�S֨�膛���>��<ΨQI�B��ڱ��S��l �4��%F���b�Ʃl,��g��J�n����2ZO���h,�߸������r��.u�����LXIE�F�S�(�n�n���a&�e:y|�{ae��Ϙ����ɸ8�v�<;׵��Fݵ|\���1�v�og�x�-�x�s҄;)�ٳ'�c�� pe��1�Uc��Ӕ�o'�����f� ���`[��J	VTLTkT�r���k˱8^l�{�c\�]N��ӓé9�r�J�AZY��G��e�h��Rc�wcn�*����Ԃ9-t�Ư~z@���v���;�?Շ�P������B�E�z�7�(��vY6��Ǹ��W�uP��H�OmH��6Fp��H����#=�W�����L3�DC�ԏ��|E��3	҉�!��`����ə�তY֠h��ˈL�׆ g�i��ш�ǽ������2"ש_0s��
�\��K�� aͤ�)�;���`���@.v�U����Le�sL���@	剪����̠����$;P�Ո�Y�sx|� ���\�P�� p�X"J�h������i������8g���y��L�7���J�of)0DY�Cɿ�&i1pl K�B�w�!�(�b�8C�i��pDilҧ����|����>f68�\��p�ݒw��c�����9iv��RZa��	m<���G��,�-
P���^;�K1�/X'�v%���Y{3i7N�d\bi��h4�hM���ű��:�x &m��+�p{�neuu%�bJ>����	��Fؖ��Z/��LU?�g�}\�ؗ����m�!�nN�>w߁�|��I
�u��:��YGD`됭R4��д�]���SE��w��;�O�[P�p��nK~��}��1΄N����qܑ��,��	=6b�x��g!���UQ��'	�f̥3��⢖���\���a�aXXa\�H]�A��p^փGħ_�/�(�s�l�L^A���.^����RA;Mq�~�X3!�ذc�!�)X��?�ȱ�<F�+�̤�g���p���V�/�$� K���终%C�s賶#87*�ؕI3 '�[]O������I0�]�+[���C������G�����x���_F"�
� �0c�����G���Blh;��-� qҳ���=�����5�N��'��ES�`ײ�c�{�A^�:=�B|\�5�S�0���p�&��|:\�v!�s�3����)��p6erS�1�H� ġ��nQf�!)�`l��z��(�,�xx|��S�߯/(R�µ�XS6�n!������A����+~J��x,"�'��/��ӂ#���}��K�G}.G�H�գ}87;�)�{ �
rni��`8����%��g�-��z��3L�|���a��sQ�\�xMO�H��̉�-��^����'3���p�9 %7�3�pSzF��4z�~�<�A�nPX9u&��.��l`��j�@ˣx�g��вxn���ß"_�>*�Ԇ��C|�Sк����Qoƣ(1C|��u�)�'����7@������Lm��1��8��J��K�r�i`jn6�O&$Ի�i+�L@�,n�v��i:�& �d�{�cm��x˞����e?9�����g�A�Ϻ�@BQ3 �/������p�h��c�w������")��绗 ���,8�-
o׶�X`�)���Y��׏�������A0h2��!���Y�	��� ۅG~�`�])}�y�*f�#4���8��1d� .#j���\�p� Gu#&8yU#�D�i��DB�H��� �
j9���*���y,��	�d��%�=ӌؑ@��ir��5�=K4�.�q�����c��F�#����{D��+E��ORc����3��o�K}�z`��`�4��LS�h�[��؟��s�My@Qư��g�[i�c��٨���e���$uɚ�{8jJ����%z�Bܒ�R3�cEX +�g)�	'󿆑c�0� sx�k)g�S��$՛o:���
�?�#~����Ө�:��z���tQ��N�ʋ�o�y�ݐ{Q�O%|(��c��` �,�5N�m*�S�~y,����3��Ď�U������~�2��թ}t�Iy�U��#��q�3;�1c��^�g� rA?����� ��0?��'B��':&�G�6kh�t�0��]f���$�H>����q���"�[v���u�U=��&�e����˰d�A;�牯>�2�vݥ%����"��}Sv�t_�OM�%�L���'K�5��w+�L^�X�r��ͻ��n~\���J�RQEbԘ�ڷo_�}���@�.��AX������d��;wO�m��]�\C$�4�s���'RJ�,�*-���=~+�ˏ>��'��)�Ӟ�F�6by	}8eS5����9�(�    IDATw�3=�g��&�Hs���<��_����3ir
GV���7N��UN/ӿ�C��(��ʹK^J����[�_{�7�����n	v
�W�c�m�9�_�hO3�6jN���#2!�q	�`��+b�@.��O"L3o[�B�)���R�Cę������#�.���^@>t�P�g��X���ඞ�z�Uw���>�X���'��/��Q�H�/��a0�"�n�A�z�mX~?�md����yn�K�e�93{����_��:�uv��=�:gyZpw����؞ECq�˜'q�)����g{����ۡ	�Z�GS��:�I:ƹ�p��F'�e���i�o�_|��#t�-NЪRF�J*i�g������J�/�I/��-��ͷ�~,���y0B ��C޶��+�(^Z�>��Y�ʍԼZ��ze���jYT��$��4�����9
O�̈P�s�Y�sC�~��^�P��ٻ�@����Tf!l��R6��@�ZF�P��R��w�h��IS8�r���zF࣏>�n~ű���*i��c-Lϡ��0Ts{w�[o�5�<�t�G�n�A��g��t��G:��G�t�a$�XDðB��k '8��j9 7�7ה�ʳ�=�S���F��i�:�*c�4͢,�Că��Q�Vz�b� �F�=��ic�*^cORz�V=U���t����;�ǂ$ft9��A����Ȅ�~�a�'�H$) �?�j����r��ز͜����Z�-�\��S���������W�rD�K������;W,�hz���+�LX:U�Uo1��P�̖�����{d��ƻ��2�	O7�lt�����Ox����/����BT,q�T��c޹/���4�§�l8���НU�!~bC�+�j��˙U�
��a p��/�l���,W�ָ�+� 	��PM���Xbu��&�'�gt�ɱ�VΖ���xl3����"�q-��	&��l���uΰ{�cS�Q��똿�Ӿ���F~��Qz��7���z�g� [���sg�rZ.e�.�Y���N{	 ��)륷��>s�Ro%�ڗ��]�^�n�z�X��b�b20�ʄ�E�����z�O=�A�!s�9����pfpi�@�Հ�� r�$7R����R
�]�܅�Q��Ʈ��%pa?w�8��[_�^`}����St�뜫� ����S�Z��=��9k������V�!%%�Fqj�-_�����p:}�SL߻@}�]�b��{�Zŝ��nڵ��q�B^']Lp�@�h˕,p�q�N�t�dތ��l �F�jԸ˲��1`<N��Q[.ӀOP�5��(*M�Dx���#�O�n�o�W�iO�U�K}��2h����F&�FFw�C-��u�������;�b���9�u�1`0��L��>�	�(�d�{y��h{hݳ����y~�zS�zU��sW�����HcG5& *��W���b\K$�J4ѨK"*�(��Lڤ����z��_U�y���y���߹߻��۩s��;��>��ϔ6�����d�}
���H���A��>�����X��`�Z���_D�}�fX�dr��#�0���+}���"�2H�hL�K���Y�u,��!F��ƕ����h@�_�}P'���|GrV�K�}/����:c��r�" ?OZ�Y�BP���R����o��%�o>�!���Am�� /}��.�ZX�ݺ;�a��G,����h�*>��(6�+;#/mCf���F�]��9X�!u�0�ԃf�*�W�];@��s8�B�-�����'���L��P<� ��my��`�[�Y���m%U��.�\ i>�я�?�]"��$劣㉇���'��/{�|�?}�����*�ts*u�G��&�,�`25��s�	�GZ^M'Ւ�P/�Yw�<n���*3x�3HK�GX rP��fGل���byy�C�� �>__��`���Y� �#dx�0�ut�����:�A����*Y!�{�=Y�ztB��]�=|�X���B�xɅ/��0ccՃp'K�z����k�{�A���6ôv�i�a�̕Z�T)�Ç���¾(�[^�)����ujXǛ�!
���������~�BwM�n�Z7%/�ҕ��a����,��Gx)I�J0֘�XF؇}�)�� �#�],q�`_J�D�ᒼ�|���W���8��4��Y||@�m��C+�E^�6Y���p����S �"�]�Jl�0�-\�E��>�7r��<[����;9B9]��CHc�apsQ�IsS�.�&�vz���b�;��D_�Ǿt�
�ȭ��b��TG�(jt�� ��.�ϰ����/�y�+b2msQ;����v�|���>����n�Y�c{e8ͪ�g��W�~�io�%"�+4��E�r��N�+��E��? �����ijހg�Cꬨ��TY)UM��?�2h�0�n:�q��4���y�9ܘh"6
�1���d�f؞:r��~�W��ѣe�]ւI�����#���Tkܫ}�I�AX�X�!��l��r]t��6�:�r�ny���e�r�0Q� �u��c�2}�f����W�z{RF�_���+3B� �HV��L"�sZ#;�|��~���kR��W_8�pǟ���뽇���,���BG�'�!���m�L8�˛Ij�ݷ;e�$��.پ�U���m��n�*èˢy��:���y�j�;��rOL,#�������B'E�Rڦqn��%�fa�w ���'�Z\��u�0�9yUW�n�2������]��q �j�`Ec��9]�X@�`�v����2��K׮č��<����U�e/׼ʅ��D�ʮ��]�����GG�����T���ػ���s��6oMn�@�7�P�z�*����k���W�3m�.��2:�$�g�}�����~qF	e�hl��X�P���Ġ��/�s�/"���D9}�s���˕�&�Z`Ak�Nw���^��˰4�,:���eǰ��َ������[{"�f���1�Ș��햺a3\�t�e/Mϸ�{#�!�{��u�|��ĸ]��2�;�}!�i!-���n@d����S/j�(i��w+�*+�~	�t�-�i�c8'���+����z���������c1���y"��qx�cg�+�Ǐr�p9y�ly���r���-.���$���π�Wi��R�5ʗ��א
�xuӮ<����s���4�2�]6�F���R��$�ӷa[�i�}�ߦ $�q`hHYt��*^<�]�f����}�K�Ɠ4����{�9ɾ�C�+tD�ܸL���!��Nr�䅛��o��r�:�� /��'��u�E=| �Q�w�{Ͷ]J�tT"h�n?u��?_֖lb����6_Z\��`����B�����l�fN��(�Q{�!W��mv��j�6^kP-�Ɛ��.����;	ri�g~�g���
��\ElJ桪��{��-�'�)w�yʚ�j˳/�o� �i�C�<Z.s����\b_ƥk�� 4&����sM����:��n�{��D�94�����:>H3���Ç�}hk��壑ր��,��$T�����0�ց(�v%S/�J�������3L����۵n��H�Ν+k�9�|��r����CW��Y��2} ����*�!U��z"�f�9�k��j�gx��z��ba�n}��s��񡺵:��g_�=>�Pg8��̛iv�-x�����`٣���ej+4XƬ�i�q��g�D���K��+E_��̓��0�[�E� ��������̙{}8��a�����s����9��.g����Ʒ<2����(\at�gEs���@4�i)��?^�����;0`yُ�7��Ȯ�� �pc"�������8Q����U/�߀�wQ&���o��j��W��u�g1Ǐ-��=��mwvЁ��n�C?x�L�f�9&������_�^˪�����<���P7/�6����	�k�l����@K����K�C�/�7�YgU�1=�V}y����Vw�[���˰�я��S=��Ą�`T�E�N�V[Ѭ�z�Z{N=û_�m�����ۋ|�k��B�?��r(�JL�\)�}��p^��Ξ.�O�D��U�9ͫ^G�3y�$�ο��$���}�;ʑ��+H!�3!��_��+R[v2�I"L;v����L�@�`cAyy�a�^$Gb��-_���P�m�~�J+����� ��	��Tש'�����	�M�4��8�4N�:�$�-R<�E:����.�a�>{��2�47��v�X(�i�$�jl#/�m�W��6PO>T"b"t�Ni6��ڲ�����P*rL�2�&��-o��<}�/�������I�_4 �M%b�_ڳw�@�0���O���{O�<�n.f��'>Q~�d�����@~���'���5�2�:��$���,v�~�V��=�t�^z�<��K����/����x5Ŀx�f��~	���[� �N�kN�;Q����~ J�]�*�b>d��5L����PnE|�L��7|���y����ܯr�������8��nB՝*��g8�t�C�i��o}����+���o�x�5.v�_3EĶs¸C%�J��6�u��"�8�m�&��m'��/���ŗJ�K%k��R����Oݟ���k�ݢ��:��r�P�rsO�*���гb	�6��@V4��Z�T�~ƕj[q�l�=={�1�q�����s?�s��ʅ%*�66��v%�?������w�Sw��,x�/�zyd�׾x�s�G�����E�B�vʽJc�܋ �
R)��@Y�I��`�(����CDs�A)�h�R$���S�J��{Y.7h)֌#X��0��@w����O�>U��ɔCls��-�U^��'�;KY��o��|����*C��W�&��%~a+<���r��G�9�����R��z"v��AuWe����~�_?m�V։NcX;>>>Ć���>��%�N����-���pC�/OdWi	e�U&��m+��U�;�5|��� �eC��C����L�S�?��?�����}eY</�ԏ?d��Ε׽�Ay��w���@F_I�JB��g���sϓ�v9{��������;�׽]��{����S�EQb�aѱ�@.���^6�TI��I#�^q�(��:wȼ�L�k����+�n��JK��bXW'}���h��\l������,&ѹ�!A)�OX���:t*�-W�y{��#�!u��Y?�j�4���0R������Ȇc�l䷧�?�����iy�E�ݕo�l<��c���u�eЁ�̓��y*&D!]�+��,T��Y{T����'��`0�At7DR��:n-EN�"�|������h���"��eq���r9ľ���J!z˃e������/3��s��+���2U�T�r����}��W���ʣo{{��O�w��@��R9���1؇c��:݄/�ϲ�zJy���j�7+� 䅀2�X�����<E��k�O ��K$�ѩV�J!P[��r��st��3tVz�Q����tF&� ����w�� ���O>^~�;�o�+�"\��)W���8�?�d	K ��[}9[��R�9� �=��Qu��\$峝�#�A:;"����n;�p�'+ٴ!�hñ����j*�[�Ҡpg��X������ڢDuO�/�����o=��J�2�Y[Z�9񥨹(
,)Pl�F��h���滩௨�* ����Q�����n~u�M��G�/��/���/�}�S���P*�"�3�z,� ����xac����o��R��GˋO}�얃"�#�tVHf�?^o��o��x��c����O~����rm���9�0˰��{._��mNf��/p�:,0��#�N� ���}��G�ܼ����"Ew�ɖx�G�}���(���,^[���'H��R����\9���{����K/���e���f�{;�+�_��vKݸ�\{m��b�{��]}0n��K�hC;�vf�-\4S�D�r�vg`�yWܽk u��%���B6>;�~dİ�Qq�Z�D,t�ӳR��t7^�B)2�/Q�	A25�.�p�=����c*<P���"{*����}��������r���${T��:Q^ϵiKW�_|�\�t��G�Rϗ�\������w�w���l��'>R�O��2l�
TR6�rm_Cj�	�$�f"�`cr��I�`sJ��O��0 @�N��t�CƼa�MU�~��s�Pec���7�8�����<Ĩ��������T.(�c Q^"D�An�����M�m <S"�~�T��l�����ƻ��M3��5l�,�z�%G9���u���SǏ��ulǛ})eٌ'���M�m܇�|
�
d�J����nW	L���~�Q'b"N��m8������>[�����_�诔ӧN����sL�\ق�MA=�{�[�¡ٹ����!x�w�G��Λ���Ēa�:y�{I�p 驏?���>�Py�����(o�?�����3_���PP��T`���i؇MV&���
�<nݘ�S��T��&�<:6³�y/������"��\g�tw���HM�����P� �U�"I��]�  vÒ�M&Z�+���7��s��t��鮞�0���6�s�cƉ�`|l{͎V�s*��r4ٹ�{뵻N��I79V��T�$��9���;
�"���B}�5n���5NB�w�R�!]�D����r�r�k���Ǹ�b���(�Oo��G\�F�D����!��}���������,�²<r��p�T���/�0�-(���j9�}	��9&u�H������3��7<ZN������ϱ�jy�=+W9�ӑAhw.��ߌS�O|���o?�ˁk�ؓƔ!$#��a�U}��xI�����L�(3\J��u_���T�������r�����Q��2�F�щ�� J:���HD(����~4K��ٶ]�nڍc=vS��}�9��:���
G��閺��Έ�%�_���.��2�d�X�~�IFD�~E�3Q+ڧ���fX�0�����=�*�13�#1pUO����z���P�����py��'�����~w�+���,z�y˛8�vo���*�s_*'9ox���T��^{����8�����ww^,�Pko�;5�t�*'�,XO������JN�7X��D��{O��������0�T�-+�$�}y�I �`*�d.:��p�m���e	�"�����˧^:_�g�<�,��ѵu ������|�+��D{����6���7��z�>m�������eZ��eD���s1Gd�c�$}� Tfo�o�LV�P��5
cO�*.%�PVJ�Dm�v�ڣ+e�2nW"�3l~I�[~T�(�tDr�wu�ӽ���Nr��;�>����������Ky���P^a��̜bE_O@��j�Uq��c����ڲt�Ry��,י�=t��6[cϟ/���\y�����پ�P/=���R��4���S\y|����tEE�PLe����HƦa-�^8_ƨ��������#G���'^g�u�P��Ti�����,{ş��/�=�)�!۔�%N�ó���
;;��x`J��H�D)���^�j���2TƲ��m�l�L?۸�f�4g��eq<6(K&q8|� ���Z�/�]�`ȑQ�cD�cI�m��ր�6�֣Q$� H����&�:��u���K��d�!ܤ�]�'�\AK�o����_�I����� Y'@��b-i�����sr�0HW�\)/.�䩻�r���������S/���@��*w�3��W��*���xq��O=E�&Fǡ�R�m7bQ�gΔ/\潝��[�	��@�ˤc�fZ��vO�-��MF�g��������֗`n���QaE�C�GϤ��e�tY�4���(��@�m��6��-!3�n��6�Ե�M���R�IħƗ�O��xE,�\y�[��=����7]�j�dV�,��d)�L� Yqu�Cy����WU��I�w۹Z���_�i�*%0uo��-����7�jG��.��|��ϕ��?Y����P.��ܸj��+� ҆�(�E�A    IDAT���gN��P� F@����l��<_��c2:V��\9��ܸ����7�7YhD7YŜ����s�8��H��YB|2��� ��-f�7�\//r"� ��g9]j_a�:�H�J�ݶ�9P|�R�*,���9l�:�УW`a\Nw/]tw����<��LFzx�B9�v�ֶ�0�}����[���]G�8^��.��h�2o��{2�6m�p'�ԺڝTJ����ws�[Zb��fp�����_2��E�xG� YH�Be%(��-��3n�FI�2
�Y�qK�3�a3�,��v��cY��o��<�������/�{ j|D�Zd&33�/�\�>�p�v���G_W^�_^���ǹB�Jyy��ԋ/�3�ȣ0�;�\ִ�"-"������(��DP��I�D�� �_�I���/�/Ҙȴ�Y$N.��s'�[sey�4�i�ʣ+��H�ZفAp��8�wA����͆w�U�-�.u�(%<��g��C�ݯW�_�E�T5���*;�J"���aX��{�`�����g�M7��g������s�v<+�.%Me8�K��=��3��qy�hYrÒ^1��5��PG������|}�xj���π�����o�x(�]3R�&��k�ȑ/Bi�.���+�)�꯳��g�=4���|\(���BL(.�RzՆ�A�oe��!��^���N�����?˼Ef�'���jlB���N���1*娓/+�Q�jV !P�P� �Qv7-��E�t4�.r�J�vt�p�wR�ak�^!��0��p�k�'=�}#�`#��ٙ�m�����b?����8�ߎʪ �
L����H@=�e�-c�7��K����9��� �=ٖ(?Q�5�ye�����?�+�V��?������/������K������\6���Y��s+�<o}�����,�\�x��]��B؄��2\:����{����8�
]f�HVa�S>_�-�)?����,���m�.���֛[������t����%j؜����*I����aGb ��n�!aM���dK�xm���p�2��8Vw�T^=)y�9�T	�ԥⰛ���������(9X�JOr!�s�4���-�,��_��Jܪ��CU��~�'p�g�8]T�Ja5�+m8K�JQR�ǧzt�g�Q1�8���>�ܽ�o�D��f���L9�BϷ������.���P��Y�d���{v��F8�
l��8M=R&���M��a3L ��%"�w�xY��-�ܩ���9�������{�l�E�~��O�i�]��4�#�cJ���Ò~���A�@��ZVb
BB;�xȦԡ���*{m�9�5Sݴ�@n��e�������}��3����zv�dKL��wQ��w+ ,�)w�}���J���BJ�3�(��
Z�A�[�K��V�\���"@b�F)��m����O�B�\
���}cg
����=Q����o�[�ϭ��Y�[ҼMj�x^�C/��j&��\8R��)�t��N�
�TX��8���D'����8ļJ�����7�ȦsP���ǿDIή8�D<���r)?�c�Z�ۑ��wU���Oص�4�x�*�OexS�El�j�ݎ������ٸl��㹣úmno�o��*�\�)�h7t�=v��䬻�J%5�ns�ͤ������4X6x��E&I��V��oL#fU������4��*n��X^gy|�\A�6��T����_�_����?�}(gO�.�؉�؛��6�U�a�;#u\F�� "a�e��]e�F�:�ԛK-���}�r�ˀ���
K��������� ��\�:�&d�
7g��bn���;�����U��;z��E|���N�
��'�/��4S�|�Jt���闝#�m�h���N���a��/����RӖ1萦:���o�D�8��u������E���YT$Wea�2�V�K����5n���]��7��)U��6J�ku��y�SDl�1{����h���r������nб�UlJ���'ʽG�!?g��[�=�L�;o�\$qQ'������y����4���*�S��Ơ_��_-�!���>����j�0{N�fC�A*�{��U��u4�d���?����RA�A�dī����a��#ᚁ�S��_�/q�vl��]w�2������#\�C�����>�����;�(�cc��½��hA4dO����UI@O
�G�@�:dIa�~-(�w%M%�<�T���wѲ�����&�3d�6�����J��O��[����N�����_����Q��F���q��{g&Ƽo|���?����E�;�I����=�����+>>5����F�o#�dס��^���� ����nܧ�;�_B�?��ߊ��D�t6����X*k��$�҅k E��7��j%�r	��u0/̱�K��Wa^�"&u4���?D$�"�m�"y�v0�TPwyQW�iƓHU���ŭ��zf:*�o#�v�$ ��O�DV�qC` ��!��>�8�5b����6I�һDp+ 5��OVl�������a�צ��n~�L�%E�R�'��&u�Ke>;T�3�Fn㛮�<s��/������gΜ������c������Q�ao���zZH���RVH��Fc������O��'�=���(��zjh�b�5�}'4��v=�~P���K��Mi{T8d���]R5|g	���j��������5t�����@�*���c��+����ddן}#�� )���$��m��k�y������T�'�X��[ [�[�e���i���	�L߼�O�����	��O�LO]������5l׸�3��|��T���g��X�W������?����q�i9z�K{R����'��?�٧�ɞ����ܕ�G�h2^ ���Q�`�Jn��d���kOU���d���!osIus�.�6�܇���/�t3�=u�f�q�!Ѵ�Sֺ8�S��e�LYj��!�^�����&�*���^J�' 2ܠ=��&r& 2^��l����[�5~G��V6���t�e���]}�9�F����'91�UV_�����^�&⎡Z9�2+�.���쮄�e�أ�NӼ���_�AӆKs�*���K�);C�XTw�f|]`+?ߔ1è'�mz��[?�ڷj���������������A�^��_䖣�h�6hn-;��g۹^��1��Oee�Z��O]�6f�S��?���xr�m�pZ5L��R��;K5��f���i��Y}�ػB�*9����e:���	}�$F2�h�և#�L�~
�q���!�1�(��[���J�Q:�UB%��D9d�z��aj}*<�/��u�6��2톷�}�DRY��S�j}2�fU�X�/�M�q�(s��Tc�_�r�az��ɿ?��]~���]���s�9�M�mj�gC�'�M	����v�\+Ry�lӫ����/"E`���ǯ�q�b��[g�~:�Ѽ|2�2Mu&��y�u�W<�s�����mʸ
Q�i	��#�a�t��4ܮp����\��D?�������0���WOs����nβ�u��8qmC�_��nW=a��{��͍�9�jaÞa��	7�(`K����j���E�/r�k�q3��Eh�68L9���값�e�z5!0�7Ӟ�U����O��=�Jaz@H�Å�:��L+�<E��V@s*��{�{=�m^��Zw�&�K������IŅ��]%q|�����=(�E�-R� jm���f>UYa�/w�+˨�#L����s�ѱ5Ww;��ѠYN6�2~��]�4�Ѫ��`ڪ��^�L3�kX�Ϩ(f���x�bBX��|v�Z����ԭ��Y�xQoF\� �ET����Ut�rd%�?+#|����&� W�A�_�N��K7����4��^�2LX���Rtچ���a��u.�T��3~WB�c�l�k��9.I��ӓ醷�,�z�!�,z��a#r��{���i6���0�M�[�6�L�����X���c���6��v��H����8ER_݅�0�5A���i�}�P��-����Tְ�"ւd�H1�ʤ	�@�_3?=ʙq����`�K	s�gx�צ��*өY�*�%�����	kqj��%�8d㛶w�YW��uO����7i��g\���n4�x����7�y�����E��dˊĎ�Z�
�d1��e���F�rZ�N��V){M��n�~������~��!I����	��cG$�m#���,O�j��Զ��^?۳��>t�׺ny��j�������<P��\,�3X�l]Av�o������w�K����x=�U�~Z���O�aURݍ�]��W@��5�z?	hv�[;� 2���0;��������h˓ygw��l�:f���i���?��iԑS�֞�|��nYu����ؼ����9��.�;B�=��{��#w��l��A����W΢ns̤O���l��Ӏϴ� �*@������5L�͘]ڤWӼݿ��2�l���DTA�n�'�i��=���O�~�K&�R_+��ܽ�<*�J���O##_ޡF�%V�L����9a�{F;�����t�������p
��̷�g�M=�(s���i�k�$[�9�-�s���޿�G�zJ��n ��Yz_@G�q}c=��d���D6��}�>���ަ���N{�F�z��0�Gu�#O"~���Ks=����Mo0��t�fo�ʹ��z*�U�ƣQӬ��􅁝�v�~���2��oX|{m�{�G�D��2�o<�-^]D�?�q�2�w�aP�7r3pX�!2��^�
V9фb�%xxL�'��*����t��v6��&P��<X�eG����Ul�x�=��|��(�e�X��W�u���������&Ŏ0w�A�Y��0���D����L���MЮ���X�z�q��Td�)��C�H��E?tpHa�k���Q���
��$��4#��tLCjN�F��p���k�;Ŷ��#��ͱ�q��|H b�k2��_��V��-��6`g�t3\�u����,�q�Ӛ�f����f���^�$�ݦ�n;C�mm��,}�j3�f�����6m�m7;�_�׬'�:_=?�I�����^"r�g�A�iH�UN,�_]j.r��s���Sn6v��ٌ���w�I��j\wY	�Qx��-�tEI�_��T�O� p/섉����l$ː�zi��|L�0.�QO�;�2���
�n�1�{�cJ͇�u�IWU�q�� ;T�	wEf9vh,��Qw����6�y3^��()�n�XuO<ݸX8*��Ȳ���!D��-¸hf�m7�)��q�46�+���*�3�����rM�]T?ջ��(�p�9����@�֩qO�׊1EV$ۚ���n�3���~ o B�8����L��Ӟ��l�	t�U5(Z�����ʙ�fy��2�H���8�ӎ�Z��܆׼��`X�Y6�e�S$g:i�-�-4믞f���a�n��mޙ�e�J���
'D�j������M��9��[�3��K7�	(v ���r�?�S(�h`�a C�.�36��į�SUy5�J#�>u��4c�e�"��VM3�l8��'����Fna����g޵�k:�Qӣ$4��1n6�øď�&���$�
�KMK���*��y�Y.�fU_��Q4Dh�l�q�WF�яol�;]:������xN��6B����V�.�zv��I�)	2Y~��l�?���1Ľ$�1b	�V�|c»1	3���L'���>�e���;��} ��Z�X���\.ͯ<K���Ͼ���,Ö+o���ڇ7�7��F�i��=�5���V�M`�/��W@�n��+�J�0*�UO?�M�C�C��/_�?)�e�Mez7�g�,�nqu���ߦ�_�������uw
�����Ջ=馞��D���,QVt���u0��:��I�gx�2L/==Q�^�U�d���k�s���w��W�^���:@��>��������,�x>�������W��=v-�Ҝ�H$Ю��T��n�})Ag�A�#T�g7 �f��;��Yw�A$FS��=�n�W����4#�.�^"{�4�����K�g��Tփ/�a@�{�O�f���Q��mq'��5t�0ӱQٞ	�-����i�/˄~��U1�tW�I�-���ԍ���gߔ����b��Ec<��}sbj�����0�N-���q(*KwTZ t��W�h�[���Ġ����z��O�q�_?�2�l�A�tϴ�[s��b�����kˮ�/���ɊDZ����]y]hD��mm|Y�ɰ��W�.����5��a�M��+�U���8��Y�{?7�΅�?�Fn6r��l��s��f��=lx��wSY/do� ���e�l� L��f�oU�{��V����8Mok�k�8:'Rg�6O�e~鿗^�!��j��d�uJ
�S{4tJ?
����� Z��1�ƿ��G���\ȴ���0�eu�U��G[~��5�>�[{��8��Un���,����"ޕr�_3�W����'O�����������to�Ѡ�B��=+�]�� �� ��4jO��[�q2��3?�f���洧�q��;����1���#�e���龛��o�i�w��nY�����-w�@���rKLZXePØ��*a�s��3~�.˓q�˯�O'㙗��i����f�ϝ;�̾w�����	��kE��k��
|�!� w0m���+IY��-x*+$���<Zq�3^\���t3ͭj�����3��gg��������j�u��#Ы��8����֫Ъ������QM6Ds�	s���u"� �T�N��{�Y��Ȭ{�k��W�����0�����ޱ.�^��4�|jiq�WW���^����=����>=�������{��Y��da�SY��J�_�מH�9��f�V�٪������3�v��~����2L��|�<&��S�i������-|�g�A=����5*��*�}�$�L�6���Dp�2n�SOx���L;�d:�J�ZV�<���'s��WVxY�(���6�yw�x �n�0�����;l�w��D�2nV����;�H�;������Z��&+Q��i'@Ե[�l����8��k�e��lt�i6|�O�uw�A��6�f�QO�O��=�S*�Ր����+O�k�]�Z���&�֎�g{�j��$�l9U�%^��캙��l\�х�W7\�Q_�H{���	s�Y�����[�M?e��؋�'M�����&��ݕ-�7rS#A6����}��\qW;(�����l�[D��$��,�.z�1,_V8�i�_�|�_���5�[�zz����"z�g�5t?����k�w�oöf�ߦߖ!��:�~��b��2d<�7�[�M{�e8�������l�}�B�ޓN�G)�hutz�����n��ۺ�
�`[=t�3o?��s�7�ή��sQ���~Y!����$�}��[ȶ���Z.g߬�ƞ�[��Q�[,w���}�[��j�v�JiDlU�=�E�گ�T����|}����i��km���-��]�i�!U�n�|!5��ȓ<�$x��"6{7�v��*���?w�S�Q�-B{@AQ�����f�x\b���)�t�7�Flg뎱aʓ���Eks��{K��BZI�Ys[�Y��E��2N��፟ȩ�ٯ��m~�� �a3�ަ�_k�<�]=�����=��� �_�u�uk�3n�հ"o *��H���4U�f�¡��u�Z?���7h�=<����|�e�2��m?�p���f��m���2�]�}#w��:�.��Ӏg.��*���r����0{���/+�{=S\�kz-u��ߡ�ׄ�� �5�ifGJ��?�ճ�GW�S"�OC�~Y]��sF��Ou�;jOe�_��q-C���h^R��"Y�$!�w�jm�ȓcWEǀ���`��0E�!BZTR�FV�<�=ͻ�����~�nʷU�J�ئ#�����Qݻʹ��ܼ����ZX^"Sa0�M�����ّ��M���۝T�I}0��(b6�'Rd��W*Py�;���|�o�t��Ӟ髧�z�k��kn�kӕ@��#ߎ�h�3����=t�&
G���Mwqƻ�Q[����q�K\I?uݼP%��Yx�:̼ⱉ��5�q��-����w�����=�ek�{}��5�E�+�K�LQBB'��T�b��    IDAT��W��)J�t��a��=���6?X	�^>]<ä��&��_��i�#��8�9/�7L�aڸ�1g�g��UڝhQ�0;x��7���a�b��q���e�v��j~�
)�69�ۺf9uKs�5J�u�C���ԭ��7�*5�=�@r_���<Y����� 2��O~�|�����!d�M.����u�;���� AQ;z`e����ʳL.��ig>�i�u�<3�z���n�{�=U��v�6��}?��13�uK�L��$�fy�rf�W����</�n�ӭ+,�=�=�gҬ����n�+��B�@m�V�i�I�7[�\;Zys-�t�FW�3�L�يe��̳"��=mȦ�w�� ��d�=��2�LW�H�yj�<#\�-�,���E�T7b��bχt��#巜���s��o8cd����Ġ�,��R��*#:�mq߉&K�Of�6��^8�~�Qe��}h��ݩ �#_k{�L!��ʔ�)e��ŝ�H�E�M;^G���ޱn�*�h��Ӱ�	��?w����V�G��g�c<���EI\b4:��L�K8R��g��ݥnsParb�[1��Z�������A$��U{ �^��'�5�t�-���8*��LO��m�̣�����3�;�J����S�3H�߽}�3M�����Z�#,���_s�1ӌ<��+P�z�I�H���!<1X��b�~v��|��-ի���9�n��;������1J�����Nv϶�fE+8'�@EW��uo�����=U�����=-wԓ���Y����y�n6��=���[�ߍL4�v�z�g����n�NSߌ�.��&G:�~��~�m:m��%�h���sϸ������[�iʘ����I8݈w�m*����L/�;�u��}gg.&�y�6���[��u��-c�ݔ�6�)d�Փ�nF]e�l�Aզi�L#�����<N{���n��,�ni[�TmY�m�8�e��O=㥮{~�z��7˒a���ކ�p����n���f�Գùx�{�B<�kO�K+�vK�u�7�f�,���
-�@^Y�M��`Da�{3�Gg��ߠ�J��e:��ֆ��9Û^旺n��n�{k6ܗ������gڷw���zp��x�յ@��n���.p6zv+�vsҚDG�b\�F�^ڤ��qSE=;Xf����'��Ӎ���CA��e�fK��KoY������U�������p{�w8��E܆���`��˟�r�z�M�
��n�m�*���	����i����2�Aw�;���պe�>�_L^6�z��i�g��~�M�dz�iΰ�[��F�z.��z��{�sl��(
\�ۋ/"�^�b�G=��G���l�ѣ �C<:*��3|l�,��\�"�*$��z�`�X���7��x�q���5L�֚�8m�m�/�l'6��2=���񮤢�u�ޖ+�Gܻ�؆������-�H�{�5�6ˮ�O�yd��=�Ͱ�u3|ύb�(�̸���'N�oO"\���I\q������:�k8��/���,������
���a'$^Gfa��<Se�'`�-èO�a4���n�t�4RL?�gx�v�F�KUm��&-�[�^�;�i�i��:�W�5�o/m<��0J�D����<������"ͮ���[�#���q�r4�a�<nܨ+��}�˼�y��>=��=<���-�l��. �������1��mʱ��@j�WP���w�~-r�/+��L�Y�4'�ɰ��f�m�~m���p��J{�մ�qSe>��Ꙗ�6�iti��ƕ27YGr�g���tul�O��[����]{}��Բꖓ��]���~v�]?���&i��7y�t��m��w.aڙ���'�3�n�;�����
��#�w�l���g�l	p��J]��zAO��f�� Q��ůV�/U�-�f�VY�T�P�3|����7�N�_�q5g|��9�͸�e�2��K�0�t7M��k�2\�����`m�����o�hnå�n'��kuˬ�1^��a#�9����X>�M��/n���=.6�"�8z(Q"'�۩,��9sWܽk��2׍L��e�d�FdFq��fȹ-[�z���]�X�p�,��Qw�*�����ӿ#i�m���2�id�hT�����|0f�W�Q�Y�^i�ѽ'�Q��t�e�p�QJ?�CM%�u��xY�t�Mw[���W:�|5e��{���OЌ�z��G��=ӳ�!m�k������"t}[�����k�q�[fW�C�܎E>�ޟ��*��Nպ�Ӭ_��ά_����=��O�i�kW�g�p�~�=�w)�H��R��}��F�rd�3��gg���ʶ#���D�����L�g2�G��+4�����0k<���ӽ ���O���D9��rAG�ۓ8�F��~w��M�y�A����K��6��Q��݁�V`d%�0VZ5<��g�3G{-�&u�MՆ�M{���n~�iؓ�*�ɖ3�o���~F�>�^c�{��i��M�L����'z������4Y�V7���Q���42^��h�n�4z�3���Twۢ�����ק�y1-ٓ���a^;H�f����FnX� �vS�h��?�k�kX�Y ��~[)����m��j����id2�`z��N�_v�to�[��t�\9,��_��q�4�U���j�Y��ph�N�֭5g�t2�z�k"��;�x?�3G"^�P�|ϴ񏉦q�s�fN$��m�m쒾��o���2 �L��`S�*�ʡX�D���pP�D{��=�5n��j7��~�3�t�3�tO��z�%�ʔz��x�z/�@����3�i�{��@:�q�+�n��-�3ʹ�H�[�4�f���fôj0\����a��+-a��%�HBҦ=�;�����b�T����\RY7�D��������������uvj�r�����:{Q"wL$1Ǎ��f��J�f�iO�hn��9������z�@&ͦ�*�2^��a�r2�f��z���ץ�i[�Vq��gm�i�����2�F�c��/�Id8�/�Ro��*����ZQ�t�,G�A��a�H�t���(o'H�?�TE���p}M��Uԉ�׷���?�FnVע��1[��f_�D��l%��d�2��,��7��Jd�Z�K���6�u�������܌�j�~9F�� \�z�x���ȇ��꣓����i�X�t�Uδ���a�׏��{2?�T��nm�Z����F��bF<��Ong^'�+oRw����6�ʜ={o���	&FK����Y
V��ʒǧ&gx�Έ���1*a���2`vTwx�A}-���2?�TO��t�J��H��3���;Xh8��f@��Xh�$��<��Ꞅ�x�c����:g�U:[U��^���"m��(ʟ{҇�q�$i�ӮDV��7yP�Gj�sNhp��/ab�=&���IbO�o�n��gE���ߠ��>��-_z Be���򧍓���=�$d(5�H�ig&�˸�Ty9�f����9_QN��k �P��3(�\[Y.ss3e��R��ˋ��G�����́�X.^'��|˷�?�_���
B{�(8>�$�ն������/���g��BL����"��yx@�R�N�\MI��܊"�e�N�^�.�:RĦ�zv$�]런�#��.�U-�zp��R��_;��٪^x5�w����Ӊ0]�v���#�|)r5�l���8}�5\~g"�b����G+
eST�'�VWI�SUJC�p�@
���HD* )�x� ���� vT������c��'�b�d�
o�;J������Җ�$�v��\��y�^N�{��ݟ��r����Ʒ���Z�g���ۙ��賵�X�\}��M��H[�?C������~�7���;��<��3��C���%�����"8��6"Ј��DT@���P��H�b����L��4-B;B�
�Jd.��G���X��[=��ꔐ��#3�4(�%(��a�_J[A\̹�p=FDPj����H���r}/EXB]6��xfud��E�j��G�x�2UT��X�A��7��n6z�3N{�~f����޵1���W�W�B{�ڣN33�m�J98;Wn޸�9U�\^ �7���گ.����<��7��Rϡ½-Q�'?��e� �mh�^�+C������,��
^���[������ce�ȁ�|���?���W�cÕ�1oG�d�qU��傲p������:�fWg�1�޵%�G� }�g��lͫg¹�h�F7L�ӯ��!�~]v�e��#ZO5�^��S���w_�ϫ()9v�X���ꐭ����`�7r��e�Ҏ���C��#��7͂����S@:+�[y�k+�@ɰi���q�EH�D��=M^C-�ٱ7��9�������R�n)0/_�P&aU�a�W�ڟ/G�,���@�Q(�X����z�*� \-˜�C�A���g׸`���h��5̲7 �ƭ����{�3��w������r��8��d�yG�/�o�*e9G@~_;Du ����o��� {e�R�@�h&�����'�G�5���7m�O�F���_m�l�q�)�!��1���F��N��B�l��������\�w'}_����������$������G�`$�L�F�2���-��#���h�
0+�{ �:� �v�!|�����>׹���ި�5�y���s�9��Ux���J�k�W
Ѓ績k�|�w��������׃��v�
H3�q�	�h9r��L"���%�����8_&� 7�Q�����́p�E?u�^�|
~��B���J6�*����4�NԵ�@�pՁs,���z
gU�b���֝�f݅M��]2�����_d�D���i��e��-ä.��ٷ�5���_~�r��щC�N�6+���=:>�q=��9�l��y#ޥ��y��Y���n�VJ-"��2\�����}*�q�*�@�|)�ʗnu�[D�0ye��0It�͛ 0�~�W~e����r�� �+\�?_�^�ä�~yy�LN�����ū���	�ݙ�aX�_�l��
H�y�3X�i؏�7.�q���^)K7��[<lt��da?|����{cR\�+���X),�p����p�}�jV���]������Cs�^=үI�~��ԺB��Ʃ�4�Î�e4�NI8Uۖ�v �;q�D��U�2�i��H�2� �wQ���/���wY��q���o@�W��V-)��[� DB�.�Jo)PV�F��dD�g8�2l�Y"�@k�䷕��_K�"��[����_*����ჇA��r`�`y�����q�M.i��ˡ�sP��6�a�౫:�/߲�K$¼��Z��)K�܌nL0�X}���t��\�l��ó����ꤏ�����e�NW[�"P Q :YH�QN��ȦN�D��	�M�
�|;'U�*탰�=ag��+͉�3R�'�[�^(Kg0_��{��c�VWE�*�
mż|�Z�����ͯ�X�����7֜Q�ܾ�><�-�D �t\j��������k�ʉl�J����D����#eowUk��,���QB�%[Q��>6֟������[ʛ����	w!�'U�2�E���;EF%¾, ��ZE��X�>�V�ɩq�?T���4(�fsk	^���n0�^.�`T���T���(������J�VaM��� G�B���+eb��:���L��ӫ�k�^�� `����#�^�nP�32`�|y����R�P�	�w�{;n�)�1jG�B�)Ͱ��+ݮ�M�]dh�ɱ؆B۫-��rk���~�j���'w���}/�/�]ʷ�l���^�5�j"����* ���q�̊Z)�KU&��>��Ͱ��d�Z��5|� ����N�$�ȑ#�sD	9�,�d,��������<W����,��+י��bbe�7���2A�SIDuK�e>zll�k X����v/��$�-�X:̱=<�F<�G>;�oxd�,�|���C����W*7�/��).��^�%�����Ab�$�� �R�	���K�΅�=��������O�M�����m�,��(}�x	�l?��	�#/�vݢ�;��a"@'����o�Éz� 6�nӔ����	=���Lp}_�}������u�n3���8�r+G����iq��ʷe�0�%b'�w�%�N��_��]�"�i~)��q�A)ȱcG�&qR����K��`�u_����Ώ� �*��X*d�1���< ��fw�1�ff�=�,�CJ7_+�P���_����cz�S%���\ER�� K���,��vbb::���f��*z��Dy��3���.��(߶����Vοr��Xܠ� -�.���9ne�E��x �λBgr@I>��6G)�U�_��#�}5ؑJ�T?�;��4���ILG��໵�YK�	�1T��<R�9Gn���m�.��U>��v���ܣ�ܨ�bi�.-l�,��������e�,`���+ ��'�&�G�L =�t��;�2h����b���PaYCj�p��bʷ}۷����{���O���z�I�*7v�ƅ� �K�  �敠֛KP�eq�2io�C#1Y�	o�L\����,ȸ84�����3����k��.W�!����]"��x��2[<^>���r�)�p�K�{(�ty��O�����Ay�%��	D�W��,Ӂ&�8Kt4���I��� K�D6F�4����p�3L~&(r�%�U6ݴ�T�q���Q�j�I�쬟��B9s�yF�ҥ�V�B�6�%���T�zcD���~7�xR����;����5��m����Hs���ƌx�V��~����0�����wѝ����}wy����C�'�]���ϰ�a�.�27;Ų;T1����-X	d��S��˅K@d�h�B�^,�K���k��LM��	5�Z9vN�'�2Y����30cS���	�1�
�W
���������˗��O-�_\�,o|���#?�����?\~闞$}�X;������M�׿��
�p�e��]�1��ا�����=H��P����v�&��4�t����6��{/��jbb$ؓ�����c�������;��ω�R����5�غo᰿�E��Z�� �պ��
��h��WO������ęu�y�zH8(+���޾���|���E�9� �6����|q�I��R�m&��K��U�����}��O,�l<�LM�Drb	ȑqyB��$4
��Mf���,)S��U`���H9��e�ztd�:2�y�tf���rz{�{˵��'˥k����ϗ�O�����~�)��{ϗ��?_�|��r��[�|>d�#�[g ԃ�bP�@�mR���RdV	����?�t�v��to�N�ȡ'çn���/:�fG`�\�9~��Ёٙ�龗ڽK����"���6��GJ��F�xR-�8+�%
��v�|\_�d�������^�5�F~�b�.J�=��"�
��р��n!~��^`�������o��߈�׮]e�u%�k]A\a�bhg'��B��SS6�|y��ϗ����@��P�u���ˡ[�c�����/�O��2;��n���V��C��3� �#�����K�0l�ְ��B����ÓX��?�X.^�h�F^�j9��d���PN�:Px�x���|-���)��jm��I^o���<�TVJˊ�C.�+��K8���O�JJ�07��F�N��btP�^۴v��sd{ն��:e9��ٮ.�u�p۫�o}+,���q������=]jw��Ŗ�]��9�$�r��=%��\[c���*H� !nx�^�V�Ъ�c{fcO~2��4�:H6��-[��tӬLԕ�{�9�$�����������A�X��K��^�>Ϟ��@�nݼP.n�օ��z�A<�ݤ?��>�b���mxk�q.E�j*C�Bg��iD
���Q�Q��%�5�F�xG�D��sK!�^����F <bL'�k[A��M�-�_x��tu�����v�E��嫿�]�G~������b���v(��P16H$L�������4'��`<����@���v5|�W�$�팧ҽ3�8��O���1��/����O?�4���&DV-.$l�    IDAT7�Qw��Bn��!����6�׷��s{)��8����%� ����Nܤ]#s^I��w� +@ԿҲD��<��I6yE��[dB#*�0������|�W�BT�P��Ef�B^�$�}쭏��}�/S�C��rm�O�[\�R�ͯm\�dM`?��k�W���4���H����Z k��3T�m��^+�ť 9�_�ޡ�%S��L[�md��/ D�Ed���|��	��&c~����jϢ�y�b�
s�f�<�j��_|��9�@y��)/�|�|�w~My����G>�I�����h��r�nHV��I�Wa���"Q$�� �A��h�!��/ʁ���eG��l����0�v�hGe�T5C �-L�9U	L,L5!� ��Y�gy�u�,o`!i�w0�{����)�V)����{����x߀2�Z�Ae�+@�Lu3�a��HѦ��җ���"�R����d	��;����W�ǿ\���7�^���<�����Di��IDv�`]���\������TtrJ�(֣��O��D�I\�2�j)�TR�ӱ���p:�Fa��E� �,;WC�`ǕOg�`�Ō��4�PpxP|@=Ţ��`��W~�V=	>5�uc婧?K�b��C��B����=R~�_�kF�U:�WaGY�B��(����Ŭ�*�M��������n����Źb{�v�i�������ؐ�z�¤Y='���#���xrr����ȹ����l�r�=��мڕ~ƦG��:$g��Z�@�[��_tW�p��pȬ���6�65�(���I>�}�(��Y���������+ސ����(tc�=�P�!�|�������XLaG�6K��K���@Mi�\����mv����bI�JLR4�Qc�� �e��ENp�ӄi��CL0ch��[��~@�qS�����(�<����a�S<��j��	�㾧<��2��������b�|�����n��-,��Ú��P�#���[��&�3$n�iɭ94�խ�TY,���Tݶ�.Zk�^�t	q���[�u�vM�	Oɢ!��ms˦���go�/����B3~J���ۊ�ږr+��u �9U�ڳ����Tm���N 0� �z�F�ڊ���1{�,�C�>���'�xQH͖It��H9�#�^�Zo,/]`���<?0 �+�L#�'�v���7��3�dug���iT�,ӆ�8��Hi��r{�4�> 9�:t��A��!6������ �=Ӭr��3�З����3��3���}��{���CgCl69����+�����}nn��c2d�9��v@$O
CD.1��N�8�Dp�+��K���l�A����3�4�ܵ�\���M�Cح��.j_�m�ԁ&�˭�e�-����.��Bν�[������+�� ��B�X5h�תL'(�'�M�ೕ�L��</��	�x���]����!b�q�z�7aC�K+,��h�[�_)����ي���r-�C(#�U��.���1��T4� �e	��[Az(R�.����\�R]`E�.��4H��q�E7y�j�+��A��l�f;�Y�|�ۊ��cL�op>�$�>T�y�Y��\�?���ןe$�����|�ϰ�q����Cl����Z+���V-azM5ipy�:_�A�{R�����5>�̿l�a�)�S��N�$_dv$"��!N�C�&�Vc�s����c��L�븳���履�[��kkt*�?P�A��Y��l�Y�;�m���G
�)�×�u��={_9{�Y��c���D}���[�!�[������^ ٖ
s�r�� �Jt��a^�`�]�`�%V���n�YCN�T
�������]��9(�Q�8yb�r��lh� ����q���g]�f�<�@��Nv�z�_D�93�\v�i�V�)�jy�u���˧>����������{��]��O�83ð)�#�&:L�6	�
�7H�c1P��S�Vm��aj�D�Ԡ=�S��6V��e9c��+��`rw}_�mRtFI�⿡���IVo�T�� k����*K���	���H��2�n��6%����
�c� ��~�`�{������C_em���|���ɣ����x����]-Ǐ��� �A^�^Y�H�r<�emyj�r_�����&���A�`��g��J#�&��Ll�E�>?|�<�0����l�9��d&a��H+�;��/U��}Q�1)�n����r�=����R�EʽȹN�K�^~�W~�E��r�����g�/�FD�u��1��G
U�O	��	e�~�)�A�У�$���� ~v��U5��K�V;9 [��&�@I`�V�bK6f��N2A�z0��j�����2T�;�(Ȗ��ٹ�J��Wi�a/e�2n@7�v�A�o^{7�n���m��w��]��q���ny��s�M��͛��~]d���ؔ�ؓ�����Ԙ}%"�Ag����xk��D�Q/��	����@��5 - "�<�,!�'�0;O�2�2���Wʺ���A�Aٙ��\��b��F�D�׺���;�?�����'O���y�N�	������g��\���O�/{�1ح�����l������BS�6"J�P�%��0���ٹ�[\/���h�ʥ_�U��/�Q����OGm�%y?�q=���V`wvNLL���
��j?�=�6��6>��uxt�R�b�ZY�1�L�����iΊJ�����_]d ���gxӏs�l��a���a�+��?��7�7�K�.���W��D3l�f+L��6�巼|��K[�� 0+�na-HP�An��A
��v˪�j��ǐT�pCl��)����J�n˜f�7G�9D}-����H��������zZv�1S�*�X�5c.�PQ�/<:ʊ&,#�>�F�*��:
W)'˛�t�|^�{U�?��)���}����);{�)���F��8Ƥ��������d8yn�t�m���*[8&ǘlW)m���VEےL?�>q�6O3�ڎ��z#����ro�d�2!H�7�˽>19�@��[2BK�l �Df+����T@�tϲ�=�t��i� 5�圣���ه�._�o��U'�L8���q�E�tj�ʱ�ocY�ɛ[W9�H'�7P��e��|TJ-eID�M('����[ 7�?1q�L�jx��Q����9���|�uB�Ȧ���4��h'"q�l���G�iE���0�\2��Od�����l���&�+�`���3�:u� ��O���K�g˻������?^>��%��
�?�.���#�u"������L۔Q�"H��"L��8�X�g�<�;d'�h��,!���숬�5��?]�1+���Ʃ�W�F�U�U�c�[_[�➍z�����È���,�3s C��9j���z��k/'�256?��ᡃ�����?��������Œ�R MI���H��1�ZE|6��P�FL��s����2�]O�ț���~%�0%��h :.,�v�!�&�P�9���a�Ρ����|�o\"�u�27�-r��$�I��ᝡہ\�h�\	�"� 4�p�rJ夤"�R!E��`;:���Y����p�C�3�����#�R������Hy��G����-��g˯���('��|� �#�#�l�+�9w�lO���C��\�T���Iwu�@"������ҏ��Re���4�𖧆�hB��Ǧ�/��?���e��*e�d�}��%Ûc�l]\ZdQgh��tH-X4J�:[ɬx">5��GEDvT�	�~�|4�p�p� �,�z�;��w�}����G�S,\�����?8;�􁳍����!6(�k�8R�^������HVDn��lَ*�ˋo������,[��{7�/�l~��+PQO�ߢqq�L�4��9 �@9��v)�&���v�<e	lt	��nd�"�Hb'=��D�ƗU[^�IǞ���eo���R9{��r���m_>\>����t\&ǫ�����_G:$$�rұ,�Lě��S"o����v�uwس9EX)w}"����ϭ���2�(��Gۻiz\�y��7��^f�X\��� o ʑLɟT�r�����Rɯ�H*U�X��J$�J%)W�"�P�%�e�%SV��bDi;I(�@"@ �%,vg/��s��f�<���}=�~3+���y�~߾��ӧO�>�M��^/�v�l�;����N�ug�;.�C�=�<rnfn
V���2�`>,+oq|���o�S��is Lt ����fD��}za!V�V�n6O�	��Y����[�h#�&�y�[�]��<�6C�G) P��w�GG<�*2�=��x���恊Р�O�@�r"�}LdQQu���@(�@�J����[h 2A�Go��6(T$�8Ÿ��9׮�-��!��<��F֜��*r���Pa��%��ҽ2tO�t�?`	R���5(<�O�m��������	;�|��OQ�s��=Ӽ���L!�调�0l�_;�4�N�{9eU6�N�&�r��A�Ei�il۳t����=	�,�����ᅭ��y�fL*��g�[7�&�ve(�>r7�m����oݞ��_�=y��=o@�1H9kﻣ"�X{ؓZ���Q��}2�^��ȓ��F�?��⥋ͯ����7�-���D�}%�����NN�Dd�-a��6,ɶ,|�{Qw=�z(�,�|-lX���EU($ϼ���-��[��a�#���\4�����8���
����.�Pw��N�ha��Q��6�ґ}:��OE��҈�R��J�Ο?����u&��P�]nn߼QXf�r�?����^C��B��<�#TN$�X��uځl�X��Du�~�v~k#�滶�8n�H�L'ڟ�E�dh�IVlmK;��R�c3�<G�c!�����ѱ���	xl7q�"(�h�v
$���D�9���`�2L0� N�6�x6�1����ͩ3�l���|�cO7�}�2�bV�6���{�E}�j��M(8�W��(��E�Z^{���Ԏ��!���@�eA��	�ڃ@�!\�)�r9�t�?'�P�-v��A��;�Zw�GAN�[	�7uDh*��@��HKG�C�$�K�и���<���vXҢ�v�P�%ٛ1�?yd�fd١,7o�`)�BP�˗?м��nsE�S�G�� ]�����Oތ �UF���Wʺb���SW�;���*oψU�r��,:(u��P�@X����~�X���";la(��#ͱ�����橱����m<������v-"V�X�w�8)p �J� �t	�� �~��,t�8����왳h�-�󆼝�a�r�Qf�U�����/��x��2������Y\hΜ>	�w�!_k�o.d�SdJ��)�cL��/�%#��l��~���8�A)��.��qO�����K�]�Q��r�4)
�v4��è�dމ�������K�c�騒���,�ad��],�.4o��Լ��+4��|ꙟ@\�d����`�9�C�k�N��v�T�إp��X?M�����^��s{�eJ��[8��H\�3���<Ta��{RW����0�Bp�]Wwzjj�=��r{�ܹS�� r�bpϸ.�R8�,���r�n��}מ��]�H��t[ʪ�H-��N[����� �V!�qa+XB���H��,γ�`��.��;�B	I^]Ʉ�>�urj�F8�t6�~��`�%��f����; �c��P�R'T\���F79�O��&�j ���K��t��u�CV����+O����� �n�����:���������&@��S�2k��.�9����=�D��}��?��\�4È�X��g�h���w`=v��'O7�,,�09��pb@�\��{ �m�[>M�A!FR|�=Qd(�3�H�J����㢻�p�3&���i(�v�8u�D�ХL�K���s+.X�#��� � s,�F]��eK0F8Df����3g�R��8[�اPD7VD���"V,�
�����6�t�h���z ���~�s���.E e�#�@�[��i"� *�Y �P%�(ťLPKQF���(ϩtF^��E���s�߆�B��6*S��vq�C)Ï��l�*utW��9�;�T� :�?� ���v"(7��23
8y �B4��x�?i���n��eP"۲ƙ*� ?����ls�6#�D��gcʹU
1���5�T����=��o�y�Hem���2;'��3�5Ri;��̢���s���T��⋝Ev��#��t�g��Q5:Jav�)>α��H2�,#��q!5�EX+��n.jԀ���E�|7��J��|+�8щa�s��_�p���[��� ����w�fc�V�`I�*�i����9���4>��{�ܹ�w��|b|�Oā�kk���e�1#���AY)����Dh��"�R�Clޣ��bv��<�vG�<�n�ߋ�Zg���OJ	B0B!���F�d��S$'t
�-�-/��Ɏx�2�_��:2�A��ANB-���6�Bn�����D\��2�n����.�?��E�9@l�[7��G��$x��ӟ�bt����DsJ�����@@�h�� âǖM�D�a�>(C�=R�3bL�����6 �N� ��&=M�~7��{��C�C�2^�� ���ab��U��,�#�6�?3�s׍TT���A�">*�p	�G������˾� *,M1�3��B�-�JKm�jzuR�P)4y���a�SyT����OY��Ő&~�0mt�B-V+	�>��&:s�@�6v�F[��03�����2Ɗ�"G1{.�;�pz���a����˨K;ʘ�dގn����h�Kw�i���u1}�vd�7p�#v@�}�+I�m�ӧXu�И�ixD6��:�.t�+]��Q<"���6(n�"������X +��P��6��ɰ��nCGÙfĜA}�s��|��*��y;,r�*ɀ=��4�i��md��6�G��eؖ�s�
�����	��ὧ�NCV�:�/*$M�3]<�`X�`�����*�pQ,[��ٜ�Dը�ҋ����T�z�伌1Z���Pa�O�Ex~�:A˦�iB��N�B���O]H����	��zz�6_�o8�������Ia���Ňn�����z�6eW��ZPT�m�)
ʻe��R$�)a�5~lߚI�m8�}l/������(Εr{�T��4��A=����@ü���,3�2�x������z�-U#�h�~����)ݲ���t3��O���5?��?��;ɋ�L��Q{��Zmבּw=&R�`qup�����BcE�@n5����O���a9"ɶTY��O~ԣ��aQT��p����ގIY��A	��^� �E|'� �!���E�^PVQ>\ � �[�-�CG�I)��0��>�(JWv\�"�^;�����7�L�u�F|��ð%�1t;�&a#,��'
T�DhB�����[�M\H�D|�h��=�Ay�˗/3�,2��'�Rn���Ly�١8|,ʽ�>�a�/z.Ƚ��||{k�}���VB"t��pZ�Z�M��=�Ha	��1��=�я6���3���po����!��q�0�Yą[��LaK@n�;(x�0�LT�%���F��&��p���d�jN�jr�4$����u�=�L5���!m��=ؔ�oa�L���f�!l{b�8N�4�$���AVo<i�g*O�\�4"�=Ԓ%7O{����T�=�y��ع8{�Dsay���'�bQ�*�֐�й��`�P-���c.Qnʐ&�F�5�1N�ܸ%���p���Ύ��,��jwr�B�*���kK%#��?�b�����ʕG׸:a�.JJ ��ʘ���!�d}a�7+X��˂g�� �vI��[��E?���Φ��=�� Ԁv�O�=F�@L�V�3��'���|�q�ײ&n����h�}A�2��RM�_(f���ڥN"l��#xr���8%2X�B��g.�qi�z�8*��:���u/�mGa~����>ق��#!'VT��7���    IDAT9x���K������M1�I�-ymD��n�Kh�(5uOc[�ư��2���m� �ߺ�"̌��ȗ�x�)��I�]�4�ys���y_���X���o�fj�H��:�a�S��<U�J��B5��wZ��~�kچ�=�����&z�N�
�����;6J ]�ۨ�2�;�t��L�c��<�F[R
 ]��e2ʉ�q�$C ��;\T�E���M'��|�GD��	�=�b:r�m(,��e]��',
rZou��� I�~G�5��Ae<�O.,�)����Uiy�g�i�M�!���z����x^�t�#���QYF��KY�;eK�l#˒����1�������^�o�gZ޶��Y7ꃈ�+�D��0r_C����'-�3[�Sc-g��mc��V+���~[�4~�O�k..�=�I�0��;4���[���"�ڠLJ2Ȟƴ��\[�6Y�ʨ{Z�}�+�U�rƱg����l��.��ij��p��#�?���~[?��~<��'UV]�j�PR4a��8�#��^`���I+�tT#M[Xy��>R�M����L,�)�?
ז'��:d���:�n���5��ER��M����zDgD&�l��<�k	�����<�<{�9�=3) �#3���,C(�`ȑ��VW�B;�/��O�uO�����/C|� ��p|psn�c���m�ڣ,�xb��r'R��,b��%U��5:�*&��o&�ml���{f*�r�ȼBtt�Q{�eѨ+eS��kaUJ}�uһԡ�V��
��>11�[W�(����&y2�
�7�q�t� xAf�&�]�,��}<�@��}v� f�]:3������Y������v;���y}s�;2]�үg��L�{�m�4ٞ��������P������N
�������H��:���%ix�,GЍ�G��4�Bn�t�愸=A@�Y!&/#]�
�,t��<U]�Ұ}D��LKMy�%D� A�)�`'��"r����P蕣4'gV����PrM�#�m$J&F�S��S,��̜�@˳(d-�S�kL:�,�;��G�2�B�H�%{ߖ��c;|�V�b��u�*�)	釭\^�{S'�Kǌ�pTsN�,�|P7�dY�6ʄR��T�<\CSD�mh�&u���< �|9�`ƝF��sQ�(T��z��z����dq�T��{n�.�D���rQnY.�ua�j���Q��#|-�I<��H!�g�Q�oJ��Wu��"�aE�%\+������sS������N���9�do��̈�R�N����V���!�4�+����)ZS�E��{O�����sT���_RBJP!�g墦C��v�����Ѣ�Q~$�PxE}�ϲ���;�<�Bю+s ���X���u���:$(G �Ҵ�@9�{HQ<L�%��1�D�w���	�|M��`"����@�"�rq^��e"��\���$"7Α���)���Xp�����QӨ�$05�ƚ���1���n%���~�"��iҶ�GX;���+�&��:k��Y?�%8"��*{Gy�6��^h6��]���O?=�ۯ���"�˟c!7WS�[2�}@���B�Jz�����i���-i�pk�@Y�LC�E�mz��9�m�p�#�;��3�2��aC^JN��#P����q�O��T�CJ��#� E�!�pw̔��"|�˚+E���Do󑅂eb�9MS��Š���14+�Sƾɉ��}�Z���a�-,*�R4�I~����P�KU�ԓQ�i��M8����|�Evق�U�H!���u5Cm����u+�y�W��(VJ?렟�6C�u7_�P�S`/2�	,��p�V�&*����oR����c!��佽3#s���Cd�H=)�����J�
�h�\|S��~�dX�h���ïMC�ՑHJ�[��I�����I!������*D�[�5�Q�g���[���>X��j:Ƭx���N�R��AS��o�u�����<�X�$�
,��P[Xm��.ۤ�C���=�x��
e�y���oE��Q*4+��z�����d�E(�4��U���İ�;I�����5$����k���MA�lӴ-�5��&�ֈ�Y6���
R��Z��6�z��s��!�
�;���f�>�÷�s,���Do�L)��܍��؈�3�JX1��0"��T*Qz�ˊf"�?M���$҄�m'b�p .�M&9�� P:w���X�	���
��~��D9�wNs�5Rs1�o���A�b�#�Px��{�_�?�%�6�L=��0ދfb���@H �H(�k<��� �;�И�2�r˺�aw�G�A�=�mD����g�=T�\��6�E.=���9�����l��fd픰d{i�)e��,�Ɖ�m/K"�Ѷ�0�/�/�Rw�g�0v<Ag��T�Q��{,�f�&fBU�C�������
[	�O��)�e�Yx���T�r�Y�"��fG |l�U�IF<�W�Q�/�����n��%��G�����>�;\h6o��ȵ�k�p�8�r������ԍ(��.T���^���ə�� ��l�l�=���-T_�,�tz��-=��хf����oI0�Y��E�ogvW;��ߜ�*�����68b:�s��&�ٯ�$���ɤR�Pz�Z�B�K�R��%�b"W�sK���l����7�.=r�(���"G����'Ȳ��v�A'���qwCQp� �Ny
���*�j�0�M�$<i�e�
���ò��o\%:��fݼpu};���3l=��'&f����[PL7��ds�C�~m�ե'��%�E��D��͆�,��] "P�l�b���qb����!l=	m�DD�:y�q6N�h�}�D�g�! ��t$@��b�v����<���GSD�w�#E٥��;�_�Z�؞L$��Id"�cg.X�1�(iy��:Y�tYv�DjY3B��<��wZ��'({8!3�[��H"��д���I'�(ID"�".�M���Em6�N�C�L��<M�a��,]y�E���tg����y}��Lr���&���E�BCxΨ}��X�mt��1i� Z\�����t�̙�K;��
P���2i�Dj�}Ԃ��	���`�]z�] �%��J��;1�q2�xC'�HFܛ(�(��e�<�[�3��w�|�!~�C�~:����O>�6��)��:�����!F�¦�.�
���"uA�9ڕ���Pg&�¬lE#qD��ә��\qRr��M�6����n-sG�s���s�����!?�B'$��0ѹ��"�,�ڞ�!��w��v���Q]	�#k��p-���k�k�vT;��Ȭ��[>��A4��{nl����׮\9�KA)5�B��ݭB"H�L	�����*�NlV��J�F�C���\R�(	?�����6���'��&�����
��^��<����g���yW�|��)��b��=�.�Ih3�����'mHW#�����b���3��ӡF<�RD��66�&(��'�D"~����וp�1���_9�av�֊F%M����G:R��d7�,����D#�(����i�u#%+JF�7g���tf��r�����Й���Ǣɏ޾��j�><�����b?�bY!�
g˒K�h+l�Dl��aie��ݶ��/r�#�������Q���eHdag���\��^j�OI���$�)YT �'��0�FK0�N!��"k~'⚉q}�$B���;�H/��˯��j�/|!�^�f2�Ss��z""�G�y��8�Ȩ�7���킐� �M�]���?�J��m�8��|�=�l^ �=p��86�Q�] +{IP9;��@O�-���䫿���HPxu��=PQ;��шJ.����5���t|�BD���tӌ̬c���G�	������$+bF�Ng++�a�pB�-[����ͼl�|t��iDn�4��[��,v.���(�q� �u�uaA��Cͱ(���l��V�B��,X*�y������N����H~[�D�H��"�)v���{F��k�Qh�YF9��s�8qT"�D��=���8S���)�G-Ȣ8y��/�{��.G>lnrq*[���\�.��c��J��a�INS�2q��TaH��,)�E=[���i@�bS^Ev¬P5�o%�iڐ"�1�4X�@���Q��d��zj�x���v:�2�Sd��F�&{�|9����qD�)�Sq XM9J�E2�v��ߦ+����iٹ,����� X�#�1�i�蚨#�n���`A�O�ώ}�k_�~����/�؈��9r �m34	4y��:����з-���!�F��H�F	�,���G?�߇Ø�@��.qè�\E��F��C�ú�����`�;��!;���skو�H���TEv����Z�6�o"i���5q��Uz{49�-.�4�(Ԛ�hv.Y�,AnǆB�ccBԫ��2��ǑN�y�ƵAE&^�.}���3��7�BI�O��Է���l�-f�4x�|.�p9ϑkȾ�޽��H��=:����w)��U�����m]�*�����m��A�����L��W4�Z�G��\{����k��&p�
16���3&�pO�~�������HN�ʕ��m�qXȾ_3V̂�XH��́��Ʊ!��&l_�#ņ���$C�p��B)ʕ}n�U��1N$���{��o����b����@!�^��}����1kc�l5c�,{�ANr��JL���z�c�b��%j�/4�����f8Ԓ2�J������FƳj�B�H�Y��]��$L���1��s����G�>K�
���z*��鹛H���<W}�ki�4W N�u�� }��Oe���HZ:UA#�t��<􏼈��mj�ac�t�.�~�&�J��8��QAB6�t��X�vwƾ��o_{��gK�tJ��=��	%����H�I�("ҩv6@ܸ6��2��*�"�5e�K�eŭP��$$Pt�I`�@Я �,�Hnh��v2�ϩ�7v�8ӈ��I�&�^i_�-,�,���'�4 �8ԛ=+���Nܰ���}+w�B�9��MlZ�ĭ
�̞k��c�">���1Z��f��Q�3:��1�$���]�h�.�s	_v�f���A���������߈''�&ᒰLb��l,#*��!,HR�Clr��:��:�
�r*�$lBBc�$[MR����]:�~u��w"r��m��d��w�X��zd݈�P�r� ��i^|����e"�},����l�&�J;�e�c52(ew�I���(��C��^j%�����wm+h:�.)+/�O�>��������i�uD�8c�qG�2�i��V9Ijǭe�"�T�]7Й�à�H��~�2W�^�֫�+n���[͐Rx{Y�l 'i8�m��'E�Y�a2��\���r�dNM{(=��)W������hٰeg��ԒNva�@#�[tB�E"M�D��C���Dh�3��hvd�<�b�;�]���]���e�ܾ�1�ʴ�Q) �?��K��!J���Y�L!����>�^MЖ�E�1M��%cD�n~H"%��K;4ǃ��]�EE�ߣ�Bo������=tg���St;�	�O��a&�J)I�`��/�3L �t��MW��'N�!��NL�q���DC�����p<YR��R�O�3�<y�@WDA\O�b��YĹ��A�Y��G��0�EZn\%z���	��q݌}���nP&�n��$'���<.��&ؘ֗���7���"���z�O���D|��'q�c8�-���xxO�݄(-��L��/\x�y��M�\o�{�&j�����{�`�m��n��m��eЮ��}X��K;�(�En����A����#w��<eD�Y� �������;*���4ul,��;�X�A�K��0�Ҕ�.}QwG��eNw� ;�=۳-�ω�îq��.���#����e{�r�� ��噳*�
���']&�JI�һh�)�i�YF���f%����t��L4; ��Z�8Go��������'�Cq���5;�z�7n�'�ބ䅎�un�ȭi��'l,O"xڲ5�s��"����4�#��D��
���0v��\��{7��Kw���*,���e�q�0���'�k��Þ ��&�L�RG����x�u�4Taʸ��-��>��yj0����ԩ� Pgd�ۍ�!�7�m(vQe'�T������~�#X�'�7���=�
q�e�k�{����/��x��AMX:?Ź�#�Om;�����C���A�\͖b�@�ゎ�x��=�_��1��v� Gc�$��l<�i~���܅'(�"��,��:/����K���-�t�����x��=q���S&�Ym�ʼ�Z٨B�^�����%�;B*ϟ[�0L�)�I8G	�Du�٠�S�����^��d,�V�zu;�%����01��k2ϴñuO�l����گ����:F����D���Q��L䎚u�RJ{�l	KڻF�
%:&E ��<�vR{�`��J�{�\)�yd��|� )��a=I��ׯ4��+���]?^��ȎA@�)�HƩ���)��EV�r�U�ˣ�CΞI/��\"�N����&��ҁ&Q�:s�C�Ň���с�&�=��N$�l�)vQ���E��J^�'4�lA4OA�A��)7T^�[&a��	�ω�:��c���(��-�ě�B��,�E���\��u�'$�� [�������g^i�-퀗0�ɶO��6n��t�}d7�ac1�bw��q�;x3�I6��8�b����]A�qVJ[	J
�u��v�����k���PC�-��I� ���Y�ҟ�<�@B�1����R����Ypmݥ{;�35<�7���!������-4.
���3�ܭh�[(qp�����in�@j����̙����G`�. w_�p� +�Fބ�g���2���(����I�`��A���T<�]Qc�t��X:�pK�y��bP����^$B�c�v	�����F��]n_���_��n��}��y x�N"�j�R�x"��O�_�e�=Cg��f'K������c����ܑ~\�&m-E����s����-�$)G�:(�JRq�e��J���iO��)Tի �ƛGX����w�0�,�m��Lە��).P]8��p]V�:�x�'TV]HPT�[9��m�R�2V�����P�Y�!��ԥ��(
�&O%"'O�cO�9�=�*��8cP�R�LP�<e=�-�,��D����}�(,���r����tA*�^Rm�6�x�RH��޽׼��͝H
�w�n܄y�$�>�A��m�aO��a����������.>h8oA����?_�#\��I�~��]�)	��v}ksdyee������Teu�P�(��K��Ah�}46RK7ߣ��y(d��� �&���8�`���mv�Lr6����_������]n��l<��T�q���͛���d�`d�f������tX�������[Pl:��_"o��ӳ=F)eA%�;exa^����Ű��&�1�.TX�ؠ~ݓ�#�|�قUP<)E|��b5��"6��c���;�����)�}K^�f�{t:�J�I"�]��L����Q^/�݁wF¨֓�B3Ǆw�^�YB�}u��3�'������j����f��]ξ��|ؤ�uGsWR!q���V	ҳc���ĄR���m#;�����M*�-��ǚ ���$qº�
�F��]gpn��؍C;GtR�2v�*m<��s�G!x!��,?ίk�jlI%��HNv��;\��Br!�<c�t"�
8���������,�GOn���#Peq\�`$�b�,�믿qՋ�ۋWmt����F�q"�`�2Q,�KB%�xS��MeH�]��>��ʈd�m��2߀L��	��z$�g���P��`Kȇş�i���k6�>�0U4*/^z����ԅ���$���M�Oa�#�nN�U�U��řy&���o4�\����*��YD�w�%Qua����#pP�L��[�m�O�Y�����Ѳ�h�]��Y��!���A�p����KKG����{S����B`��    IDAT�$�KGd������� iGl)|] ��c�
H	|��ss�{ڋ�/��x�D�_��_������.*�d�J!�E��. M@��¨�Ã3Jhԩ�(O�4j�ʜE�I�SF(ҁ�y$6�u��MeP]W,��u�c���;�*��T�{.�w��~�]VI�2�\�'�������c���/a�щ�HB�o��Ǚ#x?���o0Y���5&�WB�	�\���U���f�%�+�/�=w�0�6?z�Zȷ)�2xt�3�z8�Ԙ�ؖYN�k�ᵋt���i�����^U���K��X��mf a���~�ڸ�u\�4``�B,���j�-D|s薌p�[��X�/�`V�(c%2�av_ �G���=V�8�5FDzN�T�w'��?�����w�kv�{f�;�����j�y�y���p>���#���Aᧃ���X.��eTD��E��9�:�DӲ�	G*R���L�Ι�͛Lޖ�X���\� �,�;y����-���D�&�gf��F�;��Ǝ ��oG����`�� ��Ӽ�Y�?9E����l��A�䓟D���%�_e��F���7�T-�Ă"�\X ��>�}
���6�#�!a��#�B�4�s|GmۮB�0"�D'��0Ϸ	G��~��ܴ��5q�QU�h���&}�4+P�6~��)�Kl���cnӊk�SJ3�>G�B��<��1�a;\�@)^��������ɕ�g�]'��<���U�Qv���>Ԝ9��L�\���\�/�
��O���ocJ��NT�2Q%Uu=�oģ��0�.���B�sP�׹���������O��^��\찂��ajj͌N�����4~�<H�d=�s�	�g��v��T�مMR�Gge�͛��ߺ�d���4�$��J���?h��G�1��8���9��e!�Z+C�*mi����|k�//m�t+��7R$�q��?������o�.8�/e�VHv��cϑ���D�,[jB���c\���%B��d���x27�k�f��@.K��жW;�y-������i~��~�;�_�F2.����c�8>OX����_Dķ@����uU��+W���pr�@�=2!&x ��M&a�DXEaqc����[R7=���
��[�IK�7��P��]��Fѻ0wU�E�>�"�P"���Lx������7����Idf�`�k��me���{���Ds��Ǜ��1���kq�<�� )a��JJ
Ֆ ��ؔ��K9�� ۰V)��>Q��i��5�6팧mZOM9�)�	G�|��#����[b�Ka��Β;$�q��s�@��_p�B� ��{g��mT��M��{~g��qU�+����"������ٵ楗^j~�7�9w�Ls�!.��e���1nM�������;�_�P=�F�RZ�xd5,�`Аi%�H(4[n%��Mfb�t�^w�Fy���<+�"G٦������~��A�
�)��Ov��ń�Clʎ�e�*�y�8j�ۨ��F��L����N��Lrw�?���/�Q�v� R-?��&\:�.+��>~�[�fQ���&�}�_�m���o�u"�A܌8�q���ֱ<�!���:�z��݃	�fe���P��]3��&'���4�;��Z%�.�l�"6L�@+���wT���A4������L/Ø��%j�EKJ�a<"�IPT`��r�+��߇R�5���_r�I��	��h�$o�����3)c���U�&���1�EU`OHoTv$VT��fcɗ`h�c]���t6�Nq?��m�+�"����l�F�P�����@4	��&�O��&��0y82��8����VHE��/�ʪ"�JY;,
ua�6`Un����\���B�����b����pM�� ��
O��]��=<�����Pږ����f9��y��h�{~k�)^:E�I��c���	�԰@��v�:7n���d�A�H���~���&=I�����8�>����]l[�p߭�ᇉ��O�$����ߙ�n~g�	�T��!����`=���{B�f�/}�K͟�髰j��j�)U��b2'g��E�O@��X��V=��F�BƮ��j��	\?�LZ	MR�,\��Rz�AK�aQ�U�M��<5	����`���e���K����U�"<)���"���Jʍ���F�A��ڈ.
��	b7��[P�;ȹ��X��<�ؓ�����n�дܼ����F�
�Zmm��� �D���529G���}�d��G����i��G�u�oG ����D�b�fg�����d���@�d��1K�9&r� ������������.�.��̹��FE�� ���țk+淶F7�A3y4|hڠjT�4LY5���7�˿��(W�����g���t����ʟ� +�� �L�<|Q5^���_݈[��;HdV��
H���-/��Eˤa)�TG��Ƒ��|�In9������l���7b:��Ѫ�IY5���z8�U�ue�mpP���EF��\~�-p�nq
6�c�g����;��c�V�3�����_�~����(Hm4H);��'�ز¹�D��k�wS�]A�ҾuZ�ƒߓ�����]��ī �`�u�ub���JKd��=�2��p����u���\�cs�R�_k(P +׆����{��V�F���� 09�G��t�xh���e؈����q����o~���_�c�qq���A�6�5��Ų��<H�0�OOAڛ�ڍ��[�����#x|�e��j<�R��Ҁ��ičmf��`a|��C7�}�^C���
�È`���;2�k]5U�:g��|5�{}{y�O-��1a܃�n�������赟z�y��w`5�X}
9�è�.ѡO4_��>�#'P�� P��p/D����6(���G�z�"ڔ6���9e9��}W�Y����9=kosks���}�2��㗸$`�8�%P��ytss�� bS�ZꣿҔ셆kcE�����n	\��~~��"���X���{U��p����}���_�|�7���)9YXx�	ʇi|ON�>�ô
O(I��w�����a��My|���nj�Έ&6#L�%-� ��XDY��I��$��۰8�;e6�RﭱU�<�sU��]V��p��?�����)�ҟ��K �n���W�h���(�#
꽷;�|��Vs�:;�鬷����0�H-�(C�L$��a$�~;���Zu�8ܯ���>����u��w���V�?k94��\�u�Wp�a� �$��Z�aw������@�IdvWNj6�2��q����E�'��}�0x���e��;� $V�l*]�����H�����?��PM� ��qg��d�ć~��~���!R��<q�,�������н�v�[��"��ܥs���{��Ï����u2����*���65.�c0+G#���]v��`������b��#�A�)ܗ��������1���*���͇/?�&���{|@�6�������_i�M<dg��*K�^E��k ��bC�������_T�H?���@��S3��`���#{��b�)��bn���'�ߎ6�B��N��}�

�Td�dr����Ϊ�bA���N�$�fq��>��ne�����]��w;�(opЄ�8��dr't+
ߏj*���_dQ�f�}_��N����� ?��U��\���w�� ��`'�x�ѧX�9�,]{�Y�}��F��&���ȱQq���1�Un����ܜ��q8.u�S�.L6Y�f�m�5T����w���Q��gP�E�wuce��>���s�.�����h�\};��MM�h�z��t�x�u.oz����E���-$��� f�	�	F4��XŶRN���BJrGP��:�ui;B�ǲ�}K�O�-�<��p�� �%r,�fUdg��%E�� ��K��Or�Eg��lЁ_ܱ���4$�b�'����ɳ�8����������'������PA5�6]P�<�-W�e�(�տ�����w����/5�=�0���i�ns
����mx��P4z�����x�y��[L��u^e,tY������1�%^+�=�W�7�X��;l:VG%�Oa�I�=v����0����܅�,6�o�.6�Hw��B�ݵ��ņ�吜\x��'>
�\�	�[o��|��y��7U�3��H3Ok�+�!�Y��	:�@��p/~���1�*��'%��g4u���Qzc��%�(�lR\�
p?��?�^"9���J&��9r��{���(�OT�V�����h�5\�؉��/G!i\������X���=��6-����d'�A�<� g�"�mo߅M��6_��d��s��<G|��;�������g�����#X�h�����Ϟ�r�zIg���de�ns�]�O��7@�7��;�P��d�9F�	*T� ��1�i�w]�$�ͥ�97C�a�f�+9w��w�xͷ�����?D�{͕7ߎ=�&��kO>�qTw/4/��F�ЅǛW�����I��+�Ҳ�~�|=<�r}�Q��)��`K9��#_~�ؾd;�T]�#L��]ڿ�uf����4�`��fgΞ�=����.g?MЦ�|�9r?�4�>{ʔ�r���w��M-.���5d60̹��@H%X���-�9!Y!�!�����l�@
�O +M�H�d&Y2�/��oTH�Ѹ^�� Sf
+wʩuwO�;��c�������=�9X���z���Dl������c�lC�<�j��z�I����:�\8�p����W�ջh"��iF��<��{������wY�tTpb�̺�=Z�/�5��l�~�4�ف�G{ԳXPt��t0WYY���=���.����WG�kWO5������o�f����,�~�
�o(���@�. ���77?�Uý $��^�a�?$D �b�D��D�tp�hwޝ_y
�ߎl\&�d>�5�c�j�g� I $�ۨ&�)b����7����{I)M��x��V����\����&:�s{4Ю<�%���m��V&�0i ~�ʂǕ����6�t�_�q3��ɰ���>�	.rV��?��4�=�W���K��|��A�����2=�Hl�Z9�\{�G4�Xs��
�p$,�<���m؞E�X[]n�.�
x���N�+�q沼ƍ��|���7���4gΝG���h+�6�Ї�����eGJan/�B � �S�6��� �������lmQP'���f��׿l���s�E.���ĳ��pI�.�sT��m�|�8	�L?ä{Q�*�St\m��nJ���J�s'WkQ?�L�������W���.�n2ď/p@z��)SS,:LN��ϡ9%O�C���M"}��]V�B�ܥ�S�a|���3\�kk2��U~=fN�Ņ�(E����}&�������泟�����[�6���	��� B�Bvj�Cl1Xm3�{�Ή�g��<DgagM{k��?�ݥ�VA�E�G=�������-������2�b�����?K�@T��ۻ�2R������M�o�m�z���^|�N�$|g1-/�Lpq��$��� ܄}��>��/M�g{����SX�fy�V�r����������j;S�̇��Cn�m��$���ڙRc�Q�;3;��qoy�mH{���P�"J��-;���
kk�})nx�?�!0�5	�3�y�{��N3Ͻ�o����ΩT�|���_��|��h��ȇ����O7���������Os��$�>�\��@Yذ�����^J���i�Y�c�P>�L�yy�F�V��MOrM�z�4����+�4��WP-8*V�����I�H��~��0��0�$��M�����	�LL��L� M���s��?�J#,}�,�g�����v��~�6�)�Q��q�¶�2�r�5��M a",AP`�9.rCb�ҫ�ؘ�;�x�^�Ն��1�Z8{f������f�+����6�D쌛��1�_�|�P�W�JI�ƺ��L��.�a�������4���������qs�҅��?�)K���9��N�U$rh�`�ץܻw
����4y��[ל�r�H��]N�e�:��Y��v�F �H�2���N�
+��v��Ύ�A�]8h����2�:�5+�N>��]�Mt��k F
>��m�ap,��F�!�2-C�6)�QM?�p!}�e��H���i	=d�ҥG��}�QD���흲s�M{�ul�_o�_191��<���� A����̘4� >��w��l��-v������2\>�'���M㷏��^�2Uܨ��h�IIfX�t���o~�y���a�d������ͧ?����s��󋁬��PTTHY�]�\ZZC6~�d%�R_ܫ��6��}�.�Ŏ�]&M��W~�n�[��`����}c�C�ud�xY4 Pz(7T�r�	�&e>1w��X��Rt�K�K��#2	����^?��>*�:~�6�)Į�E�I�f<���x�s�ɺ��31={��D���<G�92�������U�d�����I��S)T#T@�Cӈ<��A�d�ׯ��V���'3��+�wӁ+�)�&g�y
�j:�lp2�z(�Ȯ��4����Ss��cPՉ���χ}
��S��4��	w�Oq}��a
EG�>ù��(Tv����x�����U��'Sy��w86&W�pQf�� /�Q9�.&Ċ��g��U�wx�������J���~�[ï~؄e�ǧN+"�?鞶Ά�W/ܤ���izq��Wp��yn9U��ܹ�9������b*�S���A��>��>׹�q �4���B9,��M
��OX)ˎ�
��+j��7�_׿Fd�u��w;���w��v���w)�[X�B��( -+�S�ҽ���
��ߏt_��o5��՟�H���w�g>��泟�,�"�:�3���Yi���&[����f����W��|�w�������C�/����,�c� ����Z�(<=|S�*��Dd7@��(����t� �����O�j��0�:��{�lZ�@{'��.Q9�C;稫��ťK�Z��^\.�R����{���݄���Z��|���)y�0bDj��bں�॒�gE#2?����2X�L?Ӎ��`��1�o��d���H�^P.�
�
�p���&��F�ӥ�<���[���4����������'>��,��YF;�g>�S�3�<K�x�����k_��P޵���p�ɝ8�vV#��V	,�n��K��� G(l!
�,�0RN+�Y.\�D�:֡�]� �m�$���%,¡�1��I?��w��3h1D�tK;��Vit���'�^g0]�HHYB���+W��?����DH���ٳ�2qF�ћ���Qj2G)�{�":�QunX�`"�&��w+#`45b�4��J��0;;�2���"�j��>�hZ+�#Vq�8�q^TF7�za��P���7/8d��׿��X�Yo��E���v���㗛ˏ^n�g	������
[�)P��p��R�3N�P���ɲ���s����������,�c8��E���0�+	ۂ8	'�M�׶���d��=��^{f܄��i"n�Q�)�u$��]�rz�W_�
���G�>Og~d��g�,�}��mB����ۂ!�Ʌ����d�V�D�t��w��&�j���>*|ݡ�8��v�x�m�2��|A��9��*Z�=K���臨5(��G����m�[yEny��^�Ҽ���܉�mΜ?�$U\(�����Y@vl��"g8��e4q� H�+�v݀  CX��C��nvʣL�$��c���w:�a�m�LC7��N�-�
��\�ZI��E��)쫣��L��`#'9�i�d��y�[����#h"���	#8��+�ʊ[�xĖ�|u�֩��;�?,�����LC ��}6҉L�����GbšR�bX���(��qM ��8i�	��Op���8���ltU8c�EG��Nz�	l��RA8+Tٽ�^��DHzY�0�-.u�N:��}3#��*a�߃��}�[�0iZ�������U�C�t��,|8=8��I���7y����
��Xj    IDAT�:.rC��!��C��ua�<.l	��iL�l��.*��U�^p�B�
F�~�>�³�1�^�wV?���~g�Ek%�_�'"_4�X�{���@R'��}��db���pl�"��;&��q�]5"�\��u�#L���HGpC1
X����7.�
��^��Rs����:f�e����0i[�2��%��ݫW	܃��5��6�n�+��V��K�d��θ¦�R��#�mK�A��$�i�C� &L�Z�>#����p ��r���e�_Z��q'���,�O11����դ�~'Y�L�p����a2��K�N�4�b�( :ÔR�/�&�ƙf�a����zxfHH[h/QRB"ew���8X'yIw��c��v �)cn����@L���|!x����zdӱ�=H4"𐟄U��U=KZ������8��{������m0|���OyO�����:��YC�(lXa�ĻKK��X�����m�Y߇�t=hjd�̘?tG��B�;�V�P��+gE|��چդ]��n�դ��2̠����"r�qZ^/´iG�d��3��8�Ӷ���r�w�KU���bCG�n��N��@:Oܘf�uo�.;}�b�JU���z��/U3n*[��-���p%���/���Z�R���r/a�	��Z��l}[�6!�K	�o#��E��N�p�'��K�|L[�W춠VO	�+��w������\Qs�(��.K��ذ!f��V�E�F���%Y|qX��hYP��6�7�a
P�=\��%��|�a2��g:�G����gZ�1J)�u:���"��Y��$k�.�L�,���cޠ��W����S3!
J����%��ɥLN"�
ȷg�n�u��qe�UZ�;ʄ-�ηv�#��"eY�`�i��0�m�.�|��p����o�k�:�~���)�Jx���/$JIHsq���YAv�mcc:�A�G�cSnϻu��������&�����451���'�/*�A(��ul
$0(��PƢ��2'���|�V����@�q(�Mi���+v3��K#c���zR�?��F �Di�2qb,�%,�hU����gWM�K#N���$p����6�Cs��V�o�X�|�쑮a=�d{��c��)BZi����nl�(�W�X�,��9ҳ�i�U1E�,ݵ~a�¡n��>��������x���i��j�Љ�CX;e(�a���w���1=JCMAw>M��nolq��̱��tjԳ�'Bϖc�(����F �S�@2�QS��w��mc x������N�&��wڙ�a��n������_4�bf��W�C؈~OvA�;�+n}� ��2�V�!���8Y ��WsX�[���{�����"��=�h� G~a�d	�`_vİ��3L:SS��A�4�Fn�p��THr"E�%��B`G�̂E#�ȝ2���)��d\W�2��h��
f8��d���4Z��_���S��0�vD�#~I�_;]�y�߃�&�I��q3~���Ҏ|�G�3��3�0{0̃����a��a�s;,��T��)ÉK>���th���0W��\܎�����ds�kJ�1Εsa������-��o�bJ����m��gE#L�,?ϯa���-���`�t7\R��C�7��|��|�ߴ2�v�+ǍΏ�TJ���Y��˸��a���ؑ/�uzu��t"l[��~���y���3���,u��1g9�Hʹ����Zx�)�	b
I<��(g��-�A�5
!{�U:Q����<r,R�g\y0wD{!E��b�nAM�':��}Lô�����dڵ_����+o�1�=���e`/�.�}�_;ޱy�?U��I��G����w'�>��dxG�ވז%��re�>��5�V~k[�(W�Ϡ_�^�G���c�sX��O^�z�K�ޟF=Ac���؅��xo�H��sQn(2eQ���H4���,MaDz*&X8+0ht��{��q�����}0��oÛ���y��i���)��4�3�;�]��Mr3ﶺ�/!�M��@z�Nh�ǰi���m��&���@^��鵟u�poӬ�3f�i�skz���m9ĝR��#d�8�3���IC��d����`��F#	!�\��D4�J$�(o)��}Ƨ6	�t�oä��T��]��p�M��W���ƩM�g����O|ݣ��ѱ*+~�1��">M�a�4�rK��Ԅ݂*.�N��D�M/�p�c��&�yT�{/^ێ��`�m��dX���Bm���������U�:�������R;+m
���0�?j�X!nO��������V4"�c�d�t��:��+ Ȱ.����3=,^ϿM �h�_��[R�K�q2�an��i�e���|������r�wڃ駻v�e�xo�2�`ܬg�>�n\�"L5�.��i)#��/��a��3N@z�96r���Ǣ�x�E6'��<��@�XU��DP����~�DA~;*���L ��v��F�����8�[8���.W��?)��d����[��������=E��k2-��t2l	���ю���6l��μ|7M�i����H�jS���W�k�`;���	C�3����7�u���Pf��u6b��Bܨ�Ɏ$�E�6h0�D`�3zk�Α�ɱ���Z��d�0���^��*JV
ju�����6��ig������8�l��x����ey��'��8�n�緋I�ᣛ͒i��g�h�ϴ�i�y�P�o���"�j;:�v��v�=����["n�Y��2����z�q��u|���[�6�)�	��M00Cb3+���=T'�����N�<�=v�CՏ0�Gnd�/���߂�߇/�&��Ii%!Y�ao��E�(!��[�S ���n���vX��������m�:y�,q�7��Q϶>�!�V��G�L���ȡ�O�ɲ�����g���̑��0!�m=3�LCgœ���x����#���p3n�+�Kăm���%k] �*��x3�^S�u9��t��tmm>�:��C����S�m6Sx+�����(lr�0�%�U�1o�5�"��
����u��/ݵ�=�]���j��{����RQ�u����ښt�w�3���:��w�ӽ�o�����^��'�M/��O�yf�����u�7�|�N�m�i��(�rd�FNU�6�+�=tq��6Ϟ�~�#�q)w+*��A4�%���}��w':N�qA�
ʬLZ1N>�1�,�d��n/�M8��˰=C���U$�&BԈ��ie�3�(i�� O�Lw���5��l1�n#�f�C�^�(s[�3~/,�,�w�[��T�[�"�-�3=��h�w	Q(k�kg���������8��'�i����m�k��N(/~H�U�bB7"�t��7��4���q&�Aa�}�2ԋ#M�GTlaő�n(�P�ر`�Q�'Y���jx�d�0����⦿����rS#���>���du����W��nRk����n��ս~L_�|�4w�=�r�������]{X�_��^�y̝+�Pn��gR�N���v���s�9�s����#��=���e��;r���	���+G~ æ�f ��F����XAW��I��6U�tO��	�L��}ϼ|�͠{��v��3�nX��c��kZ1�gtfq��T����!������,S�����]�A�����el#�n'K��9�N;�{X�u:�_/�/;v6��t�n.E���)��Z�a�����%�%��1)2�dit���g?Op������4CI�m�*�8��^������~[���w�����n��B�=�nz�QS���aܡm|�=m� A�D�*�q#m��zؐ�K~۠��Hl�@��{�a�,�@�(S����t˴�=��'��;ߵ{���Q�v��а<���a<H�F���*�r��ylO��mV�8�]��sw	�}Az8U��fشН>1�.Az?��8;R¤\�F.�4�
r*��JU�|VT$pE�NP�u����>����'�� �1��Nʘ��]SO�q��$�k6@�x��)���5�9=�ʼ���!���E`��{���*�:nl<���ٔ��:.ZT����������Y�D��8�e}�q��x�<��?Îia舔��w�a����$d�ݢ,�u�����7M��<��١i�� N��%:��B���i<`����'h��7�=����Fan�X_��;�#ڡ?ǥ�d4���w#�����y��1�q�ݲ�-�S����l����4����9�V�o���Ŗ�%�& 3��O�5��w�hIy3��3͌���4�6N��{q9�7��=�Ю��u��ޝؓX-�o��'�_��Ʃ�qZ��H?3���薝#����V�a<W~��_Q��(ܸ���N('�����t�N��b��"��a����{�8�{�S�F�KhA����I8��Ev��V��xÌ@�q̓��o�H�6o�R?���.K棝�Y�9���43�i&�3ݴ���~��ߠ{~C�	�G��#�,�0JS�+��EpM�����0-��s�Gj��3^�=N:�kAG;0�ā<Q6���3��;9=���w�}��S��|��V "�� �[3�!a��&������=��m�fƍ~2,M����_����c�A�_�0� �]����������In��v�{ �&IE�!ːiG���"�2��Rg���F?��=~�i�g�%^v�2�::�t�]��f�דw��ά7�d���~���+k������][�`�r�
��vc�o�9�D�sߢr-2��� �"���	��0 Lҽg�n�H�8��A^��@hKy�o�밙W��w������e����g1�F��i��|ҭ�3N��N7�x�D�˷<�O~����_���y>�������6M���m�>�hX�ͭe�/��R ���o��,��[5�繁��}"�!�a��S1�vff�7]*uq��*��V��d#sT�%bg�Q�ġ�Z�N�!,)H�|�6���'#µ�v���u��}��/�&�t��L3˞��u9�{�?��|�Idlᓰ�8i��.(oG��;M/�<ZO��oq����.���"��t=�L�!0�_|q�2j���p~��'NMNL�ܾ?;7�[�A����d��
���nT����:=8�6D��T'�O;����d����ie�f�t��A;��ݰƷ��������fx�A��6����f�,����a�.�;^��K'GH�5�uI��-¶R��iK�J��S�=˯�q4q��˗C�D7ÑO��g��g�ǀ96�^���8�iT��R�%��cۛ["����H�X�@��2�X�u�1#�f>R��v�eH�gڲZ�r7��mD�!?uX���7�,������6����t>P���ii�̇�9�\ƣ0QE��巔9��FTe5�4�OR{�VD��tK_Ǎ� :Ú�&Jӳ��#��Dt�9>~j����G"���Q�C~�d����P.U�����o�MLm�r��9o��P&�������J��#'�D�
�[ �0��[��_6����&��6�,�ț�~k���A�<ـ~��1}��|�]��X����I���OiSZ�h�?P$}Y͂x�oy2/�����y������]9|�P���e\M���<(��+�&��c�l��p�X.ӊ�X�./�5n��.��E�%�w���������햍����?Ǧ�Ԉ] D�u��!d���qoทh
P�<�(��T�TZ���U�����W��_do�p H��i�/.}�g�mxJ�Ko0��ʐ����D�U�ֽ ���".˘��K�gx�f�?ː߇��yfd;�>ᇝi�ݖU�����i�S8�c���e�8D��N۴ヷ�Ep��歟����2��>6r#��S���x;�<6��M]��Np^��)��)�`Q�f�WX����A���z���DP� ��� ��A�u<�3�t��=dh��8Y��/]�M��'h�$�@�#~]��;����01F
���t}w�2LFd�d��W��-S�7�M;�%d�]6_�S�H��x�W�Ɇ�ϥ������.:���C��3���].S,HvY��rF��P>"d�K�"J�SF��AjS*��u����T�4|䏏���`���2\�#�3d�V����2e���ƫ��ib�}|�?�@ϸ�^�#�z�F<M�1�D��3T?ƕM�چ�%��h�^
�-s8�g[��_��R�0?({>~˺��k��rmm�c�����t�9>rsF T�;�F<�w�߹z�����X������De������l�D^�&a�v�m���%l�Q�K�/K��6N	[�����)��?����K���o�W+�m�,g�d"^��6qL�������o�M�Y)��d*fݨQ
��&���@H���8-�5n�G;�Ԅ0�ގ<b]�׾ѐ��5�H���لrd�H�Ȟ,.������	q�%�I������C�IA2�k)�������ٵ����+U����0����zŲ�Q��!,�����u�`�H��P5������@���42�v�>��q3�ߙv�ND����&��IEu�"N�L�ș�l��_I��-�A֩��|hĤ��*D��vVM�e�O�b��}?Y�,?��I�L�T��J�,�0x�7�z;��u�v ��@s�֭��ӳ�o��Gzf�a6sHq3N��5�\��qj�\a�+�t3�Ҋ��T!:�3s+�4TVZ�6鮛<7�0ݾ����4�=����������l�3-��hg�}���M�s4����Y�^z�G
�C�*Z�!ad�|7X]'%#��w�*��k��r����\�(��3�n	�˗/�q��Ery�3g��fKN����Ǧ�c�{���b����o����Kw�./�z������fc��Ie���R�,�4� �Ү�{�~�[Z�}�L��f�A�H�u׿��<:�a4���s����w��-"��v���j��C�j:t\mөM~�~	K���#-`�H�q2������"��uGY?��-3�}v����g7ⷡ{~m���w��w)��0��p�a]�/��/4W��aܳi�VW���D��p���ͱ����nq�����?���~��G��_���%�,�xyǁ<����*^��a�he� &�cx�]_��%���W������ ��,Wc���P�D� : rn���I';D[ j\��Y3aB�,�s�D���R��f�.A��e4>�"D�eE��R,�\&��x��	�mo�f�dC�g���ˍg�����	�b*�
�4�4GX`��A �N<H������W�� ��n'�p>y����(�G^�W
#T"s�>�O�@h������RG�R7�i�4��~�R�4^|p�扽��щ���0u!�w��X����]5����޽{���8��}�'yD+���������;��O`�i�/`5�x+���H�:G�Ѱ�N��+�Ӯ��M�	�wʑ�Y�ϲi;�v�n��Y�}�ʶ�?G6�2\)���l��)<{�>4v�o<�a�?�,_�~�a���a����=3L�~�V�~���0�G�gx�&KKKA�� ۸�4���M����#��ʠ\���3���\������A�&Y�^��ʻ����~�f�0+0�,,�!X�`�
��bC
i� $�Z���/��Eb�3�XzLO�L���-�rz��ߩzo���� �}����y�ɓ'O��Pu34x �L"TXQk�߻���5͎���#��ߒwL�$H�`�.�x�E����o���ʉ_���`9vފ��۬�DL4��X\�]&j���D�d�>��s�%����v���
8i�#��6u�q�Ӽ��p���ģb��Nެs�_p������|l�;n�e	K����i:����+�m�󷣻0�	�፧�k������T�{��M�� aS��c���}C���m�[�me�9P ���ޫA�u(�� H�)��'Ț Ͱ̿�m��qC|�9�n������ST*� �'�:�yQC*W���{`���89	��	��!�\ۜeґĖ�Ɏ�&���AÅi:�$R���    IDATz2�vQ/kk�P�(~\:��߆��EF�"��n�7�#n�O�7<g��oې��?�1L=wҏ��<�Qka�ߦ���7q�l/��>�&7+��ܡ���S�o�C�
�>*t+p*�%\��@Pb�w��!��iZ 9@ƿW�Z����P���x	e{�Y_�,�'��[F3���~�%�Pm�{��y9W�v.9�:)p�D9U����(�6!l�Q9�Sۦ�G�-�Z�KyN���j�j�B$EK��N�����Z]�1�i `���m�E>�Ƚu�%Hb�q�V�k���i�!�5�_8�����e�[{��o���0�ۦ�U�
�3�7J�M��76̌:n�����FG�6�  �#�f���qr�'; ɢlP4>=x�˯?�͸��K?�I���f���2,�R�5�tƱlo+ST�N6k��v�q�[˴_W�hsnwNE6]�Q��Xyӄ�Q��<�P��5�Z.0�3.��SG�����00�I�n�lk�}/�j�*�eX3��2M�3N3�f�2���WK;Ju�R�m�E�����qk,�s[s��V;�~�(Cx����Jg#�a�9u�����lp��Ώ�>R������Ęqrk	�щ����!u<�y�1�O��wn��Pc*��w�+����Ǫ�@�Ͻ��e�Cekr@��`��D��Y���e�9�%��!acT&�d�z3g�trx5V��~�3^�H���g�n<ȸ|�T���n>�4�t�6�ȷ7FJ~���c��Lo�$l;�D�O�6���v�p�%w���/����n�_�At�K W�����M�I��?ٰ��6<1��4��;�3�j�(_��n��������-����׶3��29Zpb��1�5�#՟���N�=Y�?i1.��].G*+����!���O<W_E�����r�b-�J@I�v���8I�����('�ǯ����r��\l'��Єg���g�a�m��M8�d�(�8�.����~�4��Ҁ���靃({[�b�߈pX�m�o����Y�ܖ�����?�t�؉ٹ�Yv1T1E�XyS��_]V�J�x	�l�a�峍���3N�D�@�pަI@gj�!�s6��oE���t�k���b>!�P��E�qɸ�7*�������~���/y�;ʙS'�[�r��yzv�����Y��@T�O����g~�_��7��a���M�P�,��n�G���h��o��!���O��0�j��/jh�;@���y�j�5o��EZe)]ԧ��߰�'���y���QRF�O�L���V��h]��-#ܶ�0?yة��[��[F��z�_&Q�}hKX��s�f�gʥK��&g&O��j �ȡ1>: �uM��8�g<��7�n�����_$|!NB�� T�@�1qR�0��.D8p�]������#,�,/�I6ʻ�����|gy�����F�=���A\�f�7р�H���n��ɢ�n��Un����������/�ŏ��ÃC���7ʇ>h�)�W�];Kg����m��Ω(C쀭�&<~���o�����4��m�$Ќ��ɷ����;4�q�i-#�}�Kt��Uƈ��Y��ǟ}7[aڬRm-R� 㤳����O�M���È�@�{��g����������S�P�Վ!�3>P�a�	����9���4���c�@ME���㮬,w&4-n�],�������a�������3g�F��;������t���Ъ%AL�Z/�+Kс�ۨ�P��n�@�̗>U�㻾���o����� � ���#߸G�vKW����au��m!Ǉ�����f��ſ�ᨶ������e�q�m$����5��6]0�x�N\>F�L:��q�dX�M�d��D,A�F���x�@_�@{re�3�xß}7�!��t�{p�Ņ��Y�=������К�͜��I'	 l��?�N���̣Ǹ��N��n4�yBt0�^�hSG�8-v�&�,©����ʷ������?/���x��ܭr��edt���=�텐�Gǆ�2HPk�ۏN{��^��^,m�#��gv~�0�5������|�,΁L��H9�O�˶�	�KOo�t���:�Ǫq���F�He%����� ���[M�"�R�O��~�8M��	� P��6��f�13��X��ۺ��������3o�c>�x�˚Ag㼑`�웸U2o��ͱ����S���.]�|�����@T�Q����h�g:��8��ЩJ@����j琯�6���R.5L��w�ÕZ�u�G?2v�d�!qjz�<:V~�����)O<�tp��7����H�mM�P�����Kޜ���\j)�ss�29�k
��7�5���|��`5�P)s� X���A��o� � ެC���.�;�sQ�
\��=���6���X�
�J�D�m����a�*�/�z���:�6c���-F��9�tF^)R���0��d;���\Gn�D�ށ�m�d�Y��o�6'
��,�щ���-��s�6�����Z'^YjT������26"]�gC�?߻�6�3����8	@�ã#\?����g�BY�+r�U�?�ߖ�]�QN�8VZ�}{�vi��0�0�K�V�a�ٰ�_(�䱶��|�P������ksL {�3��.R��/����\Y�X(0� |����2�\F��n�3���G)s+(f�DR.�dm�KN�K��n£����L�y���4��n�_~�G>7t��诬��E�)�����D�:<dO�o�V�`�����'�li�966�+[V ��a$��?6��0g����{�7��"O=q�n~��Ov�9�=9�0����|��{��<������-�mO<^nܺNf=eim��,VʁC�M$ N�,K�a�Ņ��K�(tn�[Y[(K���Y����UeN:bIԍ��2�����C�-��(�T�C�O=���V,��j�=5����U�Xu�f�颭�X%��7�%����;Z������:���¹�o]���|�=�UV�6���89�J�T���F����W��{n~�d�}:�p�9�z��Iy��-f�}KK�C�����:�A�Z�d6���iX9�9��Xc�L�O���ٔ��{�,O��K��dp�<8Q��뾮��/�<��G���g�0�v��,hJL;=WO�w��6���ѰeĔ����؊&+�p}k�q�hKBd�x^ڵ��qtx�\�~���^,��?�n�zQA�]�ss�,a
{���r���N�=S�H�� "Oߌm�vO�)`[�.`%<������?k"$�vǈ|:�)v4�J�%��iį.�,�wı}�/�ŏ�0vt��2=3]&����9��훸�v���n�i��GZ;42�422�b���BD %"�UW�X��y�٨�/|�;�6y�="�'�bz�6��.��:9�����ȷ�3�;�-���o��������������-?�3��,b�8��X� ��eF��!؇ö�K�=�\�|�}�K+�c7������Pk�](]}��@��� K�uu��i�Q�G0{EDi�_�n[e�`wz��8p�<��g�����K��G?�2wg	9��ϔ2��0~`��۩6�Y��.m��+�.,Y�#����n��� M�&bL����o�ո��$�:�1L���HO��h|7�PW9���O�f4#��#A�L�[�-�����RYX\ w�V���ӲN.O���M����H�nB4��f�jn߹Ӻ35}�ƍ��rC+r/�� ���fx�U ��o��Wxm�������p�$�*/ S_*�O"�_���]�*_�~��'�SSwB[6�X�4 �A\���OȡoܜD.$��M:�~�et��������#�aq�E�ۓUMj��6S�5F��h��p9��q./��[�7^���O�x����R����-�{���0�.�=r��KmW���.᫖�F��$NF��2��h3����w�%<+�Ubn��;␮7sI��̞B��S|����5?q�S���1D�eĿ���-\e`��훸=f���2����JЃ�]#�肆�v��o�Gm�@�����{��ߘV����,�I�����|L��&��u��ˋ��������Q~���Us3�����7�!�jiK$r
��B�=��$���opS�2��YB�1��-#��b��Vy�«�7��[7��;�b�I����cTa�����9D�6��V1f�A�(;�F��0������ղ�:�:�U��-�*O<�X�uy�������k�X�Dg6V��c����d����
c���C��ֶ�D�7�Bh�1���vʻD�N���1$�T,��U;��Tg��ša�j673#�p\X�Z��T��"���M�� �1�a��X�`p�P>0q`��x"=�F�ƭ��׎s�`<�Kx�W6�����ɶl��^�t���2���P)���G�G�?�����_�;0Y�2�0
�WK����y�g��z�.�0s��M��S�����r����g�`���j��A�GN+g>����zp�"2�P\��*Q�W��[�f�p���z���/�wXb"�B]��Ï���vy�3/R�Fy�˞(�=|��?���eq���m�
m�� #��=ȩNb-��C��X!:쿙K���?q��t�߻�3V3O񞋌���nA�Ue�$甌Eݧ����R|:�;{߉�eD��ܛ�n�T��׹.Qi+nQ�S�d��eG��"�w�P�m`d��x�c��)�����5�~�cE�w/�2� �����d��gx������?�? f�@��Qg�͋9�u4#/��b9u��;dr�&����1uy�u�Y+g�?!v����˅K��(�O.�xf3Z��c�)�G�����2�`z��5��AȜ�;`��i'<|�H9x� ��iĊR.�|s�Vy���Pa.�˯�/�#c����������}���⫗�X�̈́a���KBU&L��qx�/ A�w=����t�:V#�s�?�m>Y�6����iS���$�N��By��-DV�;W������ު�웸X�:�����/�e����X�7�l�oh��B�S�t�5N ���ݶ�̼���G�SV�!�"�f��o��o.?�/�r���a]q������/?V�#O<B��GE�9oay5�mD��r�ܩ�>��Ǣ�}h�z��2<1T�f�ʵ;�����L�0�Va� ��"dx8uϘ�౔�v3�숽ě`Yd����-�
��a���4��b���+/����+o��'ʍk7�s/|�|�S_�X�E���/�Ͻ�j�7��
QJbvBg/'ﺀ+p��Y���[�k��F'yg~7��<��bĕF����S�ڕ�exd ����o�N��܍�����}7�ބ��J9�;̳S���.��u'��w���-� 8��O�]�3��qI.���څ�P*`�_#8�.�a��y��5�������-?�S�c9}�L�]���/UKw�߄p�˷~�{���$\e	�y�ܞ�Ew�����O
���W�^-c��T-��*C��f�E!���xU�ܕ	%�a��D�b�Z�Ů������ˍ��W4��3���s��XC�^@C32�.~1g�0��r������k����˷�?*���(]��_��/ï�p��MD�U�(�rw7��*�T;\Z�U"6<ݽ1��ɰL~d��M��ծ��l嶱
�@Z#�7��p^�=�&j����o���m�u�:+g,��ғ&�*ہD\i�
�X�%�jl���w�w Jw2i��8��W>�������1;����So��������Ν�ஊ+��.O��_+�,��6cf��<R�_z�|�._��_ZN�=�n�r��Zƒ����X?�ݴ`gҶ$:�256*m���+�s[S����W/�R�#b<x�zpN�A�d	�����X�^�a�}��Ce��hy��G��+����}ٺ]y������WED]߂q�F���>������X��I�:j�n9z^	cGфa��w �?�I|���m��;�o<�����̟��(�7�k��˪��ʚUP���/��6��Z��)�"	����l��y��WƬ�ĩX���� ��-�͆[�Z������[c^�E~��t�ޙ�]�?�H�ٟ�9v�� b`>	\e�ThZ��uџB�mT|�Ja�ň�z�tY�/>�e
N��?��+�g�8P��h([� �8�4;U�f�Y�\@��}>;��b�s۶�v4�:t�@���̡j��Q�Ⅸ3\����1�tN��[��}��K��.^//��jy��g�[������gXI=T>��O2�`'s{��y{��-����t�G�#�쌎����a�)q��I?���[���u�|�g���M�>DA��<MWEv+������������=�~��{A�p���k�*6+�j��k���+�	���֤k� ��d�K���۷��%L B_.g��aLy�o9��YA��s?����w��!m>�˹�t�o#W�e=�E.���_(G���G�-��w��/}�Xyۃ��o��8�(I�a���e}���$
6F�~�w�GЉ�$ƦD�nԌ�c�Ľg��5�Zc.��?:!b�,FC���e|x<��r���#��&-/~����|�|�}e9���2s{�P�o��o*�G���~��R���PAv��w��a]q �	7��O���N�8#��:�}$d]�[G����b�:0`+Yı�۷�o΀���.B��7D�KU��d	�sL����B^db��r/�  ��p3��s�L�| f.����I`{ԣ����1쒧r�:6���� �����/��������{�ɐ[����L;��=qd���xp���-�k�A�}��b5t����d�B��;��q#G�չ����$�z
���t��Q�z�\���jR�Ս���[pDH$d��6an_��m���i������c|��Վ,-!����Ĵuji�ej�/�_R.�r���G?X�|����S��O~�S�U��Uϔ?��?�6C-�փz�Is���Ĩ�p��ĭ_f�?Zx�G[�h2N�#�#.�Y@��������[�$۲�TN"�A�>6::�r�F��Hq�?�&n6�`������O�b����L(?��c�r�>I�����!>�����@�u���L�o�3�^���Պ���0;�����?F�mv{��L,���E�$�~G��ߚ���x觗]���?�ɏ K��'Y49|�@�'��׮�ZΣ��B����h:�Zȥ=|G⎉2V���D�	�
��Tn�Q�:���T�F�t�W�C3`۴� �5��W!�j\�8x�H�9}��_%���G�'���v�|�g��o�j��+���[~�W~����kl��d`n��U�J�6��u�Z�^��vV����7���o��_~'�7��;�x��0�W�b��b�żzt��	�n��=҉�S[ �" +�۳�aL�P=���q	 �l���#˩u�'����_�k~�|���N����k�c�OS���,����Q����I�\�}��[AE�_dw���#e�=SfYJ�ӟ.g:G--f��3�0�2�tKM��0�V�vG�L�Xu�@�j�f�PB���E�=t2H��U]7D��5aD�m;�E]{����z���՛�ባ�ߔu}��By�'�j��+�˥[��S_�ty��"�L�Ǟz�L�b|����u]�đP�x:�Z�V���Q>J���:F<�4q�'d�w5N�%��ȗ��v$�q���/��'9�D���k�9������[\��o�^n�7U�"�޺y+��yn/^���>1b�3r�g������o��t���w'��oôs���lC��
_pRc���7?���=��&v�L`x�b������7��FO3+!_�6#����it���aӱ�A�,�}s�:K����Ct$�g�<
D�K���d$aS��"R�7ce>�!\�Y���4��h��1;��h�cP�ҋ͈�wX=�0���{ј�o���g�8Sg��	?�Fe�<�����#�ș���W^/��,�=��5�[�X�D���?��r��l��	�čL��u�W	N&�V\    IDAT�5�6�Q�.��m�fX����;eV%@�;g���˗#^�/ 3Eq��p�pwS�w������\�p��%+t�����/z{칷�I�6R���x�w?�0�����_~����0���-@��D��?�c��qrj2��89GP�V�я�fQ�E!h���?�C�Ҟr��1�Z(w�$��r��A�#,��D|9x�P醐{GF�h^*�;FG&�ɓg!^�*�:#�;���\�[�a�{��G/�^������},"m"֬l����$WRG �^��[,r��&Y�Y�.e��>��'��s.�u��W_cԂ����uy拟.GQ}R�O�Px�q�.��q�c�B?���;:�,��W��N���V9z�(�EN^��/qc�?�C'�7����7F���g?�kiq4ڞN���\���#nd��A�lN�+�;���4i�|"��������-Ӹ+��~��2t���V`q��I���Q��}��˷Xf�x����g�!��X��d�\�q�̈�bM���G@\l&�hx)�S���hvy�6jŀ���E	C��K�۶�"$�.Dq��X�uH�� ��01�\ԛ$��!������X�y�v�ڭ�V�5aPn1�@?~��!�$��#���Yn_��_U._�T.�!���&���o��7�g<ã=��t�#]�J|�<	%NƋ| F���T�:E�d����B,��ٴ��+3��YT���g����Z�*���u�!�Ǭv����r��;7[�[	eE	@B�Qx���r����$�rFc����� �+������ �mZj:�?��B��;W�����2���Y��W�m�%�vn"�ݙ�]&O`�U�7��?W��6�c_�X��Q���e��]6lI�c�^�w!E�E?n�\i��6:f�����Uİ�C�?N�<"^L")�{�:��l���8�~���:�?�mN��S���#�SNkh�^���EwD��0�]���<�m����O�-�?�jy��Ǣ/������>\.��>�N���d5���p�zhgM1�&����#���c�S�m��4pD���G�w>�|�I��㝂6�p�g�OcW�[}23���c/��!n�cо��/qo��3����N�!P*��v�>���h����x=4��S��߫nٻk�#�W��۞/ �ܷ��&�9����uo�6պ�)�����(7��pX΍����h�����by��M6,�DgfC��u�x8)5�6D�2�\f�c/m�u�����R��3�l	T� �b�Z�,��a�����26Z;>\
z��ʜ���H�7�!g֕M:���vC5g�l��WY���|ײ�0���s�4���S�~�Xz��'Y�����0;�PR��a4H�1� (���	{�xI�gr^�����q���㛯����3/�\��"©�y���,���X�][�A)jX�#G��[�o�k �����t���[�l��l`>��o�R���@nz����\y��u:���'d}��锹gf���6�Ͻ�\y�[L�yЉO�Yw�?y�:z�u����6�]H!Zx���7���Sw�%�E�ι<h%P�u#���mq��ۦ�׽�N�5�b�[[�艇, S��c)XB���g�0sa�sw���*���F���~�3&���7nÙQM>����/>W�����(���-o������ ���%�L���n�$>�đ��N���t7��wtWI��Y��������%p�7��f���/���]0D�n !8e!r\��>�����Y���A��葮H���a>�݁c��{w���4WN$�y��?��1�΂��� �E������ٍ��r��q|�\�v�vk5�-ƙΔnV��[;<kw-׆W��axU�F$�Sk�d��VUY��w��]C�-��~�#~��
c�oa3�}�ڑW�A�����!Z�9^ �l���̅!��FY]� 
},���"������?t��ȞNl�~�����ʱ#tX����a�_x�,#�n9v��:7J�'��x��,wkP2�n<ݝί꤁��q;]0�z3�LI7�0��`�V3i5�[r�}7̢zƞeo��67��>����Y�$���H��Vmf%���[@e�0��7"��c�ݡ��}�� l{���c�c�6G�D�Z�M�sp����E������W��Ȳ9m���n�m�8�V����О���
OèM�z�,t��J����Cs��݇ȱj$MV��w�j�$�i<�P�B;W���.�ۑ���@n���!p�U/��]QN��v!�r|c��W;����=p���U^�z�<p�2�>�.gΝ)/>�
p���.q�L�^��w��q�2xԏt�eG�%n�u(P��x��X
�v�&̛���8��� ��V����`�CSiD�&r��lx����-�i�f�ɰ�6���ÕFw��)�W�D]l����! 츽K��6.��v'�g�2l_G�
\}���D�]I7�,�s!(6 �Hp����.Z}��Y^nn�`�ǈ�[M���S��'�Jؚ�
�8�U��Yͅ�d��=�
�|�����ܱ1��~h;89�Ot���тY!*�W(YWG�뷯���0�������?�YT�'����?�hy���uz�2���`OHGb�9;p��(D�S���H�������0]�c�3m��N<��ϑ݉��u�rY|ۦ�f�o�:`x�Xo��"�8�G.)wH�0�h��٘l���>�	Wߦ_5ߑJ�G��f_���|��} T 	�:�\Ἶe8�;cf�/_�T>�z=��<�!��!��%���&���e&|څT��#R�c0"'��p�t�y�ܶ�Q��<�xp�?^F��YJg`�G�uT��>�B�tT5-��:�|�!��i�o~#�@ �w�ࢢ��v\.��C���6w��E�+}���qt����:o�j�l�]��h{��� #�b�6d&��th�r��"d��|�&���?���0��3�;o�+�G:��,l�.�<�;a�{�Ľ5>�օ9�G�HU�>{�lp	�J�VT��I���ݰ�w�4��yd���%}�;�*N\u3�gjP�����nZ�V7%�m��+7/ý��Q-(�o1�rgMplf��A���JH���q�25�A�ѷ�q^q!�4���=,ǐy��4��6Z�iF�ؒ_���"C��^B4�*�ؽ�́?����+������?�8���7&�pl��HΈC��I�ѻ1�y�P/։�L��f&cdz�	�G­xPmWc����8�@Bd
w;�m��4�M�\G��1މ?�~���<���w�'��`N7n�(ׯ_�<�0m����֤M�Nw3��~��Ĳ�:���6�G��_�5_"����a�����l@�ec}g\�(��g޾M�oӛ��l�yNc�t�/���"�+;4�EC��>ȉ��h\	�=ѻ"�%�"�ݦ��/bҪ�����D
�3�4xB}�\m27:R���A�X>zQ�ͳ���(ps�N������,�ϗe&zn4�]��7�Nx�\���\#��ɽa�n�v��x��v�∓N���qք+pp��8�l(�n��,@qM�.'��{��r,�,���@9�~MՈ�OpjzM2(�(�+L+!JĆ��čp3N�ķaMB׿�.���r|�0+N�\��o�kq�'��Mܾ�{dd����JX�C� pO���$D`���� �1�$N���o�y���Y9L�f�D�q�?:ĮA�'E�(nܐ���{Y�^�xV�!�qs�c)g�CE�ї�3�`O����zƙ��c��Ǆ2���ȔWm���pkb|{k�D��Ԋ�n\��o�;�e���[lfq�>��V*>m�
���/W��W���s�F���U���n�	�~��aeՑ�c.^�j?��N�+����g���2�<�����A
�g�w�@q3�/����@ša�G��4]������m{9q,�:u�T���{i�c��j���9����z�������+fu�*���0%��}��Qy�6�FAST�Y}�f+�8�q�O��?�w �]�r�U4��4��TF�)�&�r� L�9�A���������tp��FP+�R���P��^ۼ�������7V�'����y��B�j)���W��[#�qW���.a�@Ⱥn��J����AڸH��Ȋ�ת0t��o'���K��l��r/b�O����w�	��)�8���q���\�!�	&�m���<&�k�Kݿ#��*�����r��U��N<�����������y�o'�jJ\\�a�8����\�|o��K��?��	A���}c}��	E�V\�'����9[Q������&�鯘��cK����	�R���y��7~�7F\'fZ�b[��Y74x����Јx �;h���%u-����ۊ�W�U���2��gr�(rl�x |yq�+hK}�n���y�bF���ys.�*"��q���M�Uֹ;`$����?�g�8uJ�S�{#sR^���4|��4u�j�7��G���+�ۮ��Ƹ��fp�I��y�|���娊���8��5 a�?2���1G��y���y+׌�� P[���3N�Ź����:�S:��p6:�/��s{�#��A[��pP�w�F�ج�o��ț=׼m���trg��v��3�~�y�~?��?�&�r��T��c\ۆ�8D��]PT�c%���fPNh'��Ғ�1�+Vݳ8��"����������*>*�ɟ�I$P�Ze"��i�'��lr�D�N�ـ�	)k=�YU�M�u��Q�l�v�Q��<�r����HG�u���$J�u܍�h��q�͵'Y��V�v�q�Ѓln���	�g��=|XUj�E�N�n0��¾�$��'��ﬣ�L��淿���xQ�I��n��s���n��#�� en�ەH� �;w.& %V(�+���ƷWJ|>��Cg��w>~擝i����8Z�2�zw�(Y��Z�T�\5'KL��#�0��H�dzp��,�q&6��P!����I�N��&MZ���Z�8�n�Jc����R��M�/v��:r�\���p^�#��i��m_�Q�\]QMXȤ�A�U|����Ś��C9w2ML7�f�G�!����q��.�{�n�x����ʴ�ru�M\�N(�����,]�:����?��<�-�ģ8�F�W'N�W�YY9�'q�W,	��{�u~�=NK��iNG:�p��Hl���P��F�[i+o>w�7��Q:�����mfNN�F�4z�ɤN@̡�0m�Jױـ�(�NH�[���RX�!bH\N���ejy�^L���L�B�*���N��@�=e!;�!K����|X���à�3��Lԝ3�T����-�I$�@��� `^�e������ꤒX�W��"�"�(/�����­w���z����3�Y)�=[����Z7�x�z�>|s�Q�Y��Gv�0��xO:˭e���������^��ү���_����_|8��c�$Y������so(s�����X	���y��`1�&qZ)�~f�[ �[?�C��o��(��<-[?˲�ۡ���1���l�8"ӎb����V.7�"�i�N�\Sa�d��O�S�b���y�rtȝrn�M��z�5S���ud@�ww�
O�S����@�:����/��w����\����E����aX�9��QW���>N��n�]�2X�{�$H�`'1^��cY�7n�e=�m]~�n�l��q�[�ąODʼ���z��g+�k&n��/qCT��=��+ �E58�N-q���:Z��z��)4�I�@[a'8"N�	|+l��=T=��~"���G�F�-|���f��,�Y���*�}7Co7'��[f�N�����nsvv�{�	ey�O�b	_]�`����u����6���#����G�*��?Z�Cp4�L�>��P[ro��͞�����"g�wqb�&�1�g�B���M����e�	���o%2`����A�5���vb�(&���ݎ*t:�2���ު��B�k'S����g�b s���w�GM�@}5,S���/�c�+�k�aֺ*G�]�`�1�-�"N`!>��Aa�u���l�����8�m<�|�ʫy��+3�m1��p7Y�P��5_�n�a����;	�k�8o��K�QqKN�!�H �>}:z��)FH���f/mt�SbO��~�%�$~�q��ϕ�U�\�>`y�V��.����\N�,�R+����'��7���se�x./ /[?�thR�Gʦ�%�;_�v�{�E�И�?���x�?]��A��뗣���Qb�D��f��z�͵�Ç9��)R�i<�1��-WƔ��e�����eX�ɷaͧɸ�o�.���ā�^���辐KV�K�Q�GU]�d=��H@Y�l�a�����<����	��ph���&׶�Vݰ�D��䁚�# D���3��.o+�:s21g8^�Su�+��������G_<ZEқ�h�y��n��.��Ṳk�!` 'KgX����3~�;��rP&��(y���]�(�y��+�^deG��N_�92���d��K<>�ϝO�~xêz����m&m�E�p~q-���0d����y+������}���E&�[]�2�D�+��R�\����S.gX:�� ʷ��	x�D�.���;���VW��"�H�ޭ~���,u�M����g9n8Xw�(a�Ѣ� @��{<�b�5��b�&�t�\�6L"�5�zA�Q�=�ؖlF?>���m+~A�ؙ&�u��l~7��mÞ�	3��y��n�D�@hgU1��&�Z��<��O�۰��o��x��w��v�^g�O�Ȉ�J��7o��u�4����CA�
��occ�k����܃�m�Z�X"a:���V<���o�.�ˆF��aX	T�'�;[WÀ��f��#�s�w/gs��42G5$�&r3`�p�|2�A�ڊ���"W,��rc�F�v�R���S����R� 	�oN;.�HL�сb'�F������>FM�*ڪ8$��D�-;Dc�S�c����D�;��>�%l�.�!vۤ��Q,�yZT��L���8��w*,�m?�Lox���������E5�?�$�[gq���S����^�
�{�|~X��KX)�Z�"B6��It6�	lM���8	�f��'�1<�c:;�gS�>�9�:�f��$�-��b7��� nI���)��H#�-�eN�0$A�Fs�N�S�\��9�\�O⋣�E '���{o�[�!Ĝ�R�����v]��w�0k��l�)���W���D��^�M���Y�FW	��2�ϲ�S��Y�5�߸鯟�ű�r�����/�\��IA����&xwo(�I�wP����o�c���D�E+?�L];�l��|��~� ��H��wܐE<�~�o��GU|:;�y&p��m�vܞ]�VŹ�����B�ƸA���w��B�#�ߛgٚ3˥+���{vӭ��h趰�Hul�u�o�=���(�<L�B����M'R�o2śq�pk���ٮ�.��M�c Nʹ�U�~w)����M��w:��N���?��۸Q�J�y��0���6���#������K��~K�)��s)\��^Ugeu�;��^����|���  �K`�n"�o��!V��5���tTB���f�26;;���7�-��$j��˵���Ԍ���._|���q+Xj_�6����кHt��؎h/�t�M ���	kM��#��6]�G���t�j&.5ϝ��"y).9Q�d+��S2��Q&d�M|BcB�_�3jM�IPg�a}��䍸Q�[�i���v` ��;
�ߑy*UF�u#ORo�Zܥ�W�>v��'Y1��yf4s��������/�8޹�H}�9��<�z��>����:�[��I����� ������Z1���ɫe��+�`♧H�\ì������[�٥�ȗ�9ْ�E���V]=��fh`\���V��i�>Q9�@��m���T���$���    IDAT�"����ݕ/�ԲjyvFj�����3�n���t�[�D����%6?ce��Cq��*A�&βl�0�O�ee}2ܸ:�3ν�#R��L�x:w�\�H[�np�ihMjo�{��7q�����0�b���$UoVІ����a�K�>��۴�o����P߆�N�o��S� B@��<{��=��{��oZ{���q%�2�r��3�l'����u�'W��X'�Y7�u��t��p�-�'��L�w��v�$�����2?���B�pÎ�p�5	.�aF�2��pgQG1��^�|�/�U�f�(3PP��QF�%�������W�%2�2'���O��������7q�8�ծUO"M�{��)sأG��s[)+�pW�[D�X	�C �gw��&Adߵ�TM�6-ADi��v/�-�܍���v��S��)$��DU�79��H�WC��Nc�j�U$��q�G���(/�MK��H�[��55���!
UTO�Dr���h��1�w��ζC�~7;����8v{r�ۣ�U� �э���1ɚQ�_�"t�*a6�%Y�,�r����V}��$ئ_��|�Gɜ��ܪ��ѷ�M�u4���o�^\��(�C�	���/�D-a+s'w � �o�M��?	�8����Ir����␳j��n�r��+���k�D�ܵ���G��C:9v��1ALJ�Sw���QY�C����ݠ��YO�p0~�)��=�&�7;�u�~�����L+����s3�� ��vb�D��&N;��\��E4���
�if�Ik���wʾ�\kgX�1��w>����mJ����V�Z�Y)v:*G~&?��{��ƀ�~������_�P�������d�<��y��	�b�E�Kb�m�D��x��ƿ���U>�W��p��� !"_���6/Ü���e�,W���Q}�#�>��f��s���zsø��DE���E)�H���@fT����xUd�|L˓�Z��W-G¢^�����|��+ض�d|�ʡ�ġs��\���� A{є����p���&%�!�#����E�Ο,7:����i���1�D�w:q��̷�X��K'M�kGcӰf�>�~��C6���kH�v�H`��ʲw9|˥tV2��W����4�_��6,���@棿�+7��~����y���>=����U�7/���?��D�dS���qm��[��p	X�K:��+�'�y8��m��g;��v���!�ng;v��1���,+�Q�R�ɽ%p�77�E���r��Wr��?���f����[<6?tڴ��Y^�C������u��~7��ͷ\[KԊ��,�!��h%�f���=���S��(�W�M��%2�<��F�Vfˊ4ߙ�~"/��_��~"!�d�v���Mf�٣}�]5�ҙ^"�N$��[���o��+�FԈ�h��m�ۘp�屢���+��}&�RUM�,����������`h�rl-?�_������s�K��~��X/��-A�]�-�[��ϕW���Nr���Op ��\[!W7�OmCe���#-��?�����j���n�f���uζK�rleo��S�sc�Z5{�]�Y���*��j�d�Y��w�V8e��n�nW1��(���)����Ĭ��-W��4^e�#�V�{�ز�鎥�NW�u�[�,����=q6�)zYO�ȩ^	pv�3OãL���.�f�Y��w�hr�L��������,/�3o9��6���ܹs���[1J-1�t2��1^���M���N�e5����n�5ͽ�-O�[)�]m>�0�Z�Ú���;T���g7�b���.���_*/��*�a�,CC�/w4^;\�T��𽡂�6$A[7+-&�"�2�� �����K����v���3n�nۃg>��gم�7�8����K��#`Clkh����.�Or��&�؟�;�!$8��;�1����r~��s�l�8u9������K88��
�-�ԌE$�F���s�\<`��U\,aBL�`My���E���b8�\��hÃF�7u��c���\�D'N��� �}�U��]�p�a�v�-���(ko9F�=��R9�om����x�!���X�c�1x6v�{r����N{7)o 3��^�������1�|�g�~�ֺ��{	�I�,'�^s;g�p�U�7׻p�}[	Z&�5О��T���r��8x�����aE�N��X�r�2�k������I����	�㷆:�����L˰<{�K/��<1�ɵU	Z4�����M����	RYo��\[�S��H��>�qƣܻ\v�fź�f�ߺ���ٮm����B��m]2��|"���6��e[|r4���G�˷��0�-G����ə։�pS���6��䕗^�ޗaL�N�~ۮp��|u��0}�c[��ߝ��_�8z淿~���Xݶ���r�6�=�3ܓ~����B���D���_��awۼS�(&d'�2�B��ߍh�m\�v��#�Ry�2_����/��/���8	`��=�Wm��3��2p{;�� �E��;ʈ땜��z��w
�a�躇�X���?7{�k�	gi=K}lK����lN��u֥�}g�JX�q���|��R��[<���N$,�>5�e:1t/h=�MR���Q�y[⒬��/E��<�����N�td�"�c�C�GM��v�K��߸�O2ڍk������%n�P��`*�-�{O훸ٟ�α
}K�vEP��u�vk6Ԋ&��2�͸�N.p�F'�/�Ti��s�e���O~�\�u3��L<�X�������d�"����I�|:!���p�SRo,�t���{���#�7=j���){Kt�:�V��N���#��X��K�Pm�Y�z���]�6��0|n��_Hnz��x5����M=����]:�_l��N�W^y�56>#��+w�"��;eG��~3��t@�eܨC4h'e3<}Mo3,���0m�Th�=����2��.8�n�Ľ���Ĩ}59�e8t�w�}q��L���������x	�Ls�w�y�9��〕C̡��|����=� [�Z�fc������AҰ�`�T�D���x+'ֻ3Q/����0��T���\#�?�+���X4o �>����|���}���5�a�>�\�ݖ�a�����������h��Mp�J���q<���B>|�6�w��8�[�<C��#��y��� G��Wn�Gy�|���C*�@���H�ȗ.��B��'YՇ�&������%!�q�/��;��R�b�����A�*-EوB4���7q�goO���S9۞%�;	���o%0 Aq�)����Fuz��q�&���;�gy�^�I˕s��O�4G���H���V�>��߁����|Cq�R"ϕ� (&O��}{z��E08b�]�)�.��o�^�8*�KW���[ԩH��8	�k�$s��^,$�����x98t�Ӟ����f�� �ND��#��ƅ$T�mgKD7q�p�~ �+�߆!��;�+^�Eы%8��3Uf9�����}��0�]�c�7�R;�"���F#����������C�Y7�w�=������f;$b���y�����g���O�	T���n��7O�Y!�}�.C��+	׳��������9i>V>VOi���l`�8���z����v?�@X�Vgի삯r.܊�u�
��96ػK[�8e���&ǌ�,�jb��K�%4��j�Zը��B�X��ߘ���dM��o<S�s�u!8*�-�?	���QB���7\��	d�M�!(�@I�5pD`!l��`v��-�A�V��?d����/`�_F��h�J�:�=��o��Y[\/�7�b��ǅT�}�����O�K��+Ƞ�Ipz��Й�E�#��7�	{��k��u�����;��|d���z�37pB̂a�۶�J��-�l!w�W4�$w�}s��ծNq�V���F9��7��YBO.�\�4�o��N�V��is��pe�D��/��b������K�CTpqb�[\��� �fń�yVV9�b��� ;��zk�y�X����ҍ^����ٓ���4����y��1.gT1�~�J��
qu(̥�g=Ļ��1[\�4ȁ<r���4�^��1���G��V :�suןmx@d�Yj�7��
d0���u�������E�?^�\�È�*���[��[pm�	8x,���dN'�Vyx��}��i�8�#L�����u�����8Qu�v�����豣�(�A�m��Ia������}�t�ݾ���oqu�pͳ���ie������r�Z� ��~l`r��Z�m:�H��F��.{Ɖ:p]"�k:��P>��R�[�C���<������G9t��pc� FVc!����c�M{�@*��w����pu��Ŏu&��!������S�����8|�KNQ_��1D�@$Y�Q.`�Qmp��P�H�p��IJ��-MP٪C���$x�Nݳ��+��|�vh8��ryul�`�(�$pU���)��`�(&���F������ܩs��+��3��5�U�V,�a�67�
��.I��{��r�?�q�E҄aI�$��s���o��߰��Ω6h*��Fw��������7q�'mJ����o%PN7H�Н�ԙn%��K?�t'��o��rM'���=���|��s9~}�Vs��y�h
N=�PRx6�"|b�@��$$w�C�� ��,�I�A����9�n�v"9�?Z�:Z;�Xy����^�#e���>�l,�l.s���?y�s^���yp��yʀ�b���)[{�|v��M�Y�mN
1:�)�r$�ivr..~z���с���۸�ҝ��2���+�g��d9It���,;��Y�ߖ���+�v��y��v8wG�P��B����;�!;6S���q��[rY+i�V�ڻ|Rl�W���@ɸ��f��%P׹UL �2,>��������������rszZL�Tz��\�̑����d�u�n�lCn%����X�Ȓ�VBi2R�\1@d���uTpX�.�CAf������_�=��n"�om�Cd9��8-�1�ж�f�j�!tdQ��8w���!�)u.�O�+��[Q�.
9��Ӳj9L�7�ަ]T~�Un^�,�w�}�ϕ?���X8h�1(87�pw�\�C1�_�[*gV�Z�	�23q'>$8�������ɟ&������x�]��x^o�SIa���p�.����#]P����b����������nŒ�p�����mY��w0�;��Wy��M��D���I����?��?-W�ވM�n��PH�=��3��1���9�D�]����zH�I}Sh����!�3�X$��g���nq��틤�k�q��� �S�l˙�C7�I���ř�Y43�(���V���P'Q�N}ýu��rzURS�P]�b�"2U�F�7�ˑѣ��k����2�/��"`�+����S	�I���I'��H�h7>��W��t��o]�g����߻�(j���$��
b�����/qGk۫�ݷ�Fzjr*��@>� ���D�rm�����٨�w���Ȧ_��0ߙ^��2�� n�x��������@���Ա3�[�0�����ʑ!�jXG�B��d��|j�*�;&���!W������L'��]�нn��v���9Y>��w��xf�8�gl6F{�˹s��x�<~��r��s�����^��W�"WDQ$��A�l]��
��PE!�ho��{���w��a��q���`�~���p����;��eu� ��=�\��~4I�����WGa����
|*�Hx�7\�껉�꒸}gx�i���3�j^W����}sK��)�엸i���.��Oy��ڳ0֪ܔ��lP �C��N�M�/6Қ���
$���i�y�	J���~������D��W�T�a7��=r����Ѳ:��{���P�ü�~��&�P"d$�W�"�z�I���-c�����9��'k��f	i�z".p���>B~�r��q�Q�NZ:��J�y3gyj~BI� � �W�j_��W�Ӈ�:���w�O��x�|��ϕ+���:��n� ���ݶ*;��Kg��m���5B�8�$\�.��۰ģ�����X'��L�f���X�ż�������{��f����nz$�P�S	��m�#A�!�ފ��C\6��8�Hn��q����U�19�,�i�,D��j�1�?��?���W~�����XH���c9�ti�vq��w%wX{�Z7GE��-OA�Ր��B���å'XY��q^��o$�z-7�|���r���rmu����2���7f�x��N	��8¿r�%T���@��;vŬ�Sm[��E�bI&�Z�Q%D*Vc�l=���_�T^���+�����?U>���R�c���f�GV��Q�����m�"���$��$�H��G���o�mx:����.rɠ����t��:�2w?��J����1�{�=�HA���D�C�×C��3���6"9\x��?�������f�~�q�݌�yq�x˵>�|�	��~����o�	s+�y��������s�|(�^���в'�c�d���	�3�4�Ԡ����v���u��%u��u.�����/��bl
�K���433W�0����r�0��%A�z]rdvv���	U���������gQ��L͔���'������5�E�Cr�3j@ےb��ّ "�hu����K���e<���W�/�x��t�Z��X�	�7�
06;�g�7��͹�scas +CW�)�ݙ����p��;�n�Ww@�p��
_�/�t�A����G7�Э��2�ωc/�xx�z5چ1�3��9��|џ��(q����k�ч���6K����(�����G9�Z�D�6�[foqn���4� ���Q�@u������6�*���B�J����䊇�7��� ��u�2���MN+%����rm�R�m�pV�+P=�+ޑ݈p�h����Ux�����ӣ�f�,3�`1�=�^�/�˭����semv�����~M!��N@�4B'׆���*p��l�)�C3�RȰ|�E�l�SP!R�%�@"����Ы�6�@(�Ǡm&��������{�?��EW'�:;�� n��D���M�ׯ�o�>ӷl/?~�DؖhPW&Y���I�:��]	�^L�q�.�Ѵh�qu�O~�g�@�_��B���rQ��
�����8�����`�:9�8�e�9{r�v�u�v�89���v,�$�5�5;�.���)3��<!�Ц0�BcA��m1-HOi���s���@{�� R������-N�rG�m�^(���*t�k�9���enj��$��K]��n�W_<_Μ8[�������/B����֨1�C2�傰Hx�{w\�?>��ѷ⸎>�>���7Y�����9V��.(�����k1�t��a:[�;����{{�_��F�� ���'��1>�qژ���I���.@��~r[�ɩt�W�~W�.���\�NXݩbz�:1ar�U������+��e�~�B�<�2�|��������=�=�`�eD`�l�GG<{л/����M�£���`Yx��V_�N�k���Ӻr9��tX�EMm�Ё1bূ]�T���U\R��!'/�.����L�Go�o�������3�q�do������<#&���C��,�;i�~�t��&a'1f��~g���δ�[:G�A{lR�Q��3������G��8z1�o���M���#l���Tv�+*�99���M��`)k��h�qXAiu%ʬ�iz;��@|K$	 ��[�t	��9|Y?;�������{��ʅ�O��O��|�|����Ӈ���p��5�U�O_A-ȁ�twޯ��vږX>���[�R�S"���P��z�0����j����xD��Z	Z�n!���'�[�c��hUa�dvy$1slX��D�_�*7�~���w��$6�k}hHʟ���J����[�>f�fѐ�}��}��L+>�	�8�Ig���^�y�����/=v�"�i3ú�    IDAT �U���k�sit�f��E�Nό�7��7q��9*����=0\Ua�"�z�⎎5&[]E 8�����8�k�$��0�m�,���@�5� �@����ջȗ|�5�C ����st8��|=n-'�����_�u������ϣ޷f1�Ef?:v���2�Z�
X�� ��H�؞�N2��٭���v�7��[R����TL��G�:���/Y��%�A!h��c#�GG2k��1�1	��1��0s��ђP�k��8�Z)�_�\�����l�{�'s
:ê�C�[$��wϰ��	�k�a�'�2M����,�g���t��;:*E)�_��,�tҀ�]�5��v�|L�eV�C�l�ݛ��Mܫ�g�8�v@��ɕ�]��z�Jf�k��oSQ7�J�:+nc��6'�9�����o�3�N�z��(2�#��۫���3�~�)綎��^W��k���I�W��g�?Pƹ~�{$��<�h�=�-����5B�\*�=�,�l`qG=)|{�o F$E�Q�_�.T�Zo��h�f�����ǎP�4v�vR��͌-\}��E��l�;m�V���k�[,V=W���s��P��_��r����Ԃ8֗8��z/�]K탸rgRQK�0�w�~�~	_q�8���7��UmȎ�p��0���*T?���e;�vtpqI�J��[{�}���rWo��qnr��~�#)=�Py�W������:�买U q*j�A�' û6V���1,Uߵ��jK�=q�����{*��u�1q]���8�)�1�Xj\^^�ʼ�Q&�p�|�/��q������Q�X
*��'~ۏ��ZъL��dG:mV�RdmU@�#�ڛ��8w�BB��(���3�5*�o%^\[�5�י@�[t�5881bċ���h�	��j�*�`X6�z���Wb���ѳ�y�>���,M"�@��u��4� �0b4���)�#,�Pߞ�&��*��T�Է�ť��N�藿kN���9_�<2���Li���\���ҁ
	����#��#�8���o��M�1���B�@T�B匮 ~�ӟ�=�w���!����R��p��r�^䅿=4�@��	8�@'����N'��|�r��(��	�ᳳ��� �����G~�Gʷ|�{��M�e?ʦ�1�D���̵�r�vc��$�z�v k���F�h�	@]#��#�m5Xyny\�g[i�Wީ��@�|��Z;�Ҙa"�06>`����ȝ�˗����Z�.���W���>,7�7��>^ڳca��.x�Ս�a�a�2B�p�_x��~r�7L���~���S�y&���8�R[��<E��l�oEH�9��]��1�ƚާ��ea�t�o�~��?]}��^����'!}�W| 	��9����V�r �z�(�Z���I�� �hq�S�J��-_������S�
�r�� �E��c�t���Yn��I}������s�S�Ї>T���/��� r�Tg�f��'Cf_Z熭��r��58�������!�@X�ǗW�P�y��u�Um]�(KH+hX�]���u 'J=�x��υ#���jL�jh#��ln�D�k����Y)���	X����K��Ƶ����kat�˽�aC�]�ZtU�:G�g�8z.#r)
�b�ήq"QJx�'����6f�ڜD�针�	�����myvj;^&碘�^�vS����I�,G}w:ӢAi�1�60v��M���n���Y����3����~�޳O�ɾM !"�"���<ATP?}�y~�� *���""��""jD6�����ٓٷ������NuM&<qC|/3V�s��[�N�:u�)�*��@�f̘a x;�Gf^�L1���p��0��*S�*�@)Bj�_=��}2��5�� �@�>��x��pd�����m�s?��O݃�/߇��aG�V[�S�ftӛ�E����d���0٭k{�mm�*ca�����Z-����ڱ]�M�1��W�`[حl�c��k�������]���Q�&!���m�ZI8P��.ߪur_��yb������I�_Ӈ�;�l�k�`m�?IFB�$��aX��i lh�/B\�g��B�p�>}�b����p/��<Nm�lH��Ƞf�H�c�h�g\c�$#��1�X,H}��g����&�S���(ekY*	�aS =F�o���"�}(�^)Z�8�j5r w��ÿ/ @Q�O�eQBCC-�5��&�A��YS'��l����>[�{�J�|��h_w�.v�fN1�f��i���]�ZvS�dqS;�����۰Z���F2'Ys���%�B��T��nR� "�A��t��#:�X�qc�\^����lB�����w˖��e���n�ZQ/fb$x_��̞�p&��$|2�30�g�&ZA}����
ভi��j�жCi���C��7���jy��,^��V`��<`]q3�3c�,# �i8��H�1�Y����Vk���/ܬ��(�SӵЊ�}�Ī�@E���V*��b@ݹVi��7(iQd��M�J�l�J_����>6���K�c0�9
�����>>qƌ�V._��~��t�[Np?�lft2q}�6�DeЏ��aNGsÎlھQ����."�W���+���=����y\)�s?�q��b�䎢��ӭ\�B&`/��L�F���g�*Q�35՘hOL��q{9)~����� SE�o3G��N��6��B;���#<��q^��C<��e�%~צjM
Ħ޲O�n��p�W��
�	�ia�=�Jz"��WHH���H����:/_��-~�b�: 1���P�,篋�s�#����c�$]�Oh0�6��
fqD�U
?��Nު4�5.Ƹb;�N�C��7��l��J�%H�=x=�Cq��ޙu-k_pW}�J�,?s���s���ݼ�{���R9He��)7�]m��ݞs�q[�U��ތxou��8�-p����e�ڠ&t��d<Q�~w��܅��HB|g��8i	�RK䇮v�s1U��9���[�P~>m�P?�����aY�څv`�=��N�I륞�O�����m�R6��4���%nSIgFz�I�`�`��:�5">Iw���� ��:�#�-��	����:�τ�C���/oEKATj�~��x�buS�N5=�F�D�:�dU!���*E�1B�����Ҩ�w$�o���#�.�	i���i2�X�χ�T������^a���+K���MnӺ�n��M��w�[k�Z�0���1����C�/º9��\1-4���II�T#�+�љ�&Θ,=���ս�q߿�F�ZU9��ؠ�E!�~��a�����Zo
�,���.~��扨��6Q=���.�X��-i.J��w�+�!�V�Yh7��M�=�.�!�ɕ>�х�k#��&�MB"̷���я��V<�ʝs�9�U����kj����%*�-��MPs(y��]��'?��?�|��OZGS�őz44��X/���h��o�Q�Vڈ��\�;;�����ۨ֎�v��P1��� `� [��9�Q�c�c�������#���o�{n�*w�'ϳ4k��]����gO��������uR��?g�\7�Q�2 !'�N��ܚֹ���]��ܺe�$�k�� UN��U[�
�&E��-)H���Tn�CŅ_հ�E���H�6�@�Şb�`�ޒD2h�<`����/~�oB�� �;WvP��cI�@t[�R���������l��t"�T�E��ʟI5"�?^�$K���%K0��97�V��QG�.��r9�8��׭J@yp�a���M1��c{�w��i �h�qa�hL�����#�uc���1�/6�0��â')6�<���'bF ��v���s���7�-�~R��*u�C�R�!�s����s��5:����ջ����߹��G��0��(ȵpI��d1�/�v6P��{
�ޒ�(_N� F"����H�Jڂ����q�6UlcE�1%ڏk�p�2��	�½�m�}�INx'\I��̨SFbQe�$ �j�H��N�ظq�o?�s$:y����=�z��e����/��(b7pP�v6;a�V� ����8M��8�]��ֶ���JZ�B�^T��T ��{6#�Ѷ���ѭᘦ,◑�!�_��?�-^3�#�n���#��CHMuX�@�L\�cRN�5�M��5I��I��2i�������X��1u��ݲc}�K��h
���	@2��KV���`p]8�g���"���KPZ=C�+EЫ����(O�*ՀfЇ�c��o�	�38�!��;�b}� ��ə> ~�@�ܧD{�l35#X��0���_<���;���V��^Jrx�2reQ���k��7�p�[���5����W�7vҡ׬_�h��-���/���"���C��l��Vg�ae�o}K�w��vڐ�ЩPn�Wփ�/}�	!4z��5<~�=����A���"�����������,�_���峸�ܧ��Q3`��@E�>���x/<#m~�p����.|x��)���Oؑ�o�?���������^h���ʇx!��h��Ti��$WbS(�9�|��߫�t��o��X�j-�i[D���Ʉ\��p6��N/����ښج�AS�5��w
G��\�B�^﹈�r�* �Q$�Z#3Fu+$�ť-3=�a��X>"L�#��C�gP���~� 2>��wt��<'���yx��t�H�ѱ�m�m�v�#��Joy�7��mra�@�!��^ yr/��o�B\~����|ݩM%BE����:�3�#=�>]��ۛ���Ӱ���< �I<>�r���z�z�Зs�����	�'�n-�y�<)̛����	$(-����pM:2b���2vc��bNb�R���_�����o��ں�8�=����f���_x%|uϚ5˝peU=�]��U��AE��y_܉�KF��p�6��x�w��>(�k�aT�^�A�U|ރ���u���6��H����,��
K�(�u�x��餁�ڋ�X�J��J��r��C�!ߡ�_O���	mae�1V}����O^!.�Ӷ�T�)�[�DV��t����P<{��'�hC�M�P�>y�Ev��ﾯrW\q��1s����[��Ú��[�mU5:��8��r�UϮ];<���tw�;vn}Mm�2F�R�ֹ�J�E#+ڧ�~�F\��fw�A�ʌk����D����)ЎΥp��ꛡ��*t�n�b7C $\���� �͈V����f��"U��a�B��[�6ќ
�Д_�	1�'_iWxy W�����y�锇ϋl����w>! z	��(��6��ƞ�C��w��� ��@эrkVG�4|L���ǋۀ��ߣ��_(���{ 3��4l`)�z��>@����z҉v�rq��s��3 I�XF�)�,z�V,_:�������`j�TxY��c�#7w����6o<��d���h@��߰~�I���U���f���okb2
��0�;�dxC74���}���ǎo��(1����g?�'��C��	�����j��Y�z#�3��"�~�wLLi�l�X�6ګ���P8��0$������h׏��P~�tBk��=��c(�6�x7|H���9�x�
y�+�x��g�P�@��ޡ����Fe$Yz��s���Ez'���/:�K�^�k
��4 N�晪ں<���_������դ���ƍyC[[{�SҢ�9V]���:}��ҧ��.\�����-]���ߦ��v��14J���M���#�^��>�w���\+o�	�ߐ�k�> �D	��sэy)&<;�8Ȧ�_%����-�Y�ٚB)"5b�m``v!?��(8��N2�?(���" ѰbW
�hv�����wf4"��*߭a�o��?�j�3��&m���feo��� ��� ���K���	��v��$/�� �+�o;�dw�g/27��W<�>���j-3(޺�ĮԌ�r⤉9�<���ܴ}{W�x��r�]�m��9��L�tuA� l*͈c�
�u�;����l+dt�YD��^@�ݠ�����M��ڠ
Kk���yp��SR}�,�w̀�:ȏ"+i�;�� ���K��<C�����A�aU���G:�ҳ8�2U�D�	���n�o��)^����!~�P �U��B�֞v�;�	�r�W	����!� ���g(3}����������n�=���Y�����K��!Qv�7�|_��i��v�{3�?^���&%Aa^2�\p[�ZZ�;v�ٽ�}Is��Q�s�H��l��
������>�h�N�u:[PqӒ�$�X@y=�Uq�dƘ�%�Q�0儂��*�k��`q��D���aZGG��#�H ���g"2���sI����u�Z���H�g�a,`l
3Ċ«{����G����TЕ��E9��It/�ɢu֬Y-�@���S�eq�yi�o�)92�"L;����VL��1՟�_�#	��@���o�'芪��D� �pv�ڴ�|m�(���:�Xw�g�w{/��m�l~�Ε5�Ö��C3;�I�#]�H�x����2���ZV^*7�Qinz9�������M.�w�[6o�?4 8ؾ�3�<��pS�Ls�g�v�-RJGY�F�0�v7��~mr0���(_5�"��X���8j��`<3�*O�#��p�ƥ�hX���*��.p�+y� �H�lt��k@!�cpϏ�!m���(��=/Q�0Xi�<��Ƀ4ѫ��8e������w"u���׿����/����g�,�A	��ߡ/�o�N�P���wW�0(=��>��O��|<fc�B?�:�6�����I��)e���s_�Ǚ�g�5kֹ�|����dmg��i 0}���Y3۶�m}$Z�<���QnY��@-֟��wQ��ڪ���2�jV���\�b
\�(ӹ���k)UMp�z�{ӛ�h���Ԡ"4 �)P$�*�N�s�0��������i�Iƞok�H�8hh� �F)mu6�E/
Б�7�k
���xt,���N:��=��i����W�SWD\���AG��l�|�����g+�myNOz�I>�{��&I�{���3'�W�;���#�8�����i_��,}�~xR�A�&� Tږ2��b$��7;���*7m�;>�~�N�p�:����k�ҹ��/o���V14J�=Xm���Ƽ�ql?�|w�UW�~Mn�ܽ}�K_4}����t���1��@[��R����l�䶭��iT1����ǩ�y{�ho�~$R
FGұ�ꗬ2���;l�p��5��O��&O<�[�z�Q�5�AP+ާ����AB�t�8��À ��Q���:���Ω,��-F�w�а�$�ƥ�hd��} @��=y ����8<#�.�	W� �3EB�)�����y�T�Ѓu�ƹ6�_~���ww��wՕW�����HaG�.������|��2�#mP�bEhDl��U���ȍg����>*�=Q�iO>��jm.��p�u�}����B�F�mG?.^�ؔ��򖷺����j���;����W�=��P�G\ۨYA>/3�����ػM>��}�Z�^��~�7>Y�wQ���e������ܨ����\s�Q�{�ױ�y��w��4�c��g�8��FU# $�0�
-vD��������_����V�����PT��0x�@��i:�8af!:�(�ژ�����7H�,������	K�i�{�+&���?:�}�򯻷����_��Wv�4��^{�뮻ζ�i��jX ;���U?�rئb�P��WU|[C��c�%><��M�tc |:�q/u��S^ ˇ#S�;D��>@����裌��r��c�=���/P��V�[���|�?Z=�<^��w��xACQ�b\��\ݘ�/=�賟&�%�����G9.ױue[k[l�dӔ|��( �w�,�Ot��'����u���曭�?աMXg����;42�Y�CP�!:��E5q�|�t⡍���(
��ŉ<���.    IDAT%.�f�G����%Б� �b|A\���'�&�Xo �)_1��3<�Z�����zL�֬Ycu>���ݯ���hqp�s�,H���fР���o� �߁d[�A�E<��C/�6����L�e�.�����ϭdXM�1�#.�ǋ�D����3����=��#������K/�T���;�:���M����f̘ZЦ��� H@����g�Y�mx���;���y���l\�����5+����?���鞆3**�E�C�bR���}���w���E&	�M��j��y���f��F�q��׫$?4�P5�2��K#:�1��s��cu��z	p	������ACU��iO���r>��~�&O�*��lQD���ܪE�2ҭ1^V�D�X,�ʆR�FF���$�����~?+8:��lF�r�n�H�}*�:��a�%e9�$�<�� ����-\�-ƾp�76�\aWT4k/�m�%��LD{QOlߞ���Sqi/��x������\�][����fs�{���I��<���OD�5"$H�&O�T��K>1P�~��[��X֊����_���g��w�x�#���LM,&h4kD5�Q@�l�HTԨ�xB(��;5E��Qg��ޜ�s�w�w���T�$\{��M�qM�4�\�q?]k�V f�� j���#�'Lh���Z�l6��q�[�l-�>{/4C�O<>�tu�
��>����`ĵ:���L�6�\�M�6������%PM�mJ<�Q}�<� �Clk�|ł,���3%PV�V�
%fF"��hW�E���;��$?���ޡ��*N��{��xCפM]!R�3V����np��w�6�5�0H�������96�͛z�ڵ+���/˩׍�I��7i���p�5kW�|��m[#P_�Fcuε,}n@�i ��:���c�ns�Q�.�H,���J�ƯQ����6N$CEC1��kz�, ��x{G��� �iej����R���!��)�t�kש���S��� �Z�\��2`��z�Ϊ5f&" �C�K.�� �*��cI�Ԉ�59�(,�j�~®�&�ŀ�|�Ȱ�2��r�f�@)yT�F	��D���
�;@*vN�!��A͕$�`��q��<a��C�@�tY$C�#��6����GlL�XCm֌K\T[�',W�C��3r�F�-&L���k ��|O�s---���Ǘn؍��cO8���r�-�t(���sPǤ��8��JkQ'������� �dƵt�)��yh7Q�1Ѡ�5k�{�ey�,�'Z��qXV�#�b
%�D:Kj��%�R�S�]���̵�~a�:��r��J���+��j���n��vsO=�4��u˟]a�b���SO��ɛr�'�ʠ�J���nӛ��P07��lJss�V� ���
�ZIn �� p��ʀ���{�����a п��A/W,ā-�}ڇVD�mV.7D%���&�.�\���u�N���ļ�(`O�P(�т=c�@�ȗ��]�:���׃�����'�t��h��x:z��GVJ�U#���8�U���o:��LWϵ�._��~Z��8�"0m4m���\:�Dj�:ₕ3���l�dĚ&Ŷ0ʹ���$���h8:
j�t �y\���n�k=`�uWf�h�C\)�ػ(��1u��P���E����$�$�㘖0�=2T��Fٵ�I��5p�� 5�A@]&��`�g��α�خ��j{����[�� k � ��R��g����͂�z���\J�.����Y�ԋ��} +�I޴ruf�4����f��n�?����c�-�F\ڂ6�p�M�HV�vƫj�(��)t^K9D <I�����b-^��I�
.��y�-Ʊ�2%"DW�$ �`�k��!��Ih�چZ5.�����Phס�]�N$$HS�?jx:DJ[� 
�#�M��E�i�0�����Y�� �5���=�z�f���%��QD���1t�����D`�v0��pHhc��N�(-j�Y�1Px��X��Y7u�4��_�r�/���0��Ǝ������'?$K�I�݊O }�J~�5�-��5����@�FLh�l��%T��}Zp��}�8e�;��jfEzB��5��wҧM
��7�[j�0n�
{��~��6�_��K�ɿ�׶
돯Y��
]%	Ih�����y�鿘�J^�e���p��]j�Ff;������-��M�Ċ�)M�I��]�Ѣ�]6��Fי3�A�ӭ6�.��$^b�t��Ӡ�^	�`���(W���s�6�$�|�E(ZlZR���t ¢�GBj;�:
'�E���O��۸р#`B��� ���>q�JLG!�G�.5�p�#�p9Q^[�T�5Do��c�2XX? 0@�����= N�JE��0����g��ͱn�]���� ��/�-b�4mH{�1��o�f��d�(��k3"$^[l(y23M�>]�GcV��`�x�DM��K����.BQZ�\�(�\`�Fe���W.lٲ�$�R�������U3�l�u]}cT.jeRTZ�Z��h|,3�F��(T������RZ(�t��`�|&L��R���~���M���0=�e�K' ��h %+13�@u7]nu >N�i �CN?�t���-}(8~����<�V$��g���"��Pb_W��C�7�����كrM<�H��1 "6�o��)/�@�'�$ġ����� ���m���6Ȉ��A��[�Eۥ�W3'�����:��9N�1�͊��C���ؠR��I�5U�d,O��w<3n���כ�E^rׯ_���/)BY%��?�����mk�����\���k�xݢlw�ɢ��Ӷ�nk��a�ZnLݦ#.P�ǃ���c-T������f6Ow۶n����H�; ~Ş:m@i�((� ���\s�,�`��MA�+I3�Du�J �)Q�7J�g/�"�N�P���QZ �a_��݄qM���4��*�7ʁO�dJR�'�ڀ�A��ZL�2Q�4KH
���n����OSovq I�R_��.�jm�igX!�)j�3��0��8$���?���)������(�~�d�^���꡶�k�'�� �L̫�]/�R��J�T�֦�\B'B�$��=.���P��+�z�K�m�a̸�wvl+��O��{dk����������G�����/U���Lx��5���>h�W�K�To�^%��Ɓlv�<�j�.�%a�ĩP-�Z{ń:�[G�3�|���[Sʗ�s���/��\�Z�����h���AuZ..W�%]'d����fT�xA6g�~�m@�Դ
�:ƪ���_x��c�ug�u���<��%�?�$��{���c���QQ9ׁ�񌝼s�=�(ã�:�x}�>��Ύ�ݨ�҈׮]�.=�B��H�H�2�~JN�I�����%�a�A�U�1��)�CY3�|����O�W댬6��4 -�V�*����KZӈC�����O�j�:Y�¯�b�T�Wi]���:�oK�}<�7�5�*�>>ߨ��m��=���6+�+���r���m'�,�硕�χ�C�L;h�\�O�+���@�&��9V����+n��K�I�7Zn��`���c�ĢX�L)��EK���.����Tj��9�>����\����D�8քGb��3�ȵ��VJhƃB}YC]�ĐMn�n�ݶ�[���𗀊 8���y�Fu�>ޣx�4<.W�z�ᇭ<�8s�̱��,����B~�E��A�ZҜ�҂]+Td���f$�-7k��K�s���<:�����{�ԋ���Tߓh}��y�0�K�j���r�C�B�p#wYn�>QP�JKg��t�l\9V+�A~1R����v$uPO_n�]��A�#MK�������ܟJ[�=��)�
��w�t�#��Y`a�klH�/��/!/����&���*^{�wݛ��&��J��U0�2l ����;�t�ˇK�X ��qPK�  �C�����Pe�b@��98�%-���w<Pn�!Ϯ�7s�L���'#
e��9�`]����wG[:wĦ��Y,Ԓ%:hs� >��I�Q�yqsjr�y衍A��ǻ@���!�r�O s�����r���sҢ�ob݌-����X�G^�*,� h
�?|� 
�x�� 4���$M8(nN��=t)`# -�yo�	%��yy%~�|)�>�校�(Q(aӦ-�����'� �tI����*)Me��e@��������6Z��i?+Qf$�NKڗ)$"��w�+.���۟��%-ٖ���x;�m�s��Qn���/>!�%�}ƿt:�2c@�=�U7^W<8��AS=@%.�?,(	��|� ���Y�_�$] Gz��u&�!�ǳ���fj�s��@�.3T���hv@2q�%���@�I��!�!Mޡ���J���^�k�i��6R�F!��64��+
6 �u�@��o:�3@`�=PE�lPN(;ׄ�|���i���
p�C������ȼ�=*�lİ���,bаI��t�g�P$�:3^"RN!�Ʒ���N���/I#+"���X^P� hX$@Pz��H�C�uHC������"V���g��E^��ͥ�3��f�pq
� 0A��߀�Ai��F�u�*�;���b�� =q()�!�]���� ��&�O�
� ~�(6~���9Zw�"��-x�C����^��8����klG��B9;ޡ.��@�2V��^Ң����;#�Ϩw,�#q`�Q`QUTI� ⷝգM`3�>�N���`����߻Uk�s+�[54` -T�h�u�Mۼ	@n�YX�[�~;*����\!'~^�4X�p<��g�5!,P�@+�u������}�r�!n�=�k �8`�ts]+�p��Q%���pV�6i�^�-X��~�h_t@[ݩĎ����1*������`�s{�၏n۩(��FY+�o(���u���(p7�t�Xw̴P���Dx�B��� eo�%&]@�~�9���f�(��HCڥ��L���,ΦM�LJ��%�}X �֬^m�ed`Rn�3� �*�;�Ϟ�d��P�4����iaT��gkOt�����m�1$� &	�u��Z����2")�W�Φ�C�k!��֦�	�tmã=��
Y9���Gn,����{�<w���{�9;��qh+F�ZB��cD�v��}�_@��NgD���~kQֹ���H	y�d��j����;���[�l�kٸ� �gH�P�B�	G���ni���a \��k���$�KV��i��>�ܭ�-[�g�>*����%��$PK(��ν z
�̢�{H0��h����=��Z75���1��@(��G?�Qw�܅a�x�7Ņ�By1��;�-*��72;�Y��ʿ���u�]v�{X�6꿇�v�ʐ�2</���}֝w�y�e㝔t�}�)�g����neb��AO\��&��䟐q��wΰ��W��^'�C좶�D�@� > ���������Pn��vQd,�;�F�ަ�[���S����n��V-l[��>�Ԩ���M�ɂ�O2�3(�V���� ��<��Z8_җ:��w�˽��T$��,�Gy�X�F�N�6��m�̰!��O@�O �(�z��S�l*���_�~��IF�Hν�-/��Z�����X����"+�&��� �@Q�Q������Z���}��ƣ�����������S+�'d�7�|����0^�c� WI�Vj��e�Q�a#����tg�}��C<��O>���'-(qBJV�r2U��A��y��J !���X��Td)<E˺3�¨���Z}+JB�����c�] � ��7��K��Ve���;~�K�z�7����b���� �w���<*]f�@D4����5�c3Ė`�N>�++�ɀ���+\ˆ�n�[�w������T�N>���Ԅ{��%Y��gZ�SPo$.Vv�D���AU8�W��Zf���~��!�Q�Nb/�� �`TjK��'��ԓ �o�ov.�7(��-���7��	��	X���7c��in��*v*PR����S�-X�������T��z��bl�u\���3��ܺi�啒,��.W������vȓ�*�f�D��U�F$��Rht���Xr�ع5�N#���2�
���
� �5$>fVӧO����O�4��h��g�c�]G]���OD��%�#M('�� ��a0 Ρ.���0{�"��Sة<���߈zϘ1��J� 4���4y5]>�'��*���5����	�QG���{-HΈG55ː��+`z&�3`$ 5X$$ ��1�eцd���V����~B���S�.8�A'�4	l��f@��d��>��u�ʚ�ubs�u�6�c�9h��e0���E$�~Hh`oX� ?��=���Qg~�ڇ"�(:������i����r^��m8bDՏpaԁ�>�6�[�i�����t: T�5Ā6  ���o>�\9�����($�2*w���b��b�
wđ��H*��(�=���6��#�x�M��}���~��9�����_k[��v��@o ,���x���Pf��~
;���u�;��J�(���'�RuM}�������ʡ�?���x��m� l�`ј���1�@(�"���$`���|c'���*�'��B����jݺ{�<ȏ��/� ���s�.鍗�W�0?'�Ri]r�����	�,��gH[ZZ�y}�k
�>�t)y����y����/KUM��m��,�)���/�(`�Σ�rwvV�(�RbCl�� �e( ��%�;�),
��/��t�����X��J\��Ip�;���C�q�'V��=�N���/����(�9�Am�sf�u�������#�W"��_�t�׸f�(˖=���t�^R���aK&�V��Ϣ�:�3���6�uyf��5
���E�=v��˥74s� XP9~�0�
`��A�s3��L@��eҤj;7���i �@����s��c�I��֜��!�m}��GO�.%i�P/}�Q�#L�1l]{{���?~�>������a��Y�e ��S&ҁ-!P&� [FK+�	�X1q3�L�.�Q6yaDV�/u�6X��f����=z�N4�f �N4����Pp�s_.(��2 ���eQ���ü�։bZ�:h���3r�\%]���z�׼�xnxr �T~Pc|Pm��,qJ��:�Y�ʋ�"���&�-�T6xd��A'cK� Y���C��_�.���喊8��/�mR��SH?�t�Z\D��V�]�ϨdK�2M�ɲe)&����� jz�h�� 0P��ҷ���ϻ׽n�4��
hC�wP\dɲc�)؀{��'Lvλ�G�򁠴��K�kP0S �A:�T�=J�����Yљg���~�;�)'�b��%]�9(�^��w�*y�7����c��)�H����cN��w����-�@-`se2L�PPm��xx�š�o~�ݱr������&��n�M��0 )���CZhb�3F^� dM����W�#`'z��m��D{08�9�S��4i"�����/���c@���H��9����s:VDe����RJ3�����2V�]�ψ��K�MK��,&[�7@`�
���4x]��a? $ �j����S!��}�C2 h��y~`�S�'�m�3 ��<�YCy�� $�	�}�zSV*����a]/y�>	�G:@��;Pmf ����6sDc5X9�0��:�Npo�8 �U�j	��8�{6�Q��\�o��I2e!S�u�go_�͚���r�B��u�P <��q)���R�*H�����v���%����Lx�U�ͻ��|x7H�"�6�b/��_�FMM�ޑ>yF���w�.C����NU���l�ǔ��~ݳ'HM�h%���۫�����r�Hz�G���]?�Np���x����Aq�� �3(0ψ僢c��Vrf�ƍ7���GR�1�L�8��v�H    IDAT7&����2�y?܃�����M����rK�5�<8r�@|�!>� �0;q����r9�}J�z�2BGL�#�:uE"�f�yM���G���I@����6 ��68#�����s|�q���k�I=��qFώa�<�b�]꨸H�(���f��A�M��a-���,�`�`C�Kc� �8��8���e�.��������+g�x�n��[�'+w_^o���W�eg�W�Gz�����d�b1��
-�1 �J��D���()��f�
E�
��{(*T��p> ��/����_l�S�õ�܌��5���\4���т�5z!Pk�4R�((�ɡ��r'L���}��
#�:�����S��V=gqƌmP���ޑ&3��|����v"�Ê
�C�������R.7�dݣܲJ,˩���� ��e��6`� �z�g�����u����v�m�P_n�N��a֬Yn��*��N�6�އ�ت�K0��+�ѧ��W�����s���������t!�� ���Q,�?�Ye�����#�}��,ű��@}�:��� �M07åڈ	����/��L����{�]Jz0
� %�(.0A=s�����~�=����C�����9�'.�q�i��3|���gq�mc|�
s��g�T�0�
�xoX��UU㪙CM[M����}{����;קܜ2�bi��s*U���ŧ�d����R�	��i�1r��F%�[[ӹ�s"��4�8�� `�f���Y�@�=��.;}ޱ�b,
j��i������m� �
o�Q����o~�'Mo�aM���U�V�ռ�sd��*^�ޥ��L�ރ�6m�`,�\!�V��B���ꡛ���r�3��h&��{� ���Jp�K��qݸK(AY����d|�AE���H������v~����ͻ8MFz��I"h�Э^��s�a;�l�N �,6?���L�ì �vX|:�ޤ�D9ɏ2�`�r��x�y@M��C�>�F��O��Jԯ�%R�K92Z*5F����r�?��Rp7'$��PƅS5�  P@��*I?X����:=���E��ɍ�r��!��/��s�央���������Zy[z�j��轐'�JLF�-�>��������7q����ex��V-�\�6r�f@ןH!& r)��M���F)�kd�U,��IPP��/����a�sB0�7��?���N�c�9w��S�����:m��#���~^Rxf��'P߆����|�m��T�����A~�,|'�� )UyP{@��4Zo�p~D�lJq%�)��6�T$Y����m���.F�H��{��M�:g����7j����+iȾRȨ(S	 ���&��5�^owK]�v�}w;�]���i�C��y���FM:% �3j�E�
�<H<�J��$����}>�v	�kn�s(���9���=�k嵯�&�m�( M\Ր%ff�x�H<�L��u�bq[���I��W?�w�
�E��J��H<p��;(�Oj�}>��zx�׭[�+y6σL��X` ��	��7���N'ع�0i�'����^�V_� j�q?�P����q�v�[[��Ӊb��,rB��u��%֡"�L�~���6ʆ�I`ة$����x��'��?�+��`7ؒ�?�e;>�+��b����WG�J06P�z� AG�A�uO���Y�Qhv&���;�p�u�>�Ry_�e�&�enN)�Ydq�4@"^����G#����%����n;(=~�V H�X��
~���.���,��?�pw�G�3G���@X���}�{F�;��tD��')iB]aCB� ���oE��}���n��`�1�� z�D�U�7-���B\���s�Fp�_�$��E��~�'�C ��W|���zM�<���o�E���/��G����*9��=�AP�[����tn�5�Ɗ��F�mSm�i��-J��h	b1�9������Sx�.�f�x6U(i�ғ< ��N�1ʾc�}�<ŚT�pCg��0J�Mח�=��A0 x0���;��,��PrO����p-�Z$*nWW���y�<Ɔh���Ve�8�4��X
xl���q�Ȳ� "��T;���zXy���ܿ��H½�W�34�dJ�Hm!y�8�=�o���Q	�f�+E��82T��j��"
��=؁�@ƂL���5Y��g���K+vZ�� v�O����=�K�`����t���Eb<Qc:)X���X�{ޝM�I0�'"�D�W� �HL������Z�+Gj�_A��'©�F��#�gsz��� �`[B���=)br���b�|��^�nk�]�O�X�}u䳎���P�^�"H%��P�`^���l����@�Ȱ9��=�y���?���o���x�)>a����w�ml�� �� b&``J�)��.�=��{�w@�E��h�fMW�YY�4�t��	���C�<n|���!�KN@�(� ��7΂�="¨��S�dl�1!bE�5����٧"������ )"�^D|�z�:�æK��6�Z�;񤷺3���|N�n�4�d���o~�D�u0*���|b:�<�ʒ�)��+j����J�`	� 1�������à�:�rhu�7��B���0��ފ)�Q��_��Q�!��"�����������P3> �Xr� u|��_�>���X���E���_��TR�/_�V˘ �$�{��d%���x?Ҥ� �|��� ڂ������|���皼�;!@�0�`��w����vC���{SC8�ܥ�2�¨�@!33W���C3� 0P^
�*�>5 �x��ܹ.)����o��g�=c:�����g���ȇݏ~|��#uڪ?P��˔DR���PZ4�2b/����-�m�`z�a�߸�t�!*;�2]�B����}��K�}��p_>����+w1x 8u" l��:��1�KxR�)�}��C~�U�/UG�=���� ���xh�y��^�O"A�"/��� ���k�UW]���PMT[���<p�ZFܬY�L.���,^����	u�U�;q�̙c�O��)����ɓ����a�\F�N^,|��./�(X���{���~� .��R����b21aTR�͛'絃#��-Q����Ȝa�+np �E$�ڜE)��2��x\��)İ=:� �� �/��U��I��@ ��cG��QXʄ/p�_M^�Cz�U���=�'��)7i�<���\PtS�1��|�,��#(�JpK�[�+���K4� � 
((�� ��@�~�[�j`�3{�[��<;�:PȦqM:�}��6`�o&�ːg 6y�>��;z�\y�<-l��j�b�\�QV�y���_kG?i	�����=$@�E��wKd�3ْ�47�y|�ˀ�e -W@��X �"9�+T�@@	P8e���W���u������Z��w�o�p�Q턬o��#�6?)X� #��a 1{�7���<�<#j ���ǥ�W�
F�L�B��d4���%�F�>�T�V�6}�s��@���G#�#]Cq�I	v��� "�w4��2�����׿6�>�ܪ�N_������7$1��h6i�dY�<����y�C���E�Т8�o,yB���A���P77�4�5Y_^�u��R��V�j��0X(�^r��3�$F�#崄&m0R#'�Bpۙ���NG@9��w��QP���b\���\Š�nYڰ#�+m?΢D{�Z֭qW\q�m� ��%Y\'�~�NF����h@�� -�bO)��	f��k�� ��9���(�ǈx���l��MF�I�4JJ�r30@U��@�5�C�7�U��s���ߡ�sT2~
	w��(�RM����L�4��f�mSE @M0Ê �`�P��8�?����7�k|�X �����J ���%�m $o�-G(9��������{�x�bs��q�y��,���~�ӟ�Ye�]�~J,3ԝ5 y��Wyi�J�U��
�#:Hؐ�J�e���_G����Sj�����&H��\A�?� ��ȗqd��!�e��@�
?�;T����F͗�� �8q�Qq�p����G�1!c�$b<��y�)wU�9�dNI���7h��j7t�[��1�-�}{�vw����.���::P�4X��؏��zP9�W�A�_����x*�M��۴|^)�Īd��吐�aR�^��BJ�������}9���\9�e� 0��Q9��v��x�8�u�򖷘��I'��6h�/��3��#Pl�Ǖĕ���	Py����;�^z������w���E���Or�i刉�&M0��>8��#7�%6��а+�	&��E3p��7�{D ���EF]hv�ڏ�09��K�s$~X�q?���<<n��`SPl���(J?V�6Y-,�daw��xPu�3hx�4����M�[B|���̮_ߢA�^JW�R��"����o���9��Ӄ�׃��d��z���H����ϖ"^ڮ4�X���0*)���zmF�n�'P��n v"�y�t���dܘF����N�����Κ5��	�2(ؕ������%�Okq�H㩧�rϯi�"u��ڨ��.�E^�<��r�)�u�}��ݯp���o��Zm��R��+/� '��R�4pٝ�+��r]]>&Ǵ#&�Jpo�V�O�Q�K$������\Tږ�ڂemW���=x�*�'ݑ�ι����^�׆/�M��dQ�}L�@Vi j����Vz���㮷+�>t���S�~�uw��"�3�p�v�����m0��e�0�`]�'�v���)�LJ�Ȭ��J0Lf��o*�ŒD�N��L�$)ݪ��8�]Y�d�;۶��0���ޠ(UL�~��9�sg�)½��p�2˨�Ă�%���;+`��B��x���ũ�K��&����������"�=������xu%-L��ȏ`���Ǐo���	�M|t��|� ����@�=��<�m�l���D��g�zxgW��:pO���FS/r�L�\('d���et:�ۀ * A�l�e=,�@��K��K��J��q�������e�N##����7�!��k\���ɛ���뤴-[����֚4�<���Nw�]w�^#�9����{��$#c��z��d��l��tv�[�h3Z}�~zqG��]�-�-K�5RNE��VI�c$�u��j��t�$�G�O����nE�fW��Nω�'ϡ���PIuȦs:����KX��caZQ����[����T�k_����"TT�LZ��s�����]w�Ҩ9���
l��j1�f���t%���:[�º���ڀY	�f*���/�"ۚ�4�s������ۋ���Q�͛�����������w^d� Q��. ����η�==�A*�A0)|����NV\rl�?0��@��ء��ץj���Z9�!-Ψ���eu�:x���f�2��4F�6	����D����?��ΙG�����@�Im�)b�$�����c~�F���D��=<��>���_�!Kl�$ئ�Uq���!�30��p�d yH�g|X�A�y���{��ܩ�u��`(����	�	��
�>����<�#��Y޴�o"�M�6����m�c���G|h�6�[Le�]��#�x�nxpcY�P^�[rv-j��6�["I� Y~K�""�ۨ�vu͉L��>��}�1ڃR��Ϝƫǡݺ#��搠Lw���5�����;44��^���y9���{��,��ig2#�Tݫ�j��(� ������wާM��6��?�cF��]9���MD���0�LŢU#���$Sq��)=�*��g�J�#GDƐTTŉ�b��v�MV�K��(g�>۝��[�]�����.[�����i�2�S`{����C�PZtLP�x���M(e�v+�;�=���7i�4��B�o��;��xagV^{ݺu�!��a�抂�1N�	�(�d�	�����E?��6w�7ۂ�����9e#UB��oA[�|]*�j�N���xD6Ŧ���N<1a��[��u��~�S*�� `����d�P���^�	���<+��E�<���lP��:�v�W�8���;��Gf+��W�O\��u�Yn��yn����c�u��DVi��U�쫁ǢW�M�x�I"|8�P�/�%1�C�Ć����L��zW��fiE��m�\i��|�N
���(w��<E��Ɂ*0�7����$��_��W����A�9��j��vj7�{�ᇛ�5���܁j���<x؆g�%��'�x����Ysܷ��-W%������� �o��-���ƫ��=[�9�����,1Pq��D��P}ṙ��8o�������u�܈�RG���e%�<a�ڶ�� ��v05�3�s`>����k��.�:��G��jɣ���'�x�]{�5bn5pV���.�HMM���Y N���I�y��2��<��3,�s˴-��C��"6�*�|-n�<Xi���8��*�f�2@p���1�侴K�i�%C�t@N_��F�#(�R�-y�h��W �ȕ ���9�4��z$� <+���v4��O��S�)'�͜���u����`��G�Zs�5� ����<��'+��bTP"�a��ꫯv|�!�5ig����@e�kN
V���J��d%�ā'Ѫ"j�?�!pbH�Sn�x�3b[�v4J���^G+��+)Z��I}D�<����N-����4�ۛ��f��Y\�yƙ����=��f���}��Da�lX
���HW��J��Gu�Q^�5�9�2���v���)�O�	��W��v��6v��d�<�/��^�,�a�FL����hR��u N4�Hź�������V��W%%Q�,����kT�6 �Tn�2�Y8r~#@`��z�9�8�(�;�\���w�{F�0u�]c�V�7�1�q����x�������w�_~����Ns�Y⹱��w�}L�kì�A�ƍkl	�ܤ��C :��UZ߅cK��3D�1��r��n�=/?�����QJ���'WN�X�BE��y���C���hz�+;��$��5����-�P�u�ofc˜3�<˵i�v�Drx��EÕW~��a����Xޠ�A�Ix�e��o��s�=��ħN���XHH���{6�J��dU���p�qΖ��ճ[�bMT�WR��f��^�u�Bk���.l�?*���ԇ��_�JW�uؠcz�:C�q��w��3�">��;�x3F8��%^�Y�R�&H3n��FY7�"��gFJ���/h \�^��W�Q	��Γ�p�6c ���R���g?��QO�)3;�������L�H4VҰ��P�}�`C��ŋG�٣��'�ږf�̍ʻd��L��Udق���E@F/C=��%�@�˲�߼������|���w ��&
�����E�v�Ĺ�R��㠫MhsG�'�X�5ԍuw�u���W�po��7��u���Z�x�gW>o3I��(�m7�%�ں��xB�`�s��|��L���z�r���_�E�#5�4���-#�x2'&�ɘt�����a��w�n{��A�*����΁B� ��� '.l���z�灳}.�Bг1�]��l�d�yg{�(��� �/���'L�5O�΀op7�p���n�r̙;�]t�E��s�������u�v�$۲f�x�:�ր^��(#�0ȏ@���2����l�U�Tã���������Bp�ism6VG#%����~��%�\:<#�a���W�� V� ����>QO�shp0H�o٪���J���?c�N;�Ĕ���Ci�0����f\�����=���n�����`N6�o�$&}n}�����g\�FR��2��'aP�'n(๽��zl�ʈxH�ע�T,ǤӞ��)h,�\�Ī:"��Jp�ߝ�����RI6�t<����7T �lap A� |�J�X    IDAT �/}�E'*<�j��=)�W(:���\���fhx�4��[��^{.p˞~Z��:���%��K�R��W �.�T�^����?������(0�G�K]mM���V~"�=e'��C��pWWWe�\H�k0ީr$�.E�Z���0*��hM��3#=�m�<�έ:�`S���7�̀�ā�#��ꐤ��z�H�Հ�+^NԳ��^[��A�⮮ќ����	���wP}0-TEȉ�K�ɀι;�h
�� Z@�����m
E��n�f
U�����m�P>��ͯ8N2m�SbK��k��:��}��k�L�+j�s��;*���m�O(����JP��g Sw�uD��,9r��[l}�]W�t2����>W|r�d��i&������Q�-
���#}@K�Ȫ`�Ƣ��SNr���g�#߶�E:.���Rռ��K���X��6Uq Ȥ̼B �ؗ*�Q�蠺c\�)�e#K�W�����,�4�^��
   �^��%�Q]Se�.`d L���}r�v��߶�X�#�C?��9vO�����e��R[�C�D���G^�>��=���s>��&�����%`w�w)mY���� O�:ո��$�e�-Ly[��5�$�_T^�JD�P�H�":f���F|d�Q	�������6)^!���PR� �
`r��*,2m�Љ��Vt{�O����
d?D*�F�Y��@O�֘� j�}[�=K	�d��mh�f���w��5E�{{���~v�]�*�(=R��.��7���}�B��a}!㉼�#����#bxa\G%�{z&�Jݫ�>�{D�j�
*ᯁ���5K	8�?���G�O����x�ݴxh�1t�C�O��7*�����d��b]�.��꼤8�d�_����ϓ�b�5߹�=�j� ��X\�/WJ�-�0*�I�0",��"~�"wm�5�lQ�[�dA��m���(G;Ӊ�u���}�T�o��v(�R�P�p`9�~� *�(|�:E�a{[ �k��n��y�,�p�H�{����j�|挙���	b/Z��&���m؊���\}B�B��p���p�������D	x��x���|��|B�,!�Q=�aB�5�X��∣ޣpA�"=�MD�R�X!&�-E��|�H��NQ�:p	��[�n�֢��f���p|�BXW�~�Zyb�W�d�;O
O3f4�$�o���U^F`dA*��z˛�e��#�&Y����6�p� �f�� ����)/��<5�`--�k��-+�m�����@���h�>emK��bI#�n�b<k��#��\���Wv�0
�]WΥDBc�y���$l�- 0@���?��Sm ��T�������1�EC��矅$O��8�v�-[ni� ��/`��-�k�j**�Gy��K��a�`��=��?,���~�Iw�]w��+N:�t��ծ�u���M���zK�هن4�5�����Ŵ�#ENX@�DҒr$�b���ҕ]ݣ�Kd��G�X|ugGgj	�� ,�l DA�)�HV��
���>c��'���������vy>�� Jb:���(�?	�CI�?雯o�������ڵ����vBZB3˥_��ť��o��M��\x�%��/\�A5Fik!��a`�IT�Z�q�0X����$�B��T90��{�0B���NTNVf���>��PQe� P�+!HF  2n���=V�
h�����i�l�/7MM����x���S�E&�,,�5H�ee�9���PU!�Hl�ڵkm�g@b�U+WH��j�Y���!^��l0�����M�J�����BiC�	<��i��{<�'$��+�r<�!���t��0*�].W����
���`���H ����
O�>7� �W[#����Ǐ�`��p�;��8��)�`Q3V������ g�˳ �h����cB7E����N�'�|ܽ�q�ۦ�(OR�,o`�pȃyT�AI��N �a��@ⷼ^u�;�P^�dI����6��=ɷQD�I�SH=T:�Ѐ� � �~�1`Y����D���^w��6e�[�f�tLnv���&��B���vx��`@v��C8w� ������9*��:���w����̠�XD���y��?ވ��	�)+�����������%�Ή
Ҙ�೬�93����	��r밺��i�bNC���R��xa|{���7c�$���Iz��9�Z\WG����ϚYF	_��W�;O}�9��?�,�$B���\^��;�z�������C�VEnDO��I>>k��֥H�X�-���5JLR�Vq���W)�qQ�I	�A�`����w3�f6"����LjG*��D^*�LJ��u�{ڴ���֧�W�Q(t�;���HI��~��3�k'ˁ�M7�d�ϐK��+_��[�j�m�j�'�S���抁S�8<�c���X�����Ͽ�����c�<�#��VF�LZܣ��7l����!����q�/.��u�Yc������5aԁ;��Z(�38�7F�5⇽~���NlE�:�~��6/j�V �wJ[�Ȥ��Dj�6�� ؂��OMZ�nI�PxB�;��ʎ)]�]��>V'������Z�v�`�}� x���� c� �0H������d�5�M�T���rz�܈�Ĉ�H �K]L[0����1��oѱ��eB��O�^� 8��$ ����d�	���X�[�#�wJ:��GG<�@�B�|�_�e�=���҇gl���I�SO-s��|�r�����WK|�x(JawI��@�\ ^�8~0���&�^��������.��bm�0�G�lD�V��;"P���,��5]��9\tq^,Q54�B����0��zV�<Z_�M��X�3�M&-9�E�/}�2R@>i�d�+��pw�_0�w�j�������;L�5�HR���R�ɓ��N'�9��a��PZ_�hZ�����˟��[����U� = �+�D���*hs>���W3e��R_]}�vF����Ė/_.n�(��v*tDr+n��	���v�g����S�W�F'�Ǝ�wR����y�m)��,������2�3�=��$b59���O/�0<<_u�{z��ģԛ�r��Xr�d2�)[� �$����P�ԒE\WW�{����<q�D㛡� �<�Pf�#�8��}�<� P������X�2��T��n�͞1h(#�D�-�}��J���#Ik��Kdzr�����R>Z[;��;[մ������n�xi�-X�t!� �S����K�5p���/��%��д�iӦUikmm���j���:M��������;���H}~���'F��I��hYs}1��b��Fr��&[j΢�1�.h�!Y(E�3��HT��ڷ%J�h��ݚ�d��մ;�ر}��Ha�<`6�S����렣�u�ف���G:�mj'�@��g �k�q�s�"Ӡ�o �I( �Xe�����^:"8�� .��	����4Pa,�E9�/$ZdJc�|�0��ߋ�x�K���.�ރ-	&�s.����	0/XZ�+�����-ֵ�u,�0cƪ��{L�Z*56��*�&L㸆��]9�ɕF�b,���)�E92k�>:�-�(F��h)Z,um��j!6_��do)2�M工]��N������L��4���6�reK����Q��K��������6�4�Iɪ�"��I�a�H�8�*)X.�uu�|Ok�:^��R�ڀ蕓�Bv SǙ.�BNjrZ�E�E�S�G2����ܪζ���J�\���6։���H����	�C����/O 0 pf(F�� ����I��28|��OVD�H. ,:( 0�R���-Gq��2Q��T}܄q2W�Ii%���Y�:yse���%�	�b�.y00��.�s��M�ԋ:�qݫiH�^�d�ɾ��f�ŞX"9X��z'�tQ���II��"A1���"b�
b��IR��~����b��:]9����<����3��L��*_̯�<����n���C��j�ͷ�?�����/�u���x������T$�O_w�Q�xdL��;�l\?`�%۵V:�¢���v��&W}���޾�v��<�eiF([H൰�&�^��b�!�l?ƻ6`֬��^���
c%,@a�����H�:Ǜ�������5#�[����*�:�ԩS�NUQ<�2���f�8@=tY�G�ճ{6�@2X�fx!�3&K��1 ��wٝ�^9�L,ɨ,Ϙ��y���`Io��r�<��\���j0�i�l%�A�,��d�Rn�����~�G�׽������%=V��l�rC��(e����?x0s�ո���W2����5�!������O��W�n�<�Kc^�W��ԳJ�����ҧ�N���{�{gwe}ue���{�ޓ�޹ra�����k�o��{���ǟ���o{�;~$�~L�����>�03������W�f�F^�v��3�7�����Np0�D�Yx�T�B4��R���	�m�S�N�2�A�uu c�g:S�;�B!�⊩�ػKj/m�݃��	�k�W����a ɿ�7�F6�����S�xO�L\�O׶��]_����.K���ͧ��{�~������o��L��#a��sr���A��{��*����Gԉ���Gg�����EX L�YyF,�����ԭr�����l|�<��U�C��O��4rG|7��Çv33|aucm�����pbym�On���>�zv����?x��Gn��ޓ�W&������<���x+S�^�g~���W>g�Z�gs������qi����s)z7�{�H�Ă�xn6�n�,�c(̍��`!d�"���U�3��/��o��L�
D��`ZK�)&3����~��"!w�E���΍	�$���������ۓF������w��\V=��X]XW�g=�Y�O��O���7}�7��Q�q�1L���!�<]�gTou.���ׯ�i���3�z�6�h1�����i�>����s�v���<G�-�w��jYc�{n]4�����3S�ֶ7ߟ�y��������Cǟ��C�����2���DV��Hq�K�No}Fv�y���Sw�̎��DR/L7�/��D�/&��:�b6�~�U+�a����ǃ��Pq���O�;�R��.�e��N�C��75૿���Lw<'��*���E��QgP��7|�7����������g6�	P�g�:D]�jF��Hy�t�������������u��G�o��p���aR��]���7u#:r��5|���:�bp�ŬE�z������mu��0F�)G\|M�e51�g��m����3���o[�3/�랻���ͷg�^�s=>��=�O����������/���z��>|`!��r����;T� I��w��t)��#&��Or!;H��Lg���dt�٬��q8B�D�`Vя�2IKj#:�C0&�lW�"U�T�N��O[�BMZ��ݭ`g�+}7n�t_�z��{�Sy��]�Ƥ�Ν���7���_[�8R��US�����V�!�j�`"���o��᫾�k
�����L�	��7�����8Ĝ����gŽ�/���d��w;a����dZR��x��eSc����kX>������=��c,��e-�L< �����SK�/�˶O��?~��#7���>�߹}��F:�� �@����0w�7�n�����寞���ԕ�g����9�ըU��K�d��[���b<�q7��}�6E�q�+B�Q]�i��t�ē��(�܉�Ӌ�P%�:��]Ҏ��n��<Iu���OD������|�v[�k�s��w4.��g�X�q_6������B4㊇Y<;Ռ�ˑ#7�����,�J�.���շHkV�ƭ����+����о�M�p��O޹��ңw`R'��r��ā���3^��hc�ӧ��?���x���?�1��dm���ý�ؿ�����{M�bn��N��~ڥ3g��?w!���# �6KZ"*�
�ƶ���9�T�B��;K���A>� �"C@�w^��S���b�j��Dhy�fR��H��oٮ�7$GD���,��Q��vT&:��$�W��e�{ߜu��$Tҧ�t/2J�q��+��j�H���F�ǳ�ál�Y�@}T�������c�>�|1qMjh�)w%�U�:13���w�޳z��X�g#S6��L�*�[�7��� �w��מ��~�OT�Ld��"����h��d3�&��˱)b�Q��r|]R畩;����/�����S���O�m�|��<<�������0|��ӟ~iz���o�\������?�cͨ@G$yf-�q�K�Z��C�|�h�?�ư���/)�FD��|$�W����V��C��nx�w�S*�0��`�%_�(ґ�&W��]�ӧ��x ��ߪ�ģ���W~�`��>��������8����2��˦��F-�����|���k��kU���\0�9��J"+�[�n'�QSTM����u��W�2��O����4�������)=]�[�}��* 
p�^ރwf��OV��fvh�!�ď}qgys�O�f���>r��ҍ|8HO��c&�����|��.�^�ҍ��ϟ�\�5{I�ؿc+��h� ��JAߐY�a6��pQ��Z��$�3d��^$��3�l$'d��J��T�+m{���f:3�i��]HL�Uy����^>�'RK�����NĢ=��|6�l�c+G��XC~$֍/��/�e���%/��bd̪�$���U񅬆��c
| 5����V�=)WL�Fz��ɜ�v2:h, {&�1f�\Iaeß���uBS��ta�\��q�L��oA�ɿޥ�9ݪ��$���v�2Ѻ늩{��U����҇u��/-uI��u��v!+��8p��FއƛQ�&Z��X�,������}��Ɇ��0�ߖ���r��G�6�"�E>���W<e���?�Z9��O�8�"ڎ�{
Ѻsā���QK� ���B :e�뾈�u���� <��ż�!����K����K��Y@���C�I�Kc���7��~����S�F�	$=��bz'���!P�Yx@/�c�����L�R�^����^�����ۅ����۠W���V�^�՞�U�JH���R�s�+ߙ��{x��-��<]��&$���|U��$Iǳ�z�Y�2F*���#�mrh~~vcb~�������ڔ�UE~������b~ߞ��W~����^[�x㩓��`�XWX�T	����V���vk*��׆ i��k��0o���֦�+$�N�����e�\za!oļ�������W�z�^�`
֒^7k%�C�>��R!��7d�8Y_X4�k�8����eԱSgN� �0�`
S�/=7�I��߈��p滼{��꩗LГ���;�*�w~p-��4*��+8���iq����^~%�o�kKs�z^&�X�b�Z?t뭟~�����>z�����w�N�ϋ��|��֗ޱt`�;Ο~��# r �Iӆ0�O5
y�!�*�\�#H,�.�p���+�t�.�K��8�}��l.�Yߣ�\!T�����o�3�]��|]����l��ggx�6�w!���<Lа�aYN�n)��m̷���K7M:�.�TnjU��G�H<�G���ޘ�6^ة��V�����D��+������*�phR�������N���Rz�v[���S�J�P���/�6?{h�����QM�|̘��g<�kN����;!�� j@7�QsU,̑z�@��~D�o��W$J���Wi�����Y���&/i��iDH^tu����C^D�W��ؤ�P��nԈ�&eC���1Q�9�}+u�٪�F�b��=��R�t�+9�4J��w��#7d�Υ��rąem�\T���.:�1&{cd�jvz�'0Ի��`���װG�
�����z�c�!���T&5�Z�v����aΡ���A��[��QgzV��qYp�!/�S�
F9$��_$/g�onj�ݙ�[��6~>ƈQ��œ��1��g�����y蹵}A��Pk���P�{�p��|�
���uDt��Q���
����M�;�i Z�(    IDAT�A���z��Ȇ�$����J|���r��<��~�JJ���w��T����ʵ"G�����5n�6ÉI�:�ݷ���:^֕G�Q�]�����R���|�����/�o���U�����p��{5sv:��a��Io�y���v�1�hf\�^��鹩����55�I�'�$�>&�}��Ϻs��cߟ���ni�R�9��u��{e�G��8.i�M��ّ[�tŝq��i���l+MbW���k��"�����Q��J�Ew���mq\%F4qH��0��6�D|R��b�����+8��//s������e1_``*4Ѕ��8T��Wӝ��$t<�����_%���dV�[ƣk���ge�O�j\���GȢ�<-��~י|���~2UT���V�-d���&p�A\i�+[����ixe?5�rg{cnwfϹac���6e��D�����G�.^~S/�q~�;��f%{�	T�.	 ����p��&qB@i;"E���tfw�w?�;�����g/��?]�5¶�:L�)�Y+�����K��tkR��NiH�Z�������pI���]:eˣױ�������4B7��o���o���=2K��ǵa/��_�>�wX�������Ckߥ'0�(��峇8A�<�t-�>_��>z���{����?�l��E7�U7�RKn�F� �WƳ�{'N}+a�/[%1is�W������S�x^9N<�z���x�ίK�e�.ť�^7N�ҜU��!�t/I��Ҁ�RU�Ґ���t�M3��}��W�u��O���)#ϥς�b��!ӣ|{�������M`(sq��.��ΕOz��oD7������������|T�2UL�|`wSz�C��D��HeB�D����j�=��"�dƲ��#�%W�������/6V_nj]�p�h<K�5D^y'����<��Gs߉wm^��o����w��w�(N'��n����0��4=�o���u���¤������?~�������p~�`l�Wur�)ӕO����^�t��`�^���^�w�o��;�V'sgcF�{��\Z�A]����=C93;w����ot���uC�EܦZt�_AT��`�IZ-4X�v="��b녺e�~ @>���y׃wtY��`!]�|U�k'-�밺�!��i����Ο^��ʾx`xA��_@�_+�ʧ��I�OX����
BX������y9�<��奣��������o~�!q�K���в;����g�l)+���`+��J�ȧD�6s���~ol!n�t���Jp���粠U�������&�o@���7�ẙ;@lB�[ٚ`:�P ���u�"W(/n�<C|W�C>���G._z:��8�*XZYWผ�In��iy��c�������~�
~k
�Tp���T���_O���
�t؞(�eX�m��v��zW̗:=02�:�ۜ������I��No�@>�D+�.Nm�f��I���J}�1^�N\�����a}{����ŻS�Gt�^��j�[��|Tq�_˲�n8��xTP�F����Ō�B]�.V
�#f��t���g�]�B����ECZ�m���&I+�|��fr/���t�K�$��;���D�~$E�)kE���X�Ȋ��F ��2���K�$��a����^a�n�zW)1�7����a*o���O�ޣeyU�'��U�x����l�ٟ���m��2�e[�c'ZG~�3��~�r�ک�d�R[a0���][w
[�5llm!-�OV�e�#u�"�ɐ�s�{�O�$�u��qM�^��	]���Y����[m���3�8rլ#\����R��!@Iki�$�������/smp4�,Ď��oq��v�{�2�n���'ʣ�8�(#�5䤪t�6�+y���z��(���0����c#f�7y����i�{a�\��Bُd����'}�'�5�B$�ox���t�-�Ui�~{(��])[�w
���#���Rv���+��
�v����K��ܸ�a8������2���yt��<�,�+�?ȮB\1�HH�BР�������X�;QZ-���1+n>U�ѻ˙]s#N+3�b��E�� ��	-�����S����*n"y�ǳ��ӞG�I:娑 ������>W\>���c�	���*��Cj7f��
��Ԅ���ٟ7<�YώE&[��-��ٟ�%�4�C��U����?��/�Ҕ35|K\~9����邋N-�_�|HyW��\b���'S�痟��/�;��=����u���{� �<Q��^AxG���W$w#gϧ"��H�C/�?c"i�u���L�zz�����ǻg�����Ov��Fx�l*��\O�g��`e�k�ӌ��^�h��HZ�z�)�;��ӑI�<�7&=�0����o�NX_U4r8,;���re|����Oy�𲗼�xA>�eU!��tT_&o��{�bh�ǭ����w�v��<=w�0\"���$x���ލ������ B���s�v��Y��X�߉Ț&�tˍ�*���@�˱�D-;������t����F����� �'`R3��-Sl-JqE�*�Z�^�	2'R�PD�UR�Ce�Q�'{w1F�[�3�[g"׺/"��K�[A�).���u�[?�{�<�7��I�G��+��`+�_;�/��78��-~�"e[)c�n�")W�B��tɊ(�O>�;}����9ab-�3o�M����l5��j�疲�KV-e3���f�c�����d��ȅ=sSi�ᡝll������le]ힽ{v7&��H�'���q�φ [(�iE�0g&�;1��A����K6Y>ݭ��� ���p[��(����G��2���B���9'q�tյ��*�����yYjP)^��W���z�Ԧ���=���ɫ�W�8N�(]�Mcz����p���匿c�06�%��Y>�/��R��v����<o�b5��:���UY>��ʋ鱗+�1�U�����O(�I0+Z�VC`���?���w�}�����~�44�Hh��� 9N���K�-Z`�Q���C��U�{��W�5^N/�U=�8��"��s���|#���Kc���c7.�\�ɵ���/M����h�ַ�0���n�_�ɷ4��HW�IFI�]kWhЭR�5(X9`Q	U_i����#yE�,���(�3�����7����YN�83<���*Y�iVa7e�����q��;�=}�r/n�ά��	:�$�9����VM秪�F'T�2��y��?�j�ܽs��/�Zd�W�(� DjAL��;"X�ᣡ8�	�[�b��#0I�Gtj�@��������h%y	wm��������-��w��{��(mO��G�}�KO��Elq�o��iz���޳{ﮪ�(^�#RB��2{��3ّĘ�ۦ1�{3ҙ
��=V^����7�B����+��A�͑���޷��C����A�dJ��S�;���z����<t�(��v�&����uI�ai����LC�4��q�w��_u��qF FB�[ġs6_UJ|�5$f���(u]��nZWN	��o�����<�7I��z~y7�OF�p�W\���@Z6�|�1].�*1�/߄V7���Q.�6�V�eN�kJ��N__|m�h�ԓl��M�,���T�����zD*�z��g���������uE+��.���C4 [6鞼�?���[�!��2f�xs�������`0桊�-���8F��Ȏ�Y�=�?\}�	����
Na����r�� �E��Pg��w��7D��->?�&���ɧ�����z�^;�H�N��siE�_;�^uj�V��}1��}�?�P��5p����\�~8�zZq�{?y�|����ԇ����gy�����?���W�Doy4�vOj�te���ј�ѫ�Ԫ�ұ�����]��d9{S�{����I|���|�<.� ��[٣7E��Å���_���t��U��b^LӃ�l���k#��smU���z�'U��J�w��ܒ_&�Uy����d�sT���֍w$���t�t��x��2���7��Ǔ֯O�hT�e����W��wqFگ"]�/8���Xޏ�<��n}�Ϋ�/t����H$��$梃S;��7�r�����=ç��u��z��p�Y+�y�_���Ut���7?R;���B?�<����x��Zp��=�,i��!a"[q�15�5mj":C�$ ?a�Ȭ��I�^�2lڢ�v�t3]$� �*䏈�s��ǉ�5Jk�pa�+�������?ګ�������0~�߹��������޵?K/�x�=���ӈK��W^��}�Ucz�^�g��w�{�����y���w��S[���{�N�<�#��;L�����d��w�o+5&��7�0��>�t���I�Vf/ϵ���a�����'�V��������LF��%��޾�{��+i=Lv���H���uN+s(@�y��ԯ���AcBH�Ii������xR1��+�Qِ��	ʰ� N@�N�'Mu��ֶ;"/K�Ә�f�6���Z���	����R�*[�|���;q��
�U(�Ӌ+�n�F5������|*⺧�A �ŗǇx��b�.��=XG�;�f�>�t����/�����o��on�	;�]#�-��l��W>�S��G��*{��h�����@V'͆�eUJ��V^���~���[��o�R��~fI�5�-r����u1�����`۾�� �s��*P���>�|V�v�g��p��ϛrE(��z���ؒK��8�����`k3�b�c����d���Gq�OB�LCh�{:�́���K��^���myW�����\]>Bj���z��Cބ���j��J?V����B�{�O�1���W:��!.�VY�)sq�ۛ�����~�R�߯z��>�/����}�p�����~�6���~ș8Q˶��%�jS3�'��Өغ�2<���,ip�Sӳ�Lޝ�3���Ԥ�n����m�H2"r.�B��m+8r�8�I���"�c����b�D�-�c �{���þKmr!��!H�=G��<�G'�&����-�M>�#��廸���I�&)�=y������ڽ�͓�����j�����_�Yp��P�	L Ʋ����Vޣ��>�t�}�~��|\͕�ا�έ�ɉ8�|�K_:|Ƨ~��-����=<��o�v��_���ĩ�ɣ�䟊��9`�p8=��,0]�eñ���{���OfӚ��L�'
���'�>���3�eH��T�%t�}/���uƤN ���J*cdӿ����B���!��$4�F-�1��oN�9yY�W��?O�D�
�+X{�L�b&�UNoT�`y����������)�P�?J�����.�����O��Qo&8�@�D#_���UP}m:<}H�K��;ʂWe��.������k������A��S�����=ï��~��>�6�ptq�[�e'��ճӣ�������&��ԫ�0 K�o����(���h�_��.�^^>2�8s�� ���( �����}��	ө�|�y�
\Y^�s?��>�ޓb9@(V���oz��7�u��}�~���=o�ɟ��:�#,.�+��ʸ6�r��v�Gjh�z՗�hl����;�����lͭ����֒��	��E䗷)��1��Y_Á)��P��z�����^��ڜ�.��?tl����:#k|o~���[��IɰC�i�(<ZA���v&z�s����$2&FGA#��3��չ����z��/��jHg�س1���_�_;�c7
�������{���a*k)S䰖<���`l��q�F%�]㣚���S6b���'h��N��ر#�w?�  H�!oT��Ґ��g�7�rg݀mo����l~%vR�:G�����[*	؀�U�9s�B��;|�w|{�Nk���?�#����	���ј���{�a��ī�+��+r<�E`�����J��^�A>���J���l�:��-��]��L��ٟ��÷��簊?�?0��/����_���b����3_��_>�������2%��0�������3)-����*}7pe�y�q(=���՜t�/����������-�Z"~���_��_���0Ҝ*��8T�ip5H��aS�{ev!���q!0������1���ܟ(\��a�;)�rP8`��X@b{�:�L-���Ib._��_��E��d$�{2�0x���}��8>�s��q�)i��HC�k%�r�,�G��޵o޷oms����^���d�_�_P�Ol�Ԇ�V�W�o�=��՗���>)�`r�]���O��=�)���\��;���%a�����;���m��.���ۯ��a����ׇ���/̱#�~�~��%Y��K��8T�B}�O�upO
��Fk�|3=�י��gsϥXC��l���a��g�<8�����m��c1���b5Qi�/���S�����-��nY�S驯�b_�3�ʋ�ȝܰ���G>�3�m.޼���� Pq'�K+@���y>[��ǜǬ�mo{[I�8����˾,��;r��㱶L�|�wf�ǿ�3dXItϘ���.�3�z]A`�
9�k���B���g��q��|���~�T$;��E9�:�����g���\}���r�9�I�w��g�D�x��v��������C�E �x�;�#Y��ַ�%R}e������P��?"�_���}o�+Fcʿ�Q����v~A��u_-�����w���Y�n�������E�F��,g�:9�J�O<�p��7���Anػ�+���iП}cL �&��}�}oM�ϼz���7g	[�2"����?�����?�;<���°�BL����W�{@�Kna�U�+�>����4����>�6��ew�ts�4�o��?���I�?���5$�+~���3�п����YHW#�82�V�Y��&Tp ����XjFk�d=�Cf:i���Dv��xu�ո�y���Y7�gk�����#Q��ﾲ˷�H��h���3U�m��#=���O�VNb6��ȍ�2	b"d5�|=�g� ��I\sX�c9~��>0��������^�ۤ��^�d\�V�)����k���M{΁����Hە���4��Q/Wt��������<�T�O��ό��[�\j�C�X;������7���R��TK�Z���.��M�W�I #^�f!��ɩf`m� �r�>M-�IO,%�'�yjT���_��+�W����K0��6Z��A%��ظ��a�GI�d\H��*��_(�6�7���&6���w����_ĕ��ѸH��Bڨ����׿\5��J��,?ݾ2�{�Ǫ�>}�'>88�@5p�^V�zW������o=����ܻ
tp���A^��J6ݜK����|G�Ͼ��/��M�U��n��v��ʍ��F�ꃦ�VWe;5�۾�j=�|������f)o:rc�{Q���~���9��Ï�~�A�B��W���~���6r��Ɋ�$�.�I"=�������3��;�DǛ/(2:@4���>$Q2�,W��BN��� 9J<ibU�D>���v"Q>4<�O�@�͒=/Ӿ�rP�#a4�=�z�S���aLi���eԔ.�FnJ\�����[܂��`^�o�G���nd��/����_4���Q�W^Ș1��).�	�|V�c�gd+|@@���o��OPʋn]jNf�o�*������/���w��� ���k}��~�Wf&pf��_~Mj��z�R���
�wW�m�{Ե������
���c�Y>�s>o�_��Ұ��ON��3ܐ&��<���{�뻇;��$q^����4|��}M�ٟ���͎\�p���1� W�Oj�?��)\�sOM�9���r:�v��ԃ�x �k�u1���R�[�,q�}(=7 u��W��v�l�a��� KE&#-x���^R2���l�^��/zQ��㮝��Ï>�ٯ����1��e/)"p��������%��}5�Q��'C��i���=WL��c�����%1������J{��r��w���QJ�!����=�V��_��Q���    IDAT��n����+τE������ַ�e��O���<��#�Z�VQV?��O{Z��Ǉ��h���=�%��ww�R�w�F��O�Hh����j��v&����e�K�6��~��_��_�l��^=V�;I���oƔ/]�bXLj���P4��zFǏ4&ox$l���o�Lͦ��i��̮K-�0��r72?��|��g�����)M��*�Uӯ���Ga9�2{���
�Dc#G��w�n�P�|K0�I�\�<z�C�4"HZX̠o���n�0��$��BL�4%+����_ؽ~y�K���I&?g]�G�!y#�������� ,@ӿ�Ù�n�����Տ�*����dS�R�)��kȮ�<x
]��wy@X����g�}�;��[�7�H�����|ӑ�[n����� ��F�������B���58e���3�4h�0Q`h�a%0�&ϟ�@���kH��	�ӳ����������wxg�"t���i9é�xb.6�c����o	i�S㔎O`�(���[�ի,_��y���z8��1������ǎ�i��/.�wI���%v	٪� �Zu���c\���m���5*�;f�����
�Or�߈�@Lg��wI1�wo�C�u�a�~_0���gc�f]�?���CA��p!'<��廢,?>�$���<Z�1�ܫ�?���V��	�������W?�_�x���w�u4=ȥa#B���MpX�63�6i~����п�|!��j�,K��6�z�k��_�Aazk�&�^�������� �ıJ/F׆K�DW�xG��l�܋#(��zF��3�$5pV��|{��\s��ݙ�����(�!�I%�
��ݥ��{3=�ƞIdȃ�MDZ����$����gϓ`��ݩ0�ެ��Z�r�ﻟ��&r �#���LcVVkdm��۠���t�X!�8��m����{-�*ǩ��6b����[���x�x�.~T�b:����H�{ۼ=ߚ�.i6�A43�:a���������O��텃��c�|��7Ǔ���G�j��kJ�+�yO5�o�U���i��L�����>b��9ٍg�k^�K�'dy�������H5(0��� [����(匟sΧa4o��l����IŏB�Uc��O0eNN��(X��ӱ�go�ƶ5���듄���|�ȯ��dN#LcQ`�ӽ�]G�g��C�F���I �2C!�OB�=�:9$� ݴ�]��U{�a�K��A5/�2��_���3�,^�^Z$�j1e��^8�'V��4����P0X����\��-�{���v�v�mW'Gj8���=�B��oP�"(�4�*�Ӆ�Ue��Ry+��wo4�3k��yz^m1Yv�������a��/��r��+�\]<w��P����ϖ�O>�\'�6�ԊW8����N���A819��ẘ���ޭ�L~��v$�AGH� ��R�0F�f�1k��vk�Al���a�و`�ࣙ0�v�M��t����2X���ЧcT^#r�F��b�eOhAtG-���J3B2����Ԣ��at'�Y�D�Y>;�n�r���j6���9R�zT��p1ug;/�>_�m�U���I���xR��Y'�k�Pꍾ�#��<�0k<�K7��TX�@���icN��վ�[Z��<&g�ங �0<p5�쵿�_+�_~�_�A��	g�c������έ<=�\��g�Q*'|�� ~��Ō�0 �M��Z���a��y����#�6��O�����D�k�P�0ĐĐ��v�&���d�1�JBZ뮚����#�H)��FD�+���a�^�RMO�>dq�ԨEy����Y뗆���̬�����c�vG]��O�!Y��zzj��"����A��N��/�y�H�yO��t*�qL(a�����x���𑴘�`� ��#�yYL�Ӡ�.x�Ȯ�c���0��?u2L�E������ޙ�	������	�ݎ/Я��o��M���]Ϥ�r��0�Rz@y1���2�3����'�����mI��4PyD�f�Y��[�0Uë�\/s�����V��R �}T�=qi���:~�x!q&-�ַ�đL�$�_J�O��v�g�T��q�Xf�G�ϓ��j0�/	����g�K��0�l'`���{C�W�1�&�WVNֽ�9�Ue*�85&�4ճ$�Z�Rm�qb�|���V�_Q	��`���J����d���f7L ~����}����`�)��1��W�8a�8aϬn�\��ܘټA5�0#��;����lcv�C�P�E]�7e}$�F����z�a �F��H5>��b�:w�lᔰ��	�C�r͘�"��N���p���Kq�:Xyj �"�`�Z0��PL¢g����e�F$�n.̡�ui� h��fU���~v�������r����R'}h���r���v+]�pVSS�1WL99�f����AV@��L�t ���c<�Y\j��z��c��`�����5k
�|k8�BzoԞ��BL�9�0;��j��Y��1&k�ڪ���Az��O;))��.D�.=8���2��`����$(ݐ	��;��&{ab�$�3��BL��w����1IO�b\j���ķd'�����N�lG�۹��!�.�A��Ԑ�2�_T8�j1@��աzb[Dx9
�}SW?,����2w�ڞb�Sz��J���tS<ƴ��k����R�t�1Q6�2��z�jĭ�fT�d[��Șj�b��"Q.��Y�:������� ���ވY�Y���F1��ҿ��b���gWwe#6SJ�cV��-d�ާ3y����%�4��[i�lX�өMD�xQ�lS�<gZ����)��E@I��*����	�>�`Mo��*wz衪�S����g>�`�������^����/|�pv�����ǆ����j��;�R���A������.��}�{����>��k��b綀��WN�>QL�LkSL����=�����}[	*s'N>V����%�1<P�r��0��l7�l��o�3�.ޓ��e&�U�H����B���>�qS&N�<=����(�����a)���n
��I)]lx%z��X�F��'Y�]]=Y�l��t���H��O���*��Zx,���3��G�v��
o������i1�q!2���EV��S�ɳo�!ܖ6 �VF�.����$kҊs�B���F���	*�S��S��J���|�5�:�8����>��컟�n�3Ir!|S��^�Χ�5�-.7%_�tV"�����|�wg����yN�>�y睵��ƛ�S#�Ǘ��*�iO{F���;�|h8P�W8o��o��z�~�^l��mӱ5&�:V���?����w?�h��OzY���0�t䆚�����\p�n8�	y����^�&��Kʅ��~)0���C~��ǆ��W�Z�3?��´��i�ǆ;�s8u�԰�/� 1�Y��-�^mƒnM2c`L�`����U1��g�v����dH�9I��$��K_2�쥟8�IV������m�҅��h�!`N����gO�4�7�J����|�/��Sgn��yW'��`
���c2�M�O9]*H/���2����.u��}D����Y\��AI
?���q#L���X]��5asۭwd��=��T���bq���RU�?�̙S��q;��p+�"�9w���$�:i���f2O��PT+xbb����n���9|�wwԧ#Uz7zV�O�M@���I��#s��2�����
ZB b#�"����b�����~��|8��L�F�=�����с�y�~�
?���E|:"�4���0�3�۲�s�*�y�`{�b�0	��g�df<KQi0���^[?Q:���_;<��G�,M��A�����
�r�b>3��L'�_L�B �:73_y{��j��ܳ`·���Uo��M��̴"��7�T������9�	s^H=��L�K�������?y���[���Yׯ!�z뭥_����5�u�u�Z5e�e�|��B��p�L5���� q�\[�0�5�'3�R_*����U��\z�'N��i�c�@���p��7�a��8Y���M�&&2�N~��O�˗	����Gؔ�z�{j���}u�C
&!I� I�id�� h3�����vt��<���ܘD���F��d�0dC`�+�8yr;�a��(}/�l��
.Fb�o�Yg����K�=�k`��w?>�|��B�z����s�f(��ԏT�ٳg�T
s�O���~�=��c�d0����Ԭ���յ0��Rl�Yf�05�y��ß��ñ>Tyr�GT���OD�&�KÝ�5[H�������^u�!%�L"Tc��v2,��m���a��c�c,�y�*377�0<����>������|K��&��L�W�w��a��2��c��58 3:����ܡ���L$��f,2Q7W�Ŭ���O��O6S�0��Ӳ˙�<�S��f����_��V��=q�^�����B����Ioq�'b��$��*L��Ku�Z�g�DT�)]1�kS=�L/�"�B�1&U�1'!쾬�DdV L�����՘�$x�Ɋ ����������X����E�5d��a
�D�+K�	����S78 �r���b�L��iې��Vd��'C^������r[�Nx��fq���A���ΕݚiV.?��psq9k #,8�	ǎ+�'�-q3)$?*��oU��.u�3p����'�����	�(��⻸,7`�&���F���1�vUN����S[f��?���/^<�>�53a�0r�~Uwڐ���|w}i��=t��0����������
!,�N<^����ʦ?�]=z$��ܼu�����~w��x]嫬�GW���S�����t�✄�{�J�3M�%	�2��0K����h��9q�������VT��M��3l�$]��f:��8�pC,� �<u���O�����	ʜ���!]cYy�Ր�"=S�����P�'X1�c�Ϥ�2HSf�}�3xNc=x�p5v3��F�iu����6���s�:��n�%>�Hp���Y��[�{�bNHH#W>:����Jo���*��2���䙛�W?+�>R�.涅���r�^�VP�� P8)֥���NLGVo?��O����Z�S�.� K7'YI)W�R&��1"�=�<�NBC�r��Cplj�lka�!T9�0�U<��}������M�THM�N8�����1��+���"�y~^�Z�"�M`�><���C�c�b۾AY�Y�M�M�I�;����&❧̩H��b-��9H�KM+c0�:�^������}	��|�����{��b4�o���LV5S���͜QC��Ou1w�̰�ṉ覎v4���{���C<���������=�2��~�a�������]����b�7Gv_<���@���j xf��G��Y�2vlf�w����^�BI�t���|����0�9�WQ�^��7{��/�[/�N�,8	]��g�6������E7�0G^���������V�X���%SFc�ѻ�DP��`^�k�>4.�����Rl��PK�OT_\��zZ	&����~G� ~���a�e�&��'��_��:j `0}�`R8kj�P=���^���翨����_��eW*+_���>�V>��\,A�(���E���ތ!�1/F孨�幩���6�s=v�ԯ��l��<kϓ4ДcH��Z�����\ a��U�<�q����O�8\s=zr��Cޯ�|d���X��u~f�>���0]�u���t*����}1E�I:�F��W��R轅|1%D����`�����.+�4�7��ߟ��%/yI�ʚ�f��^�3y������/���_�6�� 9ԃٽI�b�b����YPV�O�=O:0��l����Ņ���ȏ=�h��ʛ���{���(�U0��$�;���b��0����\$��}����V>�Y��A<�`�)1k*�L�p���5B��exzWw����m=�ͷ�:|𡇇W}ŗ-^��7V>�}񈑣�\�9�����<]s�&_,^ԁ��*e&Np)BE�DBc:8S�*ݺ�6���xf�N�j�'�"�H��$�쳚:̼�U���n!p1�w�nÌh�]#{�A�Z#�I|���_��@��w����z�ɟ�ɕO�@@�ӹ��2��ꩧ�^Μ8Y�l��d�88���f�FIKRo������E�^��G]����G�_
�F��t�r�fq���Ï{�[|²4:7fꖝ?���n����?���q%�)x�F{o$�Ñ�}�,�/Ʈk���tڢ�F�h\wá���_�=�|;��o&q�LzDuRi5���AF|{|ː*�t�1�4�F�c��b�cY�s��O����bHa.@���d��Fæ�U�W��K�U\����ڥ b4LAo�������ݧt�G�g���f��L�]�|L���e�|����<z\���`\�O~�X��&��V����Itp=�YϪ<xIH�/3Qp	w���;+ǽ�� ��]/�������T<��m���o��o��"8�f�/�@�s���7ɣ�r���{۱y/�G|���׷����;
�˼����H��pUpnց�����.%��RI�{��jW��������piĺū�@*���\'$�"q!B0;FAqUA߼��P� ��!A����xؚ/��aqC��cV�>�"6�)��\��������m��1I�$�;1KF^E5��I�ybd0��� a
���l 	�Sy��lM��D��q��b�^����|����/oD�_ǗzHיJcg�aF�wy��3���wS3��~���C��O�W�C����|�(̽g���+����NX��Q�$`#@�O�~��pU�<���:ea'�M�iѓO���p]�[�ssM�Z����R � ��š{A�{��'���Ge�w���U� 2奭HG�b�*?i<K��}^�꾥GX����퓢�NT��y'/��8|򐯺�/o�XC�W7���=�I�����m8j�>l^��Ă!O����,Nz�p ����\BY\�+��dA�^�Ա�ȇ����~�d���p�'��W/:�{0�]\�$���w�������#�F6��$��D<K����ٕl*㣒��~�n枞ܳBʙ�:x�@DBE��0�4��j��qk��@*���a'�	f�*KM�T�X\�e|�ffS>��Uq��)��y�-e�����
LZ`w/�l����IR��R�}�O�W6b�N��ʛXjvh������V6��[�:&��K>�3���w��3\��[�n�!���Jg6�@�����\z(*ޅKm���R	�0+�EP�^�p��}���7�T�h
�u�my�$wT2��+�oG�c����l�ds����Ԗ-��L�GՉ ��}7����B�]v㬅�?L%ﺙ;��A�M*kUղ�PHѢ1t�g>�9�'}�'U7D�k�dIX��b&?�c@f�)��o��o�Al��=��YX
8"�f���ַ2�M5k��;ߥ���㝠���it1V�&�|G������`$!)���Oy�]]2X�Ay���3��g�E˳M^�W���Yj �I孭���`J\��:q��W[l*�:;�L��H�����{S�ʿU��-l�4�u'ܔ)�{��N�i������|Wwxڌ��_TO���V>���]Y�X�Ѷ	���?���6�XP���~���mA-&aM�k��(��1{]�T�p�D��>*ܙC~;;�X-�t��Dب�،-z@8:,�ihn���1�]̔9	a1�[H���������Ǉ����wv�W��6-i�ک)�V�Dz!�ɓ���
�w/�Ęm9����F����KM�PW�~0%��zw.�򭺏��덾w�]́CL���1R����@wT���27��_�,��C��y���9e��Jởr��d~��ձ�%�y���3ñ��m�V0ƹ�Y�p�    IDATtq�E�[Io2��g"������DE����Z;u~�;D��C�tԃ��B_  A�tT�k�g|�gTe�O� l������&����@=���]�3�X����x��|�^��1-��@1���>M���ǤHغ`�p��>'�tZu��ީS�)���
�3��OY��{
i���k�]����MYʁg��h�SO���x�[���o��֞�C���ys�M��mo�����&��� .���{�a[Yd`������pZ��Qm=�7���X��wzo����%w��c��`�T̢p�X�Ŭ|���l;�=��k_��2O5�Dwm*�Jw�v�L��A�!D@Jy�ePF��C�b֡1'k ����-�p����7���n$g:�N� n����� b ��4&=�qkWV�	�p��y���ş�3�̅���Fm�6&�Z���@�Q�J�gp#��˦�� ~y�C��5ƄRW#�D]0��0K�C��&T����y��G8�=F���i"�L��S��z�%DF�tu�'8��5�&�¨�6N[�	q-��ؕ &���튛�U��&�o���%yL��[��$�Ǐ��-_�0U�	!��Co���AtSMvK�
	�G�����OG�4ߕԇiH̋ M�kcn��ʦ�RH�4�"*�aj�9?U'��4�λ�1R���a4V�w������\fW`x�N��d���*����3��{��Ge	��=�z�y�'��i��Q���]���=�Й<��"5�Ӱ|�HZ.z0x���3���k�N�h�<�盲HO�~����W�Hs���6�,��7X�0}`�Ѻ�wfӝ�����~��p#dv�\�6������^�Ե�eTN�rl�fT�������'Δ]���bOv�Bx1�R�H����2<�݉�*�Ņ�u�͍9�s9��>��>$5G��3a�������;O�ܔ��V�Ӹb	����|n1z�v$H�Do_�
3MD�υq�3���Ҫ��w�b�*ͬ9�}���po�b�����-/ݜ�"&e�հS�]l�N��l=B�Pl�f�Y0̠S���~�������`�Č؊:d��a2�;����0��fEL~���7���a��N�������`�.�g�ٔ�8��l��R����q�8��̩�l� ��x4n���HW{��/d�k�F������Mo��o$co��>4���?��GR����lK���L�"�H��R�)�H�npk���嬄��B�����[��i��Pҵէ�9>��8��"�쇇&^>��G�&��,�!i!���V�֟��Mri�Z&����Z�����F�)�߿�67S.��8̍�+�Q!��NV�H/_�%(�3���9�I���H(� +EF	׶\$O�ϑ,8eq�$��J�Eˋ�3�"7�v�ӳ�<;��t|];�-�8{��HJ6��V���y*`U��R��A*���3���
|�j����r���,�=w}cex�3��_V�\<W�� y+S��b�V�=:}t�>&��=�sa�H��������)K�Ƽ��v�ܩ�jȔ��JJ��e*����u.��_V@�id��h&W=��Ne@I��c���9����@ʣ�{��ѹ�{��H������f�z(��?H�?\/W�R9KU��S� �!�F���=�����ѧ���Q7���m���b���_�j�H%�Ę&u� f)��u��?�Aˁ}\U�{�Y�ɔ�N��EB��J��H-Ʀ�|�me�Y[��1GE���b�\٬|''V�^�g0�6Mn�Xوq!V��Y�Y*@V������]ԣZd�!n�����:�;��f���CK�5���~6W�~���b����9�6��x.���d��?�W�7�t} T7�=Aؼ���Yw&�s`x��4��e�赳�fz���Y����l|y���ИW��pg�w>4�K���2� wzo���=�3LM-��9�{���|�~=�v2��O��������CZ����a�ލ ��
���5���g4NZ�	<��q���.w������/�/rH��u��Ȉ�F�=Db|2�x�U�w��rq1��L��ed��^��Ft&D��K.�dƴI��ߎ��3�E�u���I��ﺷ�˂i
��)y$ݷ�51���
�z�ɤ�SҒi�nX����ұ��xs<�߅0��ӏş�Ψ"���I`��
���G������Q� v/0��RlõΞS�-&̪&��=qӊf'k��ѧ�����Q�Dz�Y"øi:��	�R�4�������۲��7.~YH��x������O�F!��=��͹���^?sOd,c"�*љ
��r6���~����mk��l}{`1�	�=xv2Q>:�=�����k2-�:���0� #(_Pfop���HI��@���4���a��mne����t��?�>s����ax�;ޞn�^})=J,9�g7���3y�wbVz�K��P����I�+G�ə0VtPD�@��&]0\5�FOc�ы��@=㖭����s�3֘�}���X�Ƕ����$��]	zШ�a\� �@Ofܠ+tf�X����gQ�,�)t��{"���3�bf��H���8r|������S��o"�e	�����L&C��/�˧��؊��L�;s�ԥv�M���wT_��9�+@()i� P�u�C�F] ��j����./>0�Kr4>�����~c|��L�o�?��h���6<r��4��OR�Z�Vq倥36��,
�6XL����</^��i�s��������E%��r�+�gx��o�r�����F;YW9��#�2��������i&:����$sr˗����0�D5x�4+�2pԣY�y˭7�w�T����ca�>g�!��,ڥ����o�:�K��q�ʇ�Vf�4F���Zޙ�G?��;�Q�0	�{�k�Yaz�jzF��O�e8�	����vr�S�>;���s��إ3�1�Mdq���[����h	�R%m���ۓί'�O�/�G�u>�#��ѹ�����~t8�K��f�T'���R�ŀK٤e%��\*�E��]�����GO�S�}0*E���d͆9����{�D������".y"b�ЧtK�tx�@��I
#�6�� ��/=��lu��t���><��E�=~��񙅽s+K7<����qx�����v��n�	j{`k�o���������6]c���$4;�r16ɮ�!�3V/�������v����h3�5�Lfm�Dc��>�y�3��{�}-�w�+�̰C�97U�0N��a[ωR��=��F��e�͑M�~�'~������Xh���SqZ�f�'��>t��`9��U֨g�	�24,o���ն�����R5yAR}�ę6��-}#�/�~��X��0\�Zd�>�c+N�Y�ވ�~$��	Y�#$�hV�<ЛuM�#=�h[Ic�IȽ+�Ҟ��g�$u�R������p����|��F�R7Ds���Ƞ��T����y&a���t�`y����3x�i�$Ji
m�Ù����Φ+����ٽ3{�9wr���S�-��4��7�r��I򪃺��#r1Ts��}ߌz��7����1��O8�RQi�nW����2���'>e�=)n+����'����ު{I���Pp/�ш0�F�7{���ѯ2��Vgz3�S!�3مц�`)�V���r���s��Cs1�M�ʼ�������G���<s�Ԥ��3��6����#ێ���d��YK�Ӷԁ>p7c�ë�N�����c�{����f�">�����̗��\->�U��!�$�.2��
Bd���䱱�NY����}�Y�[����k'O��̆/��A{h�-R3�ɟoFR6��K��*�_��e��7�DX�Wc��㫑�����Z]����H�Ŵq!��}ss�1�/�LxaJ̠q�I��^���������~�NoC�JRS�����=9*�9�l,�ؿϞ9�squ*�'�28���icnj���ō�?p�o}k&B�H8���p15�Lo�5&7���z"�z�7���F�+��YF��4�e��2p�{ە��?�����K۟��>�'N<~8{�L�p�fj���n�p���Bή�>���GP4̠9��Wd�2���O��g`xE�k��f�9gH�j�1� yl��mE�9���G�sf4"_�����k���Z��	 a��)h�����	�����%�r�Y��)*jCt�c��0�!�gG?/�-,��ܾ�ӳ7�tˑ�CSQO�]f<HBL���<I�����2#���ZE�q6���w��$�%P��e	J_��'Oon�.-�lLL�Lf����ٹ��{������x��K*v\����t�Hs�2i�z�Dj�SzyI�H'�6`�7ͼ)�9wv}n{ϙ�3�1�������'w�N�n�D�����֞L�M��H
k�;�'���C���춘C�G*�l7���>&���+��]��̧�΅�&�{�o,��ؙ�Iٿmfyssgn+�O�XTM��0&-���d�2:���@�����Yi�.i6ih`�j�>뛗67���OrOl���g��������z�0MB��*u�,��X0�k�tS*�XEUx2�h]8��mtm�<4����,q#߶S�����w��C�fl�v�"1�.E�f�)/���P��U.�8A
e��6��t��0���T~f�2�����p�m���^��mN�m�Y?������d�:рL�'�1S�HP'x���`���tpfѭt�'�4L���0?+�U"xY�Z߼0�x`}'{O�]�ܘ�[����{�칋w�F߿�HA��z���5��&s0�F�lF
ܙ����D��M=���5�g;��&h+Ri���Vv��$��wi�dTǙ����'�/\���[/��l��,]�w��W�^+p���|VU�����1��3���qqq��㦓S�B���$�'����8����!�y�����`y|C�J���&D�����6��:S�p���M�ܺ���?k�#7]���_��޳y��O;��Ox~I|]�AZ�!䍉����m��	�����nNC@t0�8q���F3"�b��{��ژ|���΃�k;��V'Xߞ|8��^HCٱ�K��h�=�<�ԙ�;��x,��ݲ�l�A=~_��QA6�m��>�|~����2�����(��֧c�����/�용��sv�
>���-Ѕ<���ԡ�Ϣ>.?���]:��V�������KS{�]�
+��{��ت�9(K|�k�)�\Fw�v�#�\�b`h�Z9�H��W�6�� ���������}��-��0�}�5�K���!� ���������`Ez��fPi^����)�߰6�pxmz����ҁ�#�=���LMo����̜��B"�� {|L�!)��HF��b�R>�$���\�'\^�=��6������k'�6���{b~~��lTp`F�s�i7���z����I���3��&�U����yHc��u�ңŤ~a��օ����m=�j<x!������޽ϲM[��V�0S�f�+�1X���%e4����ϺJ�Jo��?*�Y:LP�� ���,e��g�7^��l"�ށr#s��[ۓ���Μ���3�͚�� Rwu�wM��'p"�$*A���i&-�E�d���I=��'��\��/�NI `p��жPݲ����&4$v�7�}]%�?��U$��p�\Xv>�=��V���,�GzڰᔣA�À���ș�C4pv&��Q������յp���nz�͜��_�ޞ٘��<�g��b�&Y�fg�lӋ�����5fV6GT0�jp5PJ#�p�+���tM����9Vzeckw{*:mN$Y���z$��F�S�/�L�xF\f4S�2<c� ��Z(�,G|��l��	&[����z����<�F m��~��]nw6�?���/��5җ�VT#�*���p��P�{�\�C;0g�"O�k� �5�c��+�.�6��[�%�I;Ƃ�w�=�xf����uUwC�4q\uO2sy�wn��n����͘��Pj6JyVi�>��\V��:5�!F!:� ��w��t�9�C�Mg �j�L�ą�.]��{�衻�3K�w&��9usb{����|���}WO�>���ѣk$����:B���O�~�zf�^����2�8�0O]#ť�PrIqM�]�ڝ�>�y��I[�]�!�s;��/d�l�`^j�C9�u�QM��P���x�iO�k��o��{�ynImh��ɴ�)���{k	O����}γm|��ęǟ����s��#/\�p��˧�w��cύJ��^�o�:���4��^������z `�<��5��iqa�̥���q'��AO��Z�鹷����_����s�V^F�|���F��ٔU���~�g�$�V����񇫲��K�]��m����;9�";�nf�y��w�Ο={0�*�:}j>��5�������)�H��#S�����a��k����،����F��_�ar��-7�\�V��.̬onN���w{hyl����e�S�졝��ǚ2��w�k.<��&m����w�1r]�}�;w��{���7)R�$S�]S�,)N�q�T�0M�p[@MӨ�?-�4(� h�(��H[5i���Ӱv�(�r�Rd�R���II+r�%�=�;s���s�^�bH�"��V�^i8����������A��kQf�@|6�駟NLN�H���|����f�TX|Y��<s]ŚpŶ�:�-j���R�r��6�7��di���ā��X#z�R�R�<Qh&����hK	f��{����}��g�]�w�L�<��(+�1Y����Ɓl~�c�-{����6�0a�z�x���M�5k���$"�S��㮻�2 ���W�b�
p����#��J8lZ�	�?R��[��`M!{43x�?w��333�v*[�����Lk
JP�e�f$3.�� �۶�+�T}�≉Y&+*A�e�-*�yQ1?=s�Tz���>2L1u�������u�ًsBL�m�`mRb�ǶL�vY���2�9dâ�s�,�����%m�R��._�|��E�2�׼��{�'ƚ��.z��۽�C�VUe��m��s���FǶ����d��������Ǹ�ey�Ȫ�Jg�)��#O��_K��ֱl��N��.�:h�����.-�	{0~ Š�r�};�O�.�-"�^��蔇�ؘ�V{ep��6Zu�-	��	������tqr����?��W��+ SX�_�N�W�.'��8pŲ�d�.����ժ����x��iYX$Fh�iwmɲ�Rc _��2
��z��:l�h]Qq��H-5ț�\v�=?��x饗_���6�7�F���o��9�%���w��O��jd/�l�8}��#�ꝼ��٩;v�=}���f�C����"W�쌡ZP3dbX�7*Vν8���[��8�de�:yR ��w���I�ڔN�.��fd�IcWd~� ��S���g����QˊmB@�����|�TP�P��*�R�R��vT��qT|'_�9�e��G����<s��lO�K�U�v���Vl��^����?��ta�B�M��{`!��}(7A�
C���(�j�mݚ�0}:�Ƨ�)�Zd�K�ۍv�z=){��gX:mUJ���7ҟ�X��X/���Û��2���ވ�;�i�-�	����+`	D�g��R��'�k�&��ʘ��X_�M2��@Q�e���*�,��X�d��̅}A��r���7ҹ�����z�����}�*�����?���c�^�3&��xO��.,�*��v�#�`�>\D�  �l�Vm(�� ��P�h[����/��WYJ$��l��BJY�8�@ 2?��(�  @f����I���Hjm�<��c^��.y���pə�T/m��=��� "��X[Pt�X�i�)Bn�FQ
�����AQ�oY#�g>��9�W�YW����K�)9dp�P,�N6����;�n��Gg���Q��    IDAT�JF��ܸ"d��������|簢7˦�{�>�U�wH���Fkc��9�C��_d�����p{�7����E��r9������l�zǏ�,�?�䟵Bnco����{�wpq�U� �H��2?iU������w ,@ @E��+5a������}�8wN�r�8 @3��4����b��k��`L�� �g��Ŧ�)<�Hy��/�ӣ���G�w����.^��k�Zbt �k5Ŗ6��6D\�ܓ{�"K���8
�N�I�p@0� ��.s�C��4�N�h��rgK)i�L��Rٿ��=��xr�9�֥�Sw%J��c۶ٱ�b�8�I'�6Wl;۶;�����~é˺����c��f<����p�+Nx�
m�ѽ����(�6�Qz=��^\(DE�$�(�EB�;hL d}~��o:�x�_�X��������`��`3�O����6�H���f�k�3s�;�p)��i�{��#+��t��9Nw���YQ9H��v�J[� H��}3#J�󹴘�0to�$H^غuQ���6Z8d�����`�Lt��{*T��te�˱��	�}zuzЛh�N�y�<!��m&[���A���J�%�&��
�	a]��.M�#;LD�~^�]�=�y�jZ�lo��쩩����cJ���M�_%��x���ux��P������a��"�p��T=�(wϤ�n~=i�u�`u�`�NJ��/
��؁[�x��$�}�aa;yU��Rb��5����9Am�{]��Sf{]tI�b�� �{����ų�����$^_yC���f��UC���2�������:j��M�@Mp���̄�rɍ$9�IQ��xrp���tUP��G�PTU�VF�'��r��d(�!�p`�q�2bH�9CV�!x�.���Z$�AA1����L*�<(|Zb�>�)�X���:�F���җW�*�.��WBW� n�ƹ�7Kg�׆C��A�%X� �p7ZLL�Ʋ.�97jz6mjdit҆��u�����n~`~�P�������Р�g=O�p� }�3�ub��#��m�1�,x�M)��M��
�b���1y�
ղI�G7�L��.\�f3���SNJw�s#%��2o.��P���^��1P	�l�֩���Y�(�^w7�#�֕F$�_ή$N��{�R�.�T�J̠I;�x��y�եlſ9�5�j�������;����0�%B�zh��f����|�K�7M��jH6Y�Y"�XG�#ѹ?�ތy��D�
�e�k�����S�A4�J�)BeQf��z�!����������4�1X�کzB�g��\����-d��a	H�G�@�8u;������OHi<G���B�?V����6��D/GQ%|�	�*]N��P,j!�D��f��/r�1�鹚�;$�aa�nا��� ���t�C�����<@��a� ���ǔ�����D�xvv��K�b�����>��
�\-��4\��5������ {C�!�D�Q=B�W	�T:2QD��o����o�[O=�({+ǲ��k�~.�x�ƣ~����f��V2�`@��7�l��%������s(��z���n�.0�ٝ<�+��״�=`\��W�57?����%�e�l4S���~0"��ZX̜77F >��BOb.75���]��{���T��~UhVFq�d�R t֑�)�*3��c�U��0��uQdE���1��ڵ/�C� �IU#�gg*A#��K�� �-?V�L�&�5�"�2P�D��X˟6u��.s^�"5\[شS~���_���Rb���,H�fT,�`���!�x�O3Iw����Gr6�3$8|��D������`�!�N̏�(�������n6{2���J���!5S!NOh�Ta-��o����u�������
��[X��?۸�~啖 �k�[2i<P�̂V��<G��K��É5���FHǲ>&Q���u0�G�BE���X��Ua�f5��#|������}��Pa� �n�}�/�u|�2��[\t��O9&O&�+Lhd���rH��\���'�AX���n�k�5ĆB���g2M�[~� �a�qy��.c�����A g���������̉q��^?	�.oYBe#�O^0��_8�m7ܗ��ۦ���K53-^2�`��$1�M���M�w��\ψ����qect�䝤�i��}۳�@��r��ي��c/��C�/���o���n��5�\hТm8C��A&2i���tEi"���ʠ%���>��b��~6H�`@����.y�ة�d�n�<B{�攊9��Hb�@iS��C)�l���R���Ur����a�{B�ru�����K�H�0�*띃;<���۩���K�o�6َa�8�I�[����/����y����B���y;����QOM�t8�i��/I?k6�K�BXb�$Q�զ����tb�
]
�)���Z3>8�6�o�aV/�Ŋf���2kB�Æ�c��k|��մ,ސwR��$
���<�l���M^���cS��)�t�㎛g.�!D��o4�-m�%�!�d˃v0v�X�v},��1H��1!1uN{���>G�tz|Zp��<4�ۤ�t˞h�(�;�J��P�&>�F���1��m4�$l��2M�%�)��*J���\�&^˱��*Tk
"&Eޙ%L���u`z�;j�����	��SFQ��ˌ=XK�b��������2XM�a���$5!�jd!�Y��0	�jޓ���>�������J��W��;���7TD7����!���������P.��f���T�(ϷE}��t^�>C�����zG�pȭ���z��/�_4\s�R�hqD�,���A�ɞ�(���-뙨�����0�0&e�2���a�P��Ź*�dQJfy����_
z{�)�z) ���=V�+���U�Q(��Tsّ=\����ƂsLP� ��%�Bq't�Y���|�q���6��|���o2�.l ��ńQ��V���`��޳"3:�p�m�W�m��%_h�x�����xB�H}�ėT)`��r�2��wD��a�5z-��W����-��mG��YM5*���Gbd�zA�����JU]���C�c7����;ClXV��͎��6_�+�n��[�A��l涡$mh��6e�v�|*,��::��\��`+�|[��R����:d��Tn8�"�?B�#SddZA�^A*�( Xp��rQEv`���5�2 dBt��"�w�.:b�8(#�m/8�E�
M�H#G����I���*�b�� �(�^nͭ/-�(����yR	 ?�yҝ>��Q?�w����B�I187:�e�>���mE3 S Z��k K�2`��k��p�akBI��1�k����EVmO�\#gO�/��83��͇�a���m8I�y�̔�.���Ի�'�d����8��5̣�0S�ծ�������Ξ�Dz��v����ʽ�	Kus+�Aq�'',�Jbp\!e���i�W^J��(��ӦI�ע�F��4��9+��F
aO�jQ7��W!��:�yf�$i�S�πQ��2�Y��hk���U�QY��A�����6[y-����0Y�^ngK��<�G�+
+%N�a/�w�)O����fՂ�L��*����G��>%)>�V�ƆjFm�o@���˱��'�j�є�t8������A�z���]�-q�L*Ng$���@J���y�3-���l��pD�e������Q��CiӲ�C�9�W`'��l���y�-r�����2hEa ��|��6v|�S��tU�-���uܢ���v�U9��H�hP�7�4B��1t�(̈`��.�I>���ݶ5�x�2�w�ni�<��`T�vғE�TSi'�;�2��1r���uS�S\�.r4�R�~��+GA2����@����ܽ�2`�����v�R��'T6�β�[�:⻪�x��BN*@g��Q�|:���Cd$�w#l�zC��n�������Ae��D��(����$b����	�&5��*ϋ[-&CK�W^%Ï4�-�a�0�^��`���d (�MON�;�n��6���ޯk�Φ�U^C@��q��2s�2��7s�;'�#֒�܂���|��|đ����ոu���u�Xb��i�+}]e�=B�Ș7�H�)|���*���S��=�oz��~rdr��kkUo���TJ����T_�1�d��M5�Ũ��ͷ���$�`ձNg��xz��!p��U��,�Q�v^Fr=Re�%-��G�]Z��/kguX����=��'�����e��U��9y��u�)���	pQ�Z��L�0��tt=lo$�[�ʳ�;����`=l=���f�jX�aOHՇϓ"Bb�z���w�[R~3}'�NvL^QjMf��lD�Ɗ
��Ϣ��r�4�i��}�d�`�r��~a��U��)��V9�i�qy�5�R=R�+q�ɻ�ʹߠaW�)̙Ħ�{�W�H���	���\q�3�K��~n�E��-2����:[�H_1Dוt����������"�ܥC�ʪ�[���.H;��x͵���$�����;d3��u'�rhA�;+mwtO9Kj�F#_�b'�/�dN��X�m.JK�B�Ѧ�[�]]qM����]�1��̷���8*����oᯀ��7���lT%>	��1m���V�%��y�&������"m<>ː�Ȕ�!~�ȷ=�����+��
w�D�����KZ����6l@�F&%�4��N�J���T��b?��ߏ���Z�J;�wۢg�+�D�7�U�%BN�7hg"�и�իfXݲ�����x�EC+�}����sK��(S��N?���߽�p
+��%�x߰��ˇ>I���Ŭ�΋GE���{y�.�'�'����v��g;����R~-�9�Ju���@ֈG�&��] ��q�I�[���Pǡՙ%t��j�0�'n�W�cK}U�.�06�PwT�ڽky�5�O�+^��TMϖ�Ï^w�Nl@�ɾ^�j?����<Q����*�8Sã���~��d��c��;��M�������G5����r�p�ͬ}��~�~�Ԟ�z����3e�spF�Jmz����')בd�Zʒ�@��Ƌ�s�d:!�/��5�}��g����nvH������;�	�n
9����e��bڴ����#M6(a��K�F��{BJ"������T����bn0���a�[�M�仝���f\eemI��K��p� ��Q �³P-BKfL�B	Zÿ ٲ���8;�]2�m;W��n\K�RQY_�R"�p�Jy�w5��(���F�+WO|�5\r��1���l�E�Y2���^܇�`�F��ʠ2�:a�/��jR��m�T-�cV�(�@�Ռ�s�������f�C�_�"-�a���.������J�'�Q�MԴf�<hPS �W�P�ǧ���O��v�^}���J;.-�>��G�y���Y�H�{��#o��3�D��ɫة̫F�6)��$����*�vuT��j����5$f�5C33�&;󚙝�)R~HA!�'cf0I˨�J�ȔT�����v�o���x �@�YHa��f����.�O������k���<���L�,N��l��lI���j�>l��*���.���	�� ����0��Ի����C�6:��ki>�"��ע�[cCM0Aň�6�`�,��Mm��D�dx�K$M��&d�*E�w]K�K޹"yL��5n[ʌ��A6����+�� P���-�q�6h���4�I��ج5�'�=�&@o�U��y��DLB������;��:o7m�����o~�F�C�,�,�B
>ྌ����,�%al�e�����r��څ��?#考̯�=Ws����d����%�BO�_�OM��ë���K��6�����5兓�$�Y��_�c���;S2Ȱ4�7�s�/ȣ���IS���dx/d���v�H��R�H�F^���0V��ȏ�w`M����cF�`Y�C��\n>y����>j�,¼��8X4�QE�Cĥ8֛H;WZ	?I!@~x�8��F\�\M]u��`]T�o;P:�0��yE�d���|rĘ�� ��_��]40]\���.�ktO1,��, ����k/P1@�m��:�K�`
Ҁ��B��
M��b3|�v��,���΋���4�D!��F!|����6�pza\�%E���l�i�$U8D�Kϥ*���<d��Ҩ���nD-aRwE�.7aƏp�����{Z~8P_�ľ��N���B�b��品�B���a���L���ז�(�s-n�aK`��B���8j<E��Z���בJ	������	�%��﭂U�u�<�|?�bz�#��v�?>r����MA���[~;�K�
�m�p��3a�k�̬*6���l�oJW�n���=:;Ҵ�p�Hb�5�kw3?�U���ዳ�$��7�M�j'�q���vȚ��Ӧ�#Zz3>�L���$
��
�[��&7��E$��鐺ο�1����̠��b�����]\��'Us��/�ش3�DM���4�_m�M1��*� Qw~g����n{��ɪ�y���Ǚ��u�L�҄ȣ�G��Sn,5ÚX�s�_�r�dbmӗ:�x�6������'~+����Г���LU�.]�{Ԉ����h����j@����'�.y��x~�	_����MAsñ�6�<�o.�??+���Z� l����l/��R 
_�1.��x��ݤ��bVM,��Ҧ�} {�yi����+w-J:��'ko�|��#i,�j�8���qfhn��h�ٓ�Ԭ�{�a@B� �F�e
6Y Y��̷W�^��~�R3��St�M�Ɇ	z}�jw�aG[	_0+O����@0I��ק��Co-��X$ĵó�G�������?���d�"5�R�3�1�����ӑ�@��Y(��j�'4��	����@3(^bܕt��'qC��K�c�EI�Fn�����q;t��J(�t��N�ǭAO�$��JRO��'<^�!mXL����q�e���(�Q*�]�1��tC)�{QY[��y�M�/9�|*�t�QF����'��!fl�VK�zS�'�fE^�)(-�S*���q{H��`i��=�e&��֙I��l2q�zT5!���.l���@�	��޻n��&�O��1$�[z��=h|`̒��n�%�����7�,o�:V�ыB�
լA�`�aW=AZ�$���X���B���=`���F㚜Z	��T�i4�:vX'���!�R
����<;"�_�+n}�a��AE ��5��t?D��5��4'\��K3ɋ�M�a���y4O d���J��j��$nǌD�g�E��)��"�
.i��1��ޟ�Y(\����I�R����v�a�˞���x��TΥ&��`��
7w�g��-���y]h��1;�p���F���\K~���&(U&�<ᴤ����\���C�Hװ���4�	��d�Ȅ'����U���*�]�`j�
l������5��IhX��G/܄r�7>������Aoul�v�3��<�% � �:j�:����F5Kq)Bsc
zbڤ_���5ɗ� Ե0Y>��)�T�<P��gX��;��0K`2�]�����!��:��7A����`�,Y�A=���W"nC'53��,{�Ȓ�lD�F� Ib<OHA��tk����pܪ�wL����:�k����a4�K�`I�i]���v����E�'�Ze�@]�V9=�����dzB�H���g.�B��S��QU�+��Y9�9������Y�NR��t)=�C��
1�$�@6���/f�&hݼ� �̻C_�`mȏ�|�}�+��j
�d��&&~��V�]���]�/s6�S�f�<K�$s��Uڲ��sJ���0���C�P��̞J��|��2)�y u}s܀S����c�X܅G_}���O���y�<Q!��,-��?bgo��Y;������ []�gw����0�tĴ���Z�d�d�O�O��uQC/8�՛MN~���S����QW�X"�D�'��	ٵ.9���%��Xs�����/�Nw]�L��n����my���v�;dCF��C�M�1X�	%8�}�*&L��7�g �4�4�Yc�b�J�8�����^f&�vz��>�4�(��İ�|�	�@���Ƭ[�2�.�9��/�<��*n.���f��%Tg{8��I��.��D�c!�A�PRM��j�<�T�_�A��fG��U�*T�;l -�/-��*k��K9P�����^��j`*b��iv��IbAr*��y>aƘ�
5+� �sW��6W��	�7���^?�I/���}"ژ��.V|<:!+7.���r���^��Rk��j�02F?0���&��*�1�5�\&]]�+�|�' �\}^"\���C����
��oҚp"ꀆ`�K�(�7%O�a��l�����հ>64A��&��l��ee9q�G^���W��;�us?l�ɥ��1;-,S<���)���A���z���s:�f�1��?G� zd�O��6Ć4��zֽh���a0URVn6�И2�9��_��{)R,f�e=l�/���#����ل�����ʊvȂm��Ts�=Oz��B
���Ȑl�P�,���*��,DN*ZU5Q��>�:bXj�e��:O6O���
�|�J�6 L�,أ���GkϾZ�5�^\س��j�xi4x�aA>�T�zE��)6�&������%u��oy߽�ч������wF�K~�:���}
��[��D8��7��v/������U���L�t1�3�t�KT*�.\[C5�7�g��f�:�f�-@b�k�E`A�*�sd��o��%]J"���z(���Y��+0�w?��L}�7N�����x��GI�t��^�����Xmb���	qw�� 8-�9��1��j�����e�m��xUM&?2��1�⠋Xo���LPZ���C#o4Su�Ip�?u�~mg4�qb,..�9ΗKսi�XU��7⯢xU�ē�l`�3T계�����Z��~���i'�|P�T�+j׮�c	F��u��f�4�h0�X�eb���5����3�����4_��ӵ%�\bg\�� w=g�$�������TVR���8P"��䞂,�����c�83��qU��S���PC6�2<^8�{�6�Z-��y쿦ȋ�P���1+V/P�:�}�s�������,$��TA����Ocg��s\�=��� 6H�2�E{�)S$Em�D�k2�MeY=6�Ϩ��E=r������������	���
��	AG���HF>Ӵz�u^X[ȟ:k�.:aybl�voΖ�eB�E�_�z1�(�߾iB�O�@��QCq��V�L`���rD-E�b�r[�7�t���;�ۈ�^����?��K�n&:M��� HB�-�cқ;6^�6��J�̵x�����#�,�?��?gHy��'7�c|�>X�t��6�6Vr�.��9ӊ�Fvv�ˑ��L��6&����?��s�RJ7�H��J��b@�Lqf({��֨}Z�����{�@`Q�u�)��y(#A�n�����6��1�ы}cd	�!�	\]?�ǹ���'� -'��G�j�}DpM��P3ETw���x������^}�%$
J��7q�{6jQ/�b/'O��G��3֖X�꽟�����=A�j�b�! ~+�>t�
��=��l�@�`����Z��[�
3����=��4%��B>�C�C�#��Ҋc�S����э����l�*
�%��iUHu�3Z�#�7b�G�f��~��~1iA>���f"{9����V�톼o��5����>:�y)),LI����CG�֎���8�f1OO���m�&�7��G����	r���c�9�B�A�CО��w&|i񢒹ʹ��������ñ��i�闱P�d���P2h#���|�V,)��[3�����@a�2�)�������h���Â�<��zD(��D���̐H�F�X���Ԝy�T֠ՇprЎ�.��@:D��L���'g��mv����qanv��}�����
�F�^�fRi�d�\lxi1��P��+�| +�u�j��s��o��kQ��V�fR��Tjxim����f�q�&^�f� �B�JA�
�&�@��پ��ր�J��#"� (��"� �;�<��X` �؉0p�?d*@�&�LP��c�G�F1ϒ��N�i� ~���^J���n��:%�U��%o%��h�;x˔]:,g{�H �P!(�^��H
�?x���y�#%[�`�/��#�?aWuI�UY��w�͐�+BUg��TJ$,��I�ߌ�Ҋ>l�T5�C�V!\��<�z!�iw9U��/"�?�	��#��$��aK��1��4 }
�$g�۱g&�g2��B���V�"��)��j���W`X��`� ��c�$�t����I2��	�W���=�h+�41 ͹�S��B�v��A�!GeM?�s�Z�k�����Y�8�T�X=VB��9�d@�$�ԾLFυ\ycei*
^��Llbߴ�\�B/�a�5f�W�0ر�1dwi������/'�9����9��cn��%zR;M�΅���1o��i���K�XI�+25����6�Ae3V�g麕I��F;��Ѳ��J_����0�j�����5��ܺ�d;��j�`@k2	��`�֚)z����k�4�C̓T)�a30ǔT����~A�;ӵ���uϋ���Ș-|���:'{��]c7����*b����`?M*��c����9�j�w���]�B���=S�����VϱA�.4���?2�	�������2�GU��/�Y�D_g����K^7N�OO��'GQ��a��`c#��b������Z�g�l躚G�ٚeT�O?$H��f��<��GY���=����74�ۤ"��
��@��y�3Sה��q}5�[l5�K�6!j��=�����o�t��*���f;ZV9C��/���S
,�+ #�Lqc��F Y/أ�A�c̀�Z�У�n�ov�*W�El(�01�8��6� �;���l�
�ҋ*�uq��6�8Q�1a�ID��/���{c�$T7�'���0|���{@��D�0�䰉{��,�1pp�I*R�H�f�ş#�x9Y�nujab�)����6��ā{ c��_}	SR�b��Ճ ��}'�x%�H����y"���h��~��-�ZS�&�p!� !V��u�j��:�bK�*���y�7"U
5�D��}�F!��u��Z�*_mN�Jq�ke�\����|�Ċx��W����X���#	&��L�$w֩~<N��\���GL_�sZ���ǧ�s�*R�\��Ъ�e�*��:��"���Ֆt��0�;N�m!3I�j?@?v�P�H:~DK���"A���K���o�Am\���%u�j��\ދ��3�}��dq�W�U�a���X���rz~��c̠Z%�փ��i��pg�E�_0%�\p���X;ђ�.	ѱ!6�̄oɁ���~�F;0��{�D�"<�y;N�a�hF��#��}A���Ұ���r��`�ڞR���F���JǬ_�c?��'r���k�oh��`�K��델�}*�E�=��ᶨ1���|�*�iTn���$���x��#�m�������aǎ|��FH��$+�sQ3e�dХ�\���IѲ1"�?>��u)����Ĵ�6)/X 3�:���$΀򯻣����� ���8̫���N(�P��V��v����r�%�K[�m)K��b��������R �����_��������:.BmɎ��θ���i�-�y@��W�s!�7��ƀ��A5ȸݎ̙�ń�hb�4��9��4J�/,�y����-�y��z���kh��$
.��iZ�)�h�pX�5vNpV��G���x0[��7�tVj��D����/I�3�. �7H(}ͼ	,j����hx�q��OK}| #�\�l}��^�y�&G��?,�W�Sn��TU�g��	%B`���Z`��c���]|�1+C��3�8r�>iW�)=���a�?U��׉YT�r,�q1��č�k$�4�t�����ӣ���
o-�W+Q�ԉ����*C��z��&�7�qq�c���T`e�4,��zX�8������	<��\H}�7���d������0}U�&dE�����-FG	F�˩�����+�F��ؖ5:����	�����l^��NT  ��T�,cHzs��7Ե�40G�d_~�@��^�_�<��3S� �c�l D����ȹ����5om�G8x���4�� 6'��֒E��!�Ú�����Ϥ����r��'H�T�z�`5�D�?�#�S��%�U!�&%ww8�<����O������ѐDN�:��H3cd���|�&;�����C��v�Q	V��Dtl�qTd��bw�e]I���E�^�)�!Τ���.�b	��2�RҜm�r�~V���y�u��/�Ou�l,�;&|8���Ο5Rk��1tkΛ�p�*6@ƫ��y\L*��*i�%�;��������Mk��
͚dnï9im�(D4b���n[�9?W7.P��7��6��Nu% 0�G��WT'|
��p�#MW��*��X�4�BS񈉕�v:tF,���Tx#i���>�H_O��K��(�~U��g����##�a��l?�� e�g��u�y����)4�H�^��h������3NU; \��
��l��:y�D�`�����unlc���4��F�"�:Gխ��^[,��;L���(V�'1��W{_O��$���m��i�e��Z�m����Wߺ���j�L]�u+�Ꙩ��a��sZ&<��G8�6���E��?�>�;m���X�P��9�Jq��W����bH�y��HW��~�u���B^�M$I��L9LLUh�jQ������%�Z��@�/��&�[����=Su9(�A��D��q���v˩� R*��2�0`}"��V��n[w�b�i���躞�%&������<�����Ƒ��%:�OE�S�y_��|?G��{�(�ԦO¿�g�1�y��b�TIA sú�i�t\s�J�Ū¯�j�����?}C}��ǚ�}t�gÂO�un�4.M�% X�_����?�����u�2fD���LSg�8��\��.2���y�T����s�R����a����̌��/F�;3�7�Ѹ+{���#]�۶y�U!g�;�f��.�ѲK�@��[�0��H���^^>�%Ha�^��.�Y��r:�i�|b��t�ۮ�M��me��M�T�w5�����G�5��T���Ξ?���ݮ��n�9�"�}��[̑r�+c2�4��t������R�ǽUi)��&����?.�q+}����p��/l�LA��]��F��u�_k^��U�B��a��\�G{�xw���l�}�{���ZFj>j�VH�W8��P?�F������o���k9�Npg;+�ʉ�&o�Y~N�]pn|i���*�}���Q7/u����s���| �B���.�Y掏5����x55���_�x�� S|G܅ʶ�R14�ߣ�'�ܸ��۽��n��'�_����:�$��5u�(@H-7�OQϤ���[�z�7��GR/�80ʿ����qp�?ӈ;�g�����rz�P�ޖ����y2�K{�oVo]&������s��o�w�YQ�bԥhG�K���K1�܏'��s����^�-�"�4�.^�~̫}��Rw�u� �T =����b����|w�1�򫌻��[�:�)l�ޤ7^�.�����
曮:.֭m�g�5m(�� 1�Q��ۜ:�6�>#{}�n�I=ob/��/�'��Jo@SFn�-���5��Z�ٺ��J�K���6����>�ﻛ%�E�,�(��fA����Z��˨����v��J����MMmE�X]���˶{��+�e,�g���%Zl��Y�4�N�G����x_&ۗ��vU��q���y%_ga�����\��c��lO�w��Fk������k�E�?!��-�l��?���4Fybsrsrbcu�Ȉ70�Z3��]�r�5�������N�Q��\�<���V���ȵc�����۽�+��<��¡�ӦϙY<��F�O�F�[j�Q�.aC����w�����]��0F���l��X˕����������T�2�O ����Z�X�]�8�e�	������S��Y�0o�f�5~���U��ѻ�]�h�'Bi��z���N�N]~�M '�|ҼZZ�Σ��#�Tߡ[�s�(Y�n��7�X����yoB���������-��B��}�%���>V�\����$eki�h�V�s�me2B��ll�@���˅+pÆI�ip(��ϼ�����M7;�:��\�4)U�:xŊ7���Ds�m'^>ꢼo�b�iv|_�F��kE>NQ�4̾JܪܵIjj���Ճ��w�H�50�yom}��ysH慫�hIAK���緘ʂ�@�?��E����w57>��Ыv�E��(J�����%Gf�c_W�v��M�Ɲ��;�j��X�λ%*86�;9~�f1X�#��y�)]U��KnpI�R�|��� }�1�J��9u"�3��L�Ě��jl��$j
�����8�w�����8�G����MV�g'j	���r���&J��'&�h �o�J*jō��PK   T�(U]�!��	 &	 /   images/98931e0d-18f3-449f-8fca-8d5f6b2df0a7.png -@ҿ�PNG

   IHDR  �  
   m�y    IDATx���ٯ}[v��cι�ݜs~ݽ��U.W�U�I0q<�BB��_@�ސ�0!!�Ȁ�O�Kx �
&cP�8v��n��~���Zk6������ܺ.+�����9{�f�ٌ����'������n�Y��J��8"�� �ϥAD0��96�g�5�CS�)� �B��I���|=Nq��������eJ)���ExԦϷ�4L�Rw��un��p�ֶ��k����ᚇO���� �n��ϟ�{������נ?��&���#tz����ܟ�O���~͇�
m�МhT���������q��8�9�[6`_y�旿����K$���S��R�X�>�ι:����¡/�g����>NHh�Ϟp��������>�Z���n�0F������[o}	�z�,��V����X�����<�M�Q�BɅP���;��ۿ���a*D�Ւ����_�k�����D���%Թ��ȹ���iN���G�2M��	�_�w��������O^���f����~��_�*��_�m�]Թ/����E-���������_糏>��O^��i��8e�Ւ_�/�K��� N��ϱ?��<8��y�Ա+�����?�w�<f�q"��^]�ą�����S�տ�7H�)@�?���d�c�p�ه����_��|�=E:5..����5�޿��o�;��qn��)�������D��s�o��o�;����A�BX:6w�a�E����_�����i����L���b?��B>��9;	�[]{���A��m�S�������?<
�����������O������Z��t4*�?̌.% ��s *UE������z�@L��3i�u�c�B��;T�T��͌#)�c{���L���ʱ��qϬi>��?���99_�y����)?�w�������!����{>��g[�Lwj��?������?|Ϣy�����M2�/�Ə�nu�咏��,q��E�C~�{ﾇ�|�X��3OΙq��Q0�@��.��D�@+�8V"�@�>�����	��9M.��ՒO.�ay<���������'��,It�����G�{u ����{�s�������\1��/z>��w����'Jp,��i`������3:��NY6-ӓs�s�<ߝs����"u��s�up�:np���@۶�}�j�`T!�à�u��p��)H��V ���WG��f0�Sf@O)1���l4MC���^e*�C����ß��ID��9{q�`?l��-N<�E�>��1M�z��NA.�?�!M9��!�u4MChZL;�T'v�{�jޜ	!pp����Os�r�ZB�kb���GD�l6��s�9gb�x������9��0:V��틁������?+�����s뿎?��oց�{Δ&\��JA�Be�L�y23T�8o͌\
^;�i��'��_��Wy���g�8 iē�ƣ�kXh�1Bqe�Ł<l��8��Q��� j��?�Rʣ�v0&980���@�͑�9��hm��=��p��y����Ę�J3D/�b���Ū��*9g�e�v��H��p���V(f�\�C7��ѓ,YA�h�R@E(�g�3�!��Ӻ6f�n$H�֔���ɑ>�X�K�BZ<�G��6gid�O�ֱq+���Li=�������&�6��)og�%�5�!l�R����,JD΃���52��5{iq��#��	�)�:_ssǓ�W���ػ�\"9O�����L-e}J�u�b�#t�(9�_�l��MN�y�Z�:�<}�������>O?��I$Wh��5�+<�"p�k���u�U�6-�TGl��m=�WW,^}���a����䄮�Q��p;�����iK��	�y�E���J�{��A� �.`.��EB���eh�;�1�����͆��Z����(�ϟ���߽{�*N4>П�V�ZN��|��4!u=I}~J	�/�WGN����m���+޽���Ś��^,{l0���L�z������4lp��( %��� �� ���Q�^�%M8Q���KfѶ�|�]L;Yp�4L�kJ��I�[+䜑�%�@����՗�ia¡fx�F�f�*d��V�BbX�d2v��������k��;?&5��lw�_b�5"��J�ju�T�R�dC�R�s�<�xJe��)���J��A�)�!���{����e�Y^N.�Y��D ����_u�w������ ��*�`5�
i���9X�3���z��3�6C��6=���v��9ЬN�1@���6�{������D��p���,��_���R�88)P�ζ*R
��{Oc�(���eČb��8y�^�q����)󑢂D�������xþ�&%GҰ'OC�#����3yHÞ2�H�'�͏�<>灙(���H��!����ȎK S�_�����~�0�ȥ^�6;Ffz�����Rp��?��Da�6��h���LUi��64�l�<�(�.��u��#��<�8L�
�Z�Q�N�%=S�G� �t������c�JD��-��,�5���J�~0
s=~��M#���>y�E	�)"���EC(lF?G� ��B��%� Jh�㖋�s����%˳s�O����m�oZ�6�z!%C$$��8��q�R����q,�3�(cJ)�Zx���15��"x�a�n�D���iX�{|�Rv�q�1��r�e�G �T �q�F��Ǒ������q��(B�z����BO��Y�YOgK�B!��{|��o�w���2�W���$���"%Sr�sCE���8�h�5y�©g�Lm�+kRtd'����!���Hiq(��V#��=�J�IΎ�4R�2ىe뛆M�e���?�a(����P���k������>����(�;Z2L�lVYw����v^�s�B���V�g�=%f���i��ܰ�J6�У.��ړ�����o�SI�I�o��
i�����o=M�Tv,&$l�g�
�H]��OLˀ]^�b)|���>e�V�gn>����7��/�\؞�M�2��0�ɶ�Sh��֪s�&�tX��BSY������9�A}��Me*L��{���W�*�{����u�����'��u	-�=��N��-���
A�]a"P�PC����;���h���i�=9�=�ח�d�⑒\ype=ʃ���))f��Tɬ[��^t`"�a��2R��;Ԗ��-)*�x�,uU��Q�xw�a�'��b*Uw�E���q�ѿ��#Y�T�Xp)�c��#�<�C�������c3\��-q�æ=��7�Q���q�>G�'�'���H͉kzL��i&})�9��t�s�&*EjD T���n����@�׾��E��� ��X�Tf����M+���=)H*�PꠗRj?R��͞���c	�$#�4���RA�ҌMӠi�j���L��q@��z��R$�B��K�"����������T<؄S��r�i ��H�Վ,U�Qr�l�$gR��W��-�~��|(�GWk`q��#��4��SBJa��A�a��@�7�#��Z١8NL��J]H�F̔�����S���)�nO�7D���/B�����I�
*F�+jR�nQ#G'�O[bP2��y��i�$	܇�Y�%K�8[=A܎m��}��2�TC��`�w\ǹU��3ͬ��AQJ�`��&�("�3"e�H���z��%�W��'�GN��u�RX�)�����ˈfJRd(D˷�!��
r�HRS}iJ��S40LJzñx�-��r7��c����mb����G�2F:����H�9�����ȩ�HD1L4D�$w���A�'��jV����2�bÖ!��#/�������]Φ-�tS�\*���2V���5�H> }.5���I���_.�B�{��q�g%QTx�8g��m�4�𼅳�>au�)�*�\1�:�:���Uj�f��8���!�
G�o6��c�qN�Nr��H3�tH_�������LNɘ������t쬂�Y�����U�E�,�90
Ց�5s��1�zLk�pu�+i��x�xWSw�M��^������ih���	�Q��H�����]S���
�- �B��_G}X���9��̱5��ʜ�,��� �iCjxW�Q�9<��ӄMK�9�h͎��)�gs�@�Fˊց-��`OΔ)b�c]@��ޮq.� S�)1"�D�{���i�aӈ�T�-J��˃$��r,��懜��+�)3����I,x��T�C����@�S¢cS�,H)�q{�辔2{��}��!M����*F2�N� )��i�F&��1�k&[��(�X&皟wyä���ɒ*SfJ��Rzd�50�K���K6�;L��������2m���Wtc�"��by�D��ip��]��x�A,F2fM�NqM�*��٧�ݰ�����D[�Uh)y"O{�Ғ���c�f+�s�M���H�{(�)��c�IC<wi8�s�9�c��8��5ۻ{�8c!�X�i�;!�H,5��
3���ց�N�J*JA��Cihr���!wlr��.r#�ɱ����������y������2����Y�Y��a��i�@��>�ɠ(W�@5�#�}�b)�7k�YaW �Ґ�m�+���B��7��>r&욑\W�����ë��#ku|�S��h2��v�rOםs��5�x���ed�:��)�A�Ú����"�R��M��g��
 �Y"�LJ�7D�
�S*t�y�l�{��Ȣ#��0l��e`c}�w8�"~��*��H���3Й�us��#�L,�g3	��[�goٍ��zh�g7-(���j�8��H+�q_N�̟ո�vXל�ȇb9�áu��:�@�����vH���FLs��@���ˊ=��]�'ل���������jKƩK�N�%WG�L��R���1IŎ��C���?\{��t��Q[SI�YC2eQ��:�mZ\�&��g�{T�Z�oq.�B�oZ��pQ�O�"�!~���@�5�m�|h��	�=:e�i�0E!ˈ�
T������l�����#�s��^�V4DD�\�XAb���I!{,x�GHӂ��-i��b��ǩ cfX�J�'""�9_;�j�U�'�>�1f��IumP�-��=�U�LR�?O�����Qn�$�:.���r,Vʿ�VY�jl���w8[�k�9M G�U���x�@K��9���T�\bҚ��
�(	�~�m�nɥ�٢�BpӜ+w�;����Hβ_3�ݱ�r.���9��}�ܩgg���pm���RY �"E��
�2��clbh�H3UUT����_�\a��xJq=�a˔�6e��{�i��	;?ct-��(����1/i
S�(M��-1�A]��J�25kr2T�1�K�:z9#��G��4���HQ%)D1R��@��t�-Z6%J'��H�| 9�]��s!,:.�>�iJLW��{̈́n��k��&�{�&���kmp�XR����!��W'd,��N��s�S戻˽C���s��dX�T�y��=>�X�l
c��ə�m%���M(
U��Jc��v��;�LFJ�X"��&��p�%�ἱ����5GɁE�bf��#�)2�¹_��0����/
�֥=Zǔ*;�6��f�K8Ql��v풮�r!N��r��6��4�F�w�����#�B��$���R�����(�PM��`��X/.����
�4�L[��E�X�<C�H�-gmGp=wS��XU,�YEfQje/�����~�η���W�G )��Xelʜn�ѓ�UW�M�� :���S9�{/n�A��I�tݜ&8��L�FJL@!t�����=)��)d���ɜ�� �N�T)�l'[�2^R�,���مS���Ӥ��Qf�%"tW�>T������6^"��%<���:MCj���aNI��-�b�����?�2O.^i�ęO�ua�����c����|3S�T���|�.���Ε
+ӄO�j@�Qy�\��<!9R��Y����e3�9g��x��K)�9B)s�c�[������u����p��	�yp=_'�)��ɇ��G@b6{jV��X!e�Rԉ��]��l�13��1��7S���69>���L1�����yr�Rtvp��x�K��{>ʙB&�F
�t�<����~�����)%V����,�q]����-g�'�3.6�!�%���ŞL��s�~�-��mj,Զ�GTH�	����3�R:�`�5\o�1��4��A��%|�x�u��&%4E\�jD`�Ü�ep�гmF����[�#R�2��MN�T��햱�����G�����%.���R"�#)	ΠX�@h��dQ�O�W� !���
��pa���Z����{ٳ�+�
�0�<��-"Ɇ�os��
y�h+�Bֆ�F��A����,�5n�8�&l���W,:�E�Y/zV+�4������w������5js��Y��@A07ӛ�j�W2�`�%��͟�v�w~�)m����XvkĿA����]��Ʉ�H�Wla:��7���:(#���j�r�����Ĳ�~�a��=c6�Ĳ�9��!����\��*HR2F<F�N.&�Ug/�RR��􏑒aΐ���R��e\3"��#������$�ٍJ��D�]��r�V ��x�;�Ԭ��p��!&�T�AM]�uW
�@9��T�j��PQBM��q_EEP@%��dTb��0��S��oʕ�*��ʂk�1h�1���j�c�U�>~R
�N����.Tvufzf�D	�+U^5���!vۿ=���j�Y������9��ʜ�.TQ�F��kEP.��X�c����-zJ���8m�\�Bu���ӎ�n�G��VՅs�H��<�p^]��a��%F�&�S�[
 u5wR����RE/�P�S=G�6'0�� �cn����6;	:G��� 3��!G�ёN���R;�?]'��?sz@}�J�<���Rr�i!;R���]vL��)A�TwI�Ql�mǮ^_'u�P�.-�U�(K��'�)�u����ߎ|:DJ������h),.����YO0�{J�t�������w?�#�@w3�kx��W��e���̤BRx�������u�$�u5o��p��(X)����~�v��L;J�4��6p�3�������ky��9s��.H49b@����]3u=w��}�f�#愪���D����L�pn+��1�&�o���*/S�zm
�͊7�L�E�i���#q�!�4���֌Ϧ�&+��Iꘆ�S�X���=gz�4
�̀�H\GB46�;R ����9��3:��IB?)�ThJ2e�Kųw�-�4m�O�"�zG[de(BX\��}�e��!�Ϊ�#,p�����&9�(|i�b���pZ�5p�����g���͑���H��g�3d�m��z��C�s��H�asw��g_�֯sռK�1�t-��E�2Ӭ`��b��Ȅ��[�d�)�bx��GD�Z��3Fi�Ii��uӲ�n�c��@4ϵ�r�eM�0���h�!U�����<�E(�c��y(5}'����i϶i(�D���K�빿����&E��kLMëAXJf�Z�n|�3sF���f���	��x{ F;����t�������pW;U�a)���0��0�ڮb	��p������*!h���DMs*��	,S����Q5��S�&w�g��D��1M1󢘝lvv=E�1�ef�~ Q�c1�!�~~����ˉ%@+5�K�;�1sQUא=��s��#4��sIh]F:ǐa�������c>~�熕r�4�b=�_�r�?k}�}�r(i)FN�]�SʄZ���ܼ)N��9մR�3��97ԟ�rf`��=8XG:h��c��q�[�L�j������g
��M����:s~��/��ةj�� �A��r|o�S5-13Ԝ���w�P��Ww�;ϔ���}/W=Y�M�T��1aL����yk\�%3�����%��L��O��KL�]�4�%�2UJy�ś�K\εL�<w�;�c+��n��Qʈ�P�
�nx9N�����W�2����    IDAT�)��q��*��G�D��!k�uB�	#�_�^��L�On�� ]��.����u�`e����$\�&>���h2�&���<ҩgMܓs�+�L�[��:q�>��K�9{)ܥ�o��2��M捅���V�Gae¢q$`?�:{��*���޳c��K�zC&v�g�L|�_q�lY��+_�;O�Wжl�����pyǓޱǅ��ղ�L���8>k:6ŸN�gS�6g$L�f�a�O���Q\�\2���j���H���
Ʉ���I>�^�5kw�[rE"ј�[&dΟ��_eS
W�x�`SJ�'�2R������鲰����]�I�ݾ�ɂSp�s^����j��by΢�ƏF7�r2H�EYB��tY[='�����n@r�c��Q�=6fB߰-�q�-�����o?�[,�(/�%�B��g�a�\�82N�F2a޿!R()��X1�LR%�sG���	�����oo�M�=�_2MB����ptl���ϑ'=qJ�fᙟ e`�I�;A}��͌6=�g��k� 6Y5p"�7�qG*; Z�D_�C,C)����h��L�\� �\�7*4V��u������PY�C�a��������Nf�Z�y�U���dRg�攩*���jv�����Df|��Q���lZXu��R��pm���,�����^�c�
(�u]���æ-;K�Y�?�p����*H�us'�\1�BN����R�P�f��r��+�lϹ�a�0�f��ۀ,��tRVd�|��+��v���p<�9��p �CT<���I�q����9&��P˪j�8�����y"豝��;��B�H|���ǩX�(�R��\�y�
3�\�� igE���+�|?a��Ɛ�g������;��~����K��`7�1�l��4���o��?�{������Hd��ifD�kwt,-��t�д���o2���C�X.�4m�k׻[6iK2�6��g�#��9_y�	Mp\]]r���]�nJ�)�	��,`x��:�eG��Ojޔ��%h�0lHe�\[��;�6w,�\�	|���|zY���&��Y�F�f��Ò��vSĹ��{Rّ���L��[��7�|�1M�y�1�����
}
�Z�n���g���4����V_��#i7R�5��5����W�|��p�����H��z^�#�@J����zu����bMC@]�^v�Y�,v?���G�-w�y�B�|mu�WC��%_�k�.,x��||}�g��^=��~�/�L'���i��e�\��f,�����Lnb��[������;�g�x7]�rT��*o�-n��L�ܼ�������y��CSFbU��s��ٿ��m���mu�qd���]\��qB�c���{>��y���7�|���C�_�ka���X.���Ƈ�u��������n�%O#nV_�q13���z]X�S�e��eЉaJ�����Վa��������g%ƹF�Y��ı3aߴ���v��BqE�)ML6bR0�ȟ�x�<?_�v��#��}J�N<y��}���VI���Ο�|y��}�k��|�`��D�L7W-7���;;U v6��ϟ�Z�r��nf{1���hqvT��ys���x�ڣ�%"�Ӊ����R��FƵ��������,���`w��i�jy�s����{�Ĝ)�!O��y�(S�spQ����%�P��(9%�k���F�<Pw��2Fe�x�8T��Y����$?�����x��i���pQZv��0��B.�r�w�R`!��D(�㞈&3�},�8���9������vl��	(kDz.��!3U%@���IP�?M�?8�_��W}�ó���j���͞X�Ϸ��{9N��a�h���|����t�4��F��X�Z���+�#3�\��s����z�������+,���l�;��x"��v�|�����[G�e��HD\�x�'��11i���z�V+.oF�8�Z-�+�С>�4�؟1F,dB�T2Ӹ������ʿ�?�?�!����17L���+�N�j>�BT+8�Y�K��E�����=9����VOx��5�y�C>��CBhx�K_b���L�[�#S���+�_��W������}�w#c�DfGl��Y�g�������4�s�������l�`s�g�߲Xtd��� M��dhi����7^���ow|0\m6진��VF�RKm���6��Y�Um�Sd��!��id3m�03v�@*�����Q��|I�n�Y_A�4�}͖ͫM1RӀkqA�nDfcEA�⻖,5�C�l�W$;�EOӵ�zu�vP����Kv��Yvąp�xB��,��;޿��2�"dW����s��W�M�#m�3;V����~u���]̌���jÇ�7���=����C�~?�x����n����l&&�;�S$Fb�5�ͼF������H��_ֲ.���\�ݲ�ݰ]�a&\��WCC/���1.n�wyy7p3D�$PG)��D�BˮR���i/֨w�]K�Z���~�	V`��>�b{w�X�Onw<])y��m[���ŉVg[���cN�`w��';��S�urrP�NL�ц��Ս���ˬHw���R���?��pN�6�D)��>���f��P��d)2ofS˫W}�L���Z˟sƒ�]���:1�"m��;b)�o6<�e��蜮�X.s��gr�aWO���f/���'�S͒��.HF��Zi�G8B!K���z(���b���bN�5*`c�z9ֈ(��J��V'����[(�Ò�#~�睢�Z�2�<1���� ��gG���G}�Q'���E�8M��5���Ŭ���Zt��Z�����;�`]8��I�2�p�뙾��
s�dV��πł�H��j��_�X�/q��_棗�X��6��l�����G?�17��.^�6a����Y�dI�B���;�j�������+���隔���(f�)�*4�'4Ӵ�~M�x�o~�!%~���}��g/�nk�9�'�T��T-W�l�Z�@����X-�<~�j������8;[�|����[6������?G���?�>�����a�!����͗�UU�\pt�#��J�JA��K�sL�O�W�SJ���QI���@p���?��������~�ۼ��p�۳-0��K�h�N�ֲ'U�q���n�j�̢	��/�q����`���e�_�H��hp������q$�W��_�2�O�|��w����U)�!P�-�z�jJ�iD����е<��ct��m_��O^]b��.Ϙ6;�\AۖwQ��g|�/��k����?���;S��PZ<u�,U�LPM��:�����b�fL#Y@�c3�2H�s��=FG�	q�rߴ��cݚKu���w�H�CաX5�N�PiԶ����m/��!�\���Eц���iV+\�f����8	ow-�o�Zŀ��\i�G7�܏#�@hjj�D��P#h�{�j%a�Ⱦc��_f�����Ħ[�|<f�����e2�z���#,c����,NT����!Ӝ1�ǁЌ"��A_t ��ח#x5����Y�C�k��sm����2�^���T)���P�%�Gfת�O���-�{$<�(�o�@{�Ô)�,/���I���T���5�b�64�rb5,+V�.�"B7�	(�� ����0�?��&�Y��Dg�Zͻ�o�C�RS9Z%W�/u#6���<8�i����A�W�� �O�w�G�i�h��_�pV�m^,��+�IUy�j�t���=�4?T�;	%~�^v�������>����|K�F돢o=h����V�㖴'�*G�8�/َO�� >Pa<l�\b��#�L<%à�ܮ��������k>��C����;\�ܰ
Kv:�I���:��(���O�i�q��B��«��lE�{.��q����a����;������i����7Y_<�����֏���/�߽�68�F>�Qp�2��5����׾F���xƛ_~��?���Պ���G�������x��^��j�|�=~��w�-��)��[Ɣ��t��1J�1G�Ο1l7�������[����W����p�ȢܺD�;�Ӏw�l�X��چ���������t�i��8�r�R `h|ӠZ�Ip��o�,%����g<{v��Y�ۜ�V+�67�)�G�)�}�H]��O�&.�s�g��_"��-�8FR�������qJ,���_�a�X�|u
���W+^�zE�-�E��J�[�e`'�8V��^���|��+>��ڎ����y�\jy��RU�J�Z�EeUV�m��O�-ȥ����'�XS��t�#�����I���������}��������!�4��	�k)N0M�?k���Yv��}N���'n��)� e�hɩ����%���v) 	� ���0�;3;��n<�?�{�{���T�SS���Nx���>!�ۆ�b1A�%uSBc���l^Pu[Qv-I��{O��J�|�:�|����I�X�zΓ�WT�$� �l��6�s��I���� �����9��`�d��ޞ#�(�-�i�W��l*�"�	H�EI����!��3҅�k/G|ގ��o��;N1b*����"mm�� �|�CD4Ds��8ki��Zӳk+�ᑺ�����	���L%�������R�-�ơ�:��m	�3�rO�������{�"�
g��#<�^'(I��r�8B�@�M�<
)b��
�u�h��5��xgB��S����\c�7R�:������6�C��f}�l���|_�է����T0&������^?Ɵ�C��1�|<��H��UT�}�{Xl��7x+Q�Km��\��$q��fh�p}8� *����f4�9��D�8~���@����4f��C����&>���d��-���=��O?���l����g�����͚mSK\(���(�l�l6CX��j�$�(
�y�]�ɟ�1W�5�y��w>`6�a]�q�/@�G�d��Qnj>��N<Bشh����g��/t0�T����QKE۵h�麆4�����i����GS[T�����?��@(�D�-;2�PZqv��=Y�"\ƽ�]�p�_�l,��g 
*OYn��9�ł��ɧ9��.�vK"G'��e>�SWN_='�@c)�E�eO�y�ݻp^�op2%O,릡u/$z(A�vl -i�ɋ�6�f3>|H�VEZr|'�]��b:����quv��`��C�3��W;��9�����	tM����S��f*��V�9�/YS��tXہ�d��������W���w��n:�>x����/��eY�|��WOp���ŁUL� Wo="	�;cmh3���{	�;��!�d���'Ֆ<S��!,�����='�򜮭� XW���L�G���k�C�i^��	M�O��Y���iQp�< ���1˦��%��.�����A��D�,�qƓ8ϋ6ᢙ�g
l�;�V%���=��%x}h�3���cڶf6��u p���]�)�w�T�@�4	ev�q(k���H(RZ�z`��ľH���Ԃ�/�P�u奊��X��l�2�p��dEDo�Z�a{���o����^�w8l0~���2�����u�d�)�ڕ�U�d� MvuM�r*�Ҩb
*�4W��xH�ڶ���|���hۖ��1S)�	���)P����J.��~O�1M־��:��	
��ӓ��#���s�cݟ�}+T
�a�ayp�"��-*������y�ȷ����̝_+_�_�C>��b��>-�[|X4�
2Z_�s��%F�{���>"�l\�ױ{�fT��?��V���:�7���u���{_��n���� �U�7�@	�tL�cc[���4a׬y}��/�>�C�"Is���I� �R�Ԥir�Z�uOg-iVp��}�i�|1%��U,�4M999a�m0]K��䓂�g�y�>'M5�Y���f�K桜S��#cF���O�f�u�j����1�[���X��U��'L.^��	Bv�-�^���?���g<�xŽ��`Rx^�zA�uHB6o|�怴H���b�r6'U���S�=�Ǐ�c�������ﲘ2?8d��	��+�ph�1��v���D�Ȕ$��sh�x����2pUkz6/�����9���?��ѵU0Ȗ=x��٧���������OxCSm�w��,4m�� ���i����KZ�Q�`8���dRTUE��p||L]�Ȳ�;w���C+x����^�(�Ie�i;���y��8��@J�|v�f��n[����
���F�N$���G�|�{�������3��=���he9}�r}��-�`$�<�V����彷�fw���l��U��^��ң�Г� ��t���L�����?�ږ4�`���e�����C����Sv����ˣ��η�Y���sLՑ,�Ts�=���ִ� �'I�p}�h�C
K��,�s&y���=l۲Z�X̹l��vK�k��&��1�%Rv�?��#LSr�ې(�Lt���{nOP6=9�^��!�!�/U 
d(���� 5z����>�A)z��y�	^�N�R����&Li��
�e苹���YJUUH�ɳV)��Q�R[�FO���wx�����a�+i�3)ft"Ȟ�nX������뚺�9T5g_>����!O/9R�B�$��ڄ���5��t-=8/{��h�8:�P�b��v �G\B�>]�]9�A�����*���ZD�X�~�k�����H��A�~`#��]W��{e"	q1��#��H&*�x��C�k
6>�p�ލ�i�&}��h���W}�h�J>\�+�D������P�)�;?��*\�?���G/���4Nk��©����C����dΫ�j[���L�X/i�Vo�����H��%$�/��]@Cg9�|A�ͨ�-y��������)�{d���C& U(�L��<��������ìH���ł4Mq�!�$�3�$a�d2�:�&!�&�EN6ɐ6E�P6-Ƈv�����6��n6��v�g>Iu@�v߈��_,Y����6�Ҿ9���`�����'��&MC�$�	D�鄶h�"L���O�[�M�?�0���	�+���>m�BW[cZ:�2��x�[�!%L��ɝ{d:�}�y�"�#��ڃ��-���S�~��Slۑ'�Ty�?z�L���a�t�bڀ>N�kU]sUW�����]6��r���Ϩ���|��K�#�RR]�y�V�Ֆ�N_���C(8I�݆�5�B	��rJ:t�W�I�1��'�dx��#�|?���F��4q��_�G�L&9Z&�"�k���5/����ՆDH�i)�kL]j�i��A�8�>��f(����w��w���̖3�'���[l�g��x��-]��F��r��P=x��dN�NI��W��ݮ�u�<Z~�NH��$�@�*C״�;ǴuM�u,��"LC�����C�ʩ�k::mq�bv��T�
_]�/^!���D����B_���5�{$�o��C�mpC����@��zY��U�H-�Dm��do`D>��`��5�u��ù=N�h*�]�P�De�$�q<oŃ�y�?�уw9�s���{�ON�Ӝ]�ruuEYU��e�YV�-�U贘�9������\s��]��P}����/�öb�{�O��'���I�7}��`�<3���ÚP�J,��|@{�o��������Q�n��Jv����׽����p��=c�����������i��2��3	/�蘣�9����_=��)��;�r��� �>&��8����DP�5/�/��}�z�S5��(��	3�C"-��KD�H'�ͨ��i�ٶ�f��w�ń�	�T(��6������"�3&�	�����i>!�6mMY�$	t�%�2�ے��fEhT1�Ni:A�ِ�х�Ϭ�a\ [ҢAx��fm��G-&�����T�&��3$Yʝ��8���ͮd�Z�u-�̱Vr8YR]lP��0/�.qۙ>��W� d`�JҔtRP�tU���%�������# .//�u��ߔ�錺�R��y�� �%I�v��uM���\m�h��&���M��K��-D�#����)i�Y,�x]��7LS�d:�ZK�۠�&���;'خa�l�v �@s��A�mUSi)��    IDAT����	�;ʦ��f迀V�:�:^I�~�������k��9��b6�ryy��lRк�@�͋/x��y6��0:	5�^�|��sf�@K�����sx�$K��	�9��;��]�e�I&�M�b����]g�+G�=O>��O>��`>��t-uW3���t5N8�D�UPB!ʖ�E������|�מ��#����d�sy>��� ���ѩ�KM��\o��o>d�N�X���pvuI!Z�0t`j��$Y�Jl�iMCY>!�s��	:My��x��������������$����j���R������͊;M�ۉ�Ӯq���Bg� ��k���O�����%�Mc��#�"V(�k-]��xk�#Zj�*p�ۇ��k��� �>4�F�J,E6a�m�U��;�������$w�q�{�O'L�S���/^�����/�mZ��sp��*C�!!��i��T��Ӕ�2���]f�哯����z7���P���p}�����t=��C���)�GE���_����0G�H����Bn�D&%R��QȆ�S~�Bˑ�s���@�BJdC`�J'cN�wأ���zo���t�=��`e`u�^ỰhT*Z����~i��x�+G����}�G�
X�O��uX�1'�F��W�2x"�h9X���ۛ�Bt4���95x��{��Q�����Z��H��5�z�;C���n�8
��x�3$�;FIO��J�i�{'C�VY�x��!�^�)H�b����PT�3��)�kY���Ԍ��D�V\���a}%C}��o�#I2v��o�hk-��=�XR+v��bF^TMK�$8�pԠ�u��&�]��ؕ+��lw%��"f�!�B�̦iȲg<���F�r�����I�Ѹ���C�d�:��M����3��Ϲ\W���6h��I��|��y�=.�}��t�]����Ӡ�
	*Ѥ>�XLX/�n�x%�YSd`�,ϸ�����#.��w3�\]]�$�8$�4�b���,�6`+�$�{*X��=(f���霮�m��,'��u��k�4����GW?G���,�P�J�$I���ٞo����D��Exo�A�T-�+������{�c�Za(H��1�t+Φ$B�f%xO]�zC.���2�´�iȵ��㲡�LP8�$˂+&9<`6]���;�ܽCZ,����#�MK.��∫��w�Sp���9+6|�[�mX��WH��
L��@)�$/��J�?|����8gX]�sr�?}�m9>)8�+2�`��=^Xr������Hu�Ʈ�N�YF�k&=���C�A���7䙿|��|k�]�N��� DY��(Wc�҅C��wv /%I�t�h$6�T�$�)t�ٵ[:�9u]1�Mظ���ۤ|��w����>��d1g.eY��/~�W_}��O�Q�%������|�H�~)��6������_J��dJ��ȴ���'��b�-��H�E����ȴ@���!�~�E��6.̍st��iI�Rh�2,��+��I�p��u􃻼��BG*:���Y��u����q�x9*'�Xr1Zo�|�Ml���{7�V��T�:���_Y��Wz�N�ka��5��r[Xh����U�2���׾w[T">��A�ct�m߹�}7@Vs�i�l͖ �� �"���J%T=��ZKS6���%uc����G4B�R)�����5��4O(�-^i�|2G+�v�e�Z��c��!�*�B}<.Q��0u �Zk��%��r�6k��2)
D-PiB�'t�Ex��)��4ϰF�fI�oj���W�hh���d���!i�ruuE�6ܽ{)�_���J����)��j-X�6쪚�d�v�BJM�u�����AJ�r����P6�mK�u�Z���,��J�*�	y�4�AK�x�~�L��	IֲݔT�s������a�^���@k=��g��t����n�֚gO�P7;<x�h� �H�u���@���VR6P\[߷��o�C��4��k^�z���n��H�ВX	2�;�T):-pe肨�C�.����\�\���{9�)��wam�`-���䰶�jvxip6�/9�^[�c%5Do��q�Q�K�I(�������3�D�f9���iC�ll	�e	McpƆ��I
B`[�i�N�}N~<}�r|�O>���f����-l?���Zf�%u��ؚ<�(/1�B�9�i��������`��?��&�{�˃C������׿�5����	RK�BIK���$:�������=����CZ/��r�z�e�Zqq����9m����G?���S֧gd�AIE��$��4��s��u*z���8��\O��:l���m1f/�Ǉ�80�ư|T���m,Ay����a�W?VB��\�{��D}ӤŅ=^Cn�o2�������Д����$���co������ߴ(��uK���h�?"TaS=�m�)�G�zr�2ѨD�mm5B'��;�|��gϞS�Y>^a^�"�c�eY���b2���
�rE��\�רD�t5W�,�����rM�d��Ek���p��sE>�<��b<��Q*l�J��a�XPU%��:x�^����M����Y�פɔ]Y�ٟw<�qB���d2!I�.�R�޽�5��,9<<FAӒ�J�ФIhN�/ٖ-:ͨ����@�yC���5|QɎ��9G�e,3��K��Ѷ-�X�]I>-�:�
^�:��tE�v���k!�o�	�ʾ�D|�i#4*����{��}�V���K����,s�7��8���;�(�KL�c��S:+��ӷ]o�^8�ł4I(7k�INgj� U�s���%�.4�ބ(e�^����a�0���@�v�r�~VeE��Ӷ�$�F��|��J�VgH	��2+�ɗ�)ʛ����̒R����������$I�-�Ȳ�������j��_!bU;� UB���5�ٜ�4G��̓r�b�A�EoC��9�!�nzHV�v����:�lɮ,1�R�9Meh[��3�(6������Dw�����#U	��������/^�Ѷ-y^����<|�6���c�^��'���÷��m����)����)B]_R�5w�~�ښ�披�3��N_<�$G-��+6g����,��x�`}�"��+W��:>�'T����hq]�ao��@z�A��p�冹e#�K�b�W �9o����?bӻV���w>�������m��vV���<��J�К�Xg��~��R~cQ��oT��Ɵ�&~ |7�7m���k�|��[������ѩ7oo��g���J�a�F�ŇҔHH�+��tJ�=W�@�+<ִC���i�Ri�R�-u��Y�t������HtF1���l����/^rqqH��3ᮿIH�4��l��sǉϟ�)O�<���+�<��Ζ�l�8|��c�,G�z�C�j|��5�s}�^��$	J����׬½Um��	'''�����Z1�Nq��dZa]�'�{�j�C�c�%����?(��>�1��7��.��tm�凶�]ױX,��a(���mI�*����ϸ����Ɖ)4m�޺R�u�Q��&���TeGW��͖�bA��Hf�yN�*�`:>{�5�MKQ�L4ee��vH���~�애��<�����ښ4M�s爦����8�X.q̺�Ͽ�j�B�s�w���y����PJ�[�M��g��{��-\.�LӜ1�:�I�f����+���f?��4VTC�T)1�bܾ�$G�iO��0G�R���f�������yG��n[q�ڠtJӵX�Wk�%�`:��Ť ъ���辩�E���1^[��J��E!��QZ��g�ɒP=���Sf?�!�I�w�=`}~ɿ���y��1Y�8�s���#��������l��2.OOy�?���{��Oz�iYoV�z���_~Ƌ/�K� P5k��$��|���;�y�}��w��:�z�%��Sj�~���i�K����LgC�\H�XbkL���F��}+�P�G ��aJ%���n��X�<���� �{��a!n��5��us!�����(����w}�߇�t`]�C�֑$����֒$�����`���`���oz���
�� ���?o[��H���a�po�g�{%��J�V/�J
ʺ��R<:b�xZ��I��,G)9xwQ�l�[:g�r�����9(�SR�X�w<}�����@���b�AH���֚��[�=�&rg���4a2�!t³��s~q�b���v��ū<}���uA���k���+����TTm۲��k��?>>��:~�˿e�Ysxx�Pppp���)����ڣ�N3�>k!�0b�pT����7o�c�۱Y��f�6%���$���e��&��K����ڐ
麖��0^W��?��YL[ �P��!w�a�4��X��=�3-���O�'�����_��%TuCey��4`��ƢX{Z�~���~�?��-�V�i����͊b:a�9G!8??��ӧ4�!����o�A���P�ؾW�^1�׃��tJ�c����$IC0��������E`�%�Y==�{Л��W�{�vlp�fiV DK'��m�n�cHӔ���������B�X��BZ3�
���IU��d�D[l�C��s��{�o���^��i�=���18F�us�{��_W��H���y2�n�����6˟���O~LcCc������_���xa�|�>:���~����(@(ʺ��\st�����n����|��ox��K��K6����
�-�m_�7-&�99b�\���?��'�{oQ�t>��4�<}B]�dҠ=h$�3��PڧY����>M�슰/I��!����,D��Hi�+�X���B��L��9����8�������X{N����?�s��b7�����t��,Kt��p���I�W4��K"��p��5����B)�Q(+$�|\7V������W���Y�{GP�} ��a�G���?�!�XZ!!Q(��}'��vKWWX��B�"����M*�$�1�d�u.Tmn6(��珹��������9��Xowl�6xQt=��g���8<Ǣ陯�в�碬��^Q�&'��Ϟ���SV�U�'�/������)I��ޔt]�tޏ��cAs�㴅�A8G�@�4H-C."�-.W\^^R�J?~�ג��N_������=ۘ��r���r�.�`�4M@�������*���Y޿���+�<�2�l��
���ׯI�9�P	ɵ0�s��q�p�N)�0�i�Z&�	ƴ�m��rNUU|���c�Q������|��K��!�m��)y6�n�ў�ݨ��t�ǚ������>M�����Mɝ;G(���ً��:=G��B�w��hO���8��3>�͈BY�Czc>����K�Ԝa:�����XoJZ#q^^��zsƀ�q�'�r������rN_<�5�ɬd;����|�ٗ����l�y�h�+��-i;ѡ��v5�u ���!b��H
�䳿�J2�n�!��i�b���O�9����/�5s�z�]>�����_��L(|���;�������er��	eݰޖdY��`�s�������o��7|���֒Ȍ�1x���%[W�T�`('I��W���3^~������wO��g�,��WO�2��Ȥ"���@��ߣ5iM�%��뛣��E�v�#5,{����[��q�pC������h�����M��)�h�TA��E鬠�#Kd<�4�88:�����Fts�����FA�}z��.Q����(��.Ⱦ)�p��x�{���g?t��i��ۓ0�s}pH�
�Q:��z��1�+��iB��:��8�sHc,����:�`�]n(�הe��AA��!<mW��� �����1{�7��9G��U�4�y���d�	�mM�R�9�]�/[��A��r:�ݘ�q�f�>*X��L�4��oۖ?��]��v��zM��0��ij�z��9JҬ�v-YV\{��8���`�D�U!eYrp��z��g?�mېjI�%X#�-ʦb[ux�A�-�s�ТaS��p��!� �B)eT<Q�V�$ih=��9O�<a��QS��wLK����mMәO�(���?���� ʚ�w�T�s���{t�as��nJ��p�<(��>~̫׫�i|h�26��#���8>^7�Vc4�����9=}��`���EH��_���+�^�lt*�+�qz,^w���6��!���,�K�;������d�zuI�%�W+>���Ӂ�K�6��C�*d�P��L��\
dۑ�X���:���`o��m�Λ�������D��\77uEW�O���E>�����O�9��c���;��o~��_|E���d���?����O�J���)/_�2_p��!˧����7����?c��ѵAB��(����H�����/m�:�,�P��ٓ����`����9|��L�3.�S̗�`�5�������7�ҍ"��2�7���A�}���z�H���=C[�azJ�'��Ľ�4��9~��C>�W"�ҵ6tI�iB[wԭ�[K!�7��a��с���m����D����^<Ͼ�Ի�E��i�k�9lp��H�{V�}���t0����
3��]��A@7>�I���xi�S��1���B�E�e<z�)9>>��$�������	Ϟ��9G�44ME���7��^Ր7�v�蜣m[�R,�,3�$�1����szq�)K�Nؖ;��X[S�%ǇGׄ'p�{�׉G4r�,�m�AQh�)��d�w4��j�u\�%��:QiG��M�d�h�=ݽ(uOOO���T�"G��_��%<m[3)1_�Z]�^wL���PW-Y:}C�h���jx��aLH�x���M�:(^C���Ǐy��9R�ʎb1�Ν>}��]MH�4(eH��g߼=?V�q�\wRN�&9��/�ׁ���;�L�K�%�[��q6��t�MoYa-��<q.i��B������>��l�Q7�pq^�?��U;������mF�M�?�����2�W�|�R
�<��Z���]my��5i�Q�QZ��L��鐲�Lf$Bb�ٶpZ{|Э��x��P����o� -l�Q 5����mNێˋ׼�,��_���_|�-2�D��?���ɏ�+�MC>-��z�'�~ʣGo���..^�˟������٬��ݔ�+��(�@n䤃��ˎIqL�T�U�5�2��Z�Ʋ^�9H
l)Ț!����޺��o��l����l��ė%��C���y�~���g_�'à��Mc�m�[�ֹѠƓ9�:�_����/�и��&����gJ�{B���'�Z�� f�4T���Q����{0�q$B�J˫'����s5�Ѩ��'9.
����!�C�@�r���o��"���$��u�q}�J��9I�R�~�q��s�������6��H��<��zsk-�N��3�Ɠ����(���dy���(hՄ��`6?�3�j(1>p�+��U��b���ۏ?C���!�%�o�"MS>�������>�R�-IR����`��*��l>��R��Tu�c�I�^��"���<I���&�IXo�v��6��G���,��c�Zs��	����f3ڦi��tb���Ѱe6�����劷>����g�X L������gϞ�g�ބ���z,Qy�OpTJ���!��Q�Ʉ�n9>>������/�2t�+�*�:%M<]`t	�.�Z����7��n�2��XĔFܛ���$�?�)'''|��G�e�NUU�W;>��	����r�P:�m�����X�GC">����]�v�P�v����/._����{wO�l>���j�h��D�&�΃�#(���C��[�����0e�%MS~�7�'(����ٜ�n���0��1v�s�T�ȡ1Bߋ���&^���i��ϴ��bz0�����m,]�0��Lg�ْ���૗��Z��j��:����J����;���t��d�i{�=:2�����M�&��6�~����C�ػѹz9��2���M�̩�N
i�ڢc���,�����QO�]~�F�˗kʋ�dAUV�7�~���-�i��2�ӿ�w���;<�w��������Ƨ���y1%�g�X�Q7�3}�Z"����'    IDAT�5uհ�O��MӔ�t>TedYƅ�QVS[S���l���9�i��O�����RlZt��IO�:�W����H��@xM-=��v£�:rCS���O�>$�F��C
>�V��wmBś���<��,؛yCF����+θq�go��6����"��6����w~E}Y������{��,-�7S�0���o��o�}��m����xR�SVkÎ��%	^@�6̲�<�N_pVK��+�T�hI]^w���K������<�͆�
��� �ggg}��&+r��a���4��0�^(�8<<��p>B-MS����8l0Tϟ?��t{��1����l���HDT�u]�eِk�׉ ���#2�{?({!IB�WWW|��G�5���i���Z����{�yo��5�"��N1�/�{��TU�j���}������H\�1j�6q~�e���U)%�x��p�������1���������#e��S7��=�ۼ���hL��>J#BAyn�k.//+�%�3�>��%i��]�f�(�M�!w3��g>�\�Z��4�����f�n�{�<8���7J<�H~Ƶ2�8/RJ��{@Um��S7�.4�r;϶ڲYW��_P�u��v��,�0HgCٱ�L�b�r� mh�u[Z�c��ߧ�ǟ�&����õ4���� }��.��s������?�}��OY.ζ�a��_��?���'�]�Fx�RͿ�?�W�K~���_|�_��_p���I>���j�eW��k���\{�{"tl�C�Ά4c��ߝs�_�RR�:�bۆ��=��9��|��jK��SvMKB�o�Ь-b�`������c �yݢ�mBƊ�^��$��J�nN��>�mo	k�?��؉}��������I��Fl��O���8<>����/ٽ>6����aD���K���Q ��׼1>��[7�M���Fc���<��I������n�$=�C{�R�7��zAWbL�N�s+A�Q�o9A����Z�d����WWW(�r����l�e��4�	X (e�U���d�r���?��ٶ-�_��I� ���jW�t�^�s�Eq��i��b^<F"�&*�(�gj> 䪪�ZK�����4�?�����gL�2Εg�!����Z��là�:������E��>X���N�Ьh��_�' T<{���o�o�����n�DLM3\�O�x��e�k7����M"��muR)�A����C)J�J�{����ơ��5���mȑ�/�͊�� ��ȪT�e�n0�@Ƹ������|�qzj�������
�H�4�զY��)BZ�z��V�MO��h;�����6�YƝ�	-)a,Bݼ���v|/���m�o:��8>�?$5��Լ�a@S_Iԏ�b���񺳼���8&����	������gXk�M�������_�'?�g|�����/�ӯ�pttD�����$@���j\?�RF��= �i�aM9�����u���U/c���t�}����Zq�B��5�}g ҲҲ��zC��~�)��D	����ȋ���>I��;�/o���������>Ї�����㚸}Q�`Y׊�NBd���uf�_Ӽ�R~�5fS�OB'��֜s��5,�pS����h��a��k�{E��[�9~��&�A���c�b[��j��(�i�dF�*��+��5S�I�	Y��	�����|�z���*T:�J��>�u�N��%z�Y�R�u��d �^�X��i:��CX<zӑ�%	I���{��E�ړ���C�]�rttD��e9�����<td3k�������j5䨣A��B�$I�9�P5]���wY�C��@��t��VJ�Y3TD�����0�4tߊ�^�6`/��4�w�=�����7㪀��8??���<<{opYk)�r����\���9Vf�~��̧��Uy4��vm]���Ȩt�A���~�7��Z�ӛ�9�S[�ڊ�j�:�X���n�g�"���,z1euӈ�׎�<6�ocW�-�I����+�CU�BԪ�B���j���X��Α
��bƝٔdS�%B�i`������f|�����͏Π�e�V�%V@�%;�3{��|��gte˪ڐs
R���.�v���k�z�?����7��}��z��?��˫i����)���t2�|�B%)]/[�Q�-I2b��#wB�A6�gPJ!<�c�h�r[qz��
M>�1���ts�k�z����ZۋPj޷r	X�K����]Կ���s��c�nv�	]���8��q8EPH!~���[6�m���c|.!D�g>Z<�bmMG!2_��?�eY3�r�1�����%e���l7�x�X	�Ƒ�m��ߴ�o*��c3�h��}���� ����^�3�4A%)�4�65]�q���n�v�Y>eW7�uM",Z*��"p-3�Х���,�ȲP��4�3�3zԃb�6�"�i(��=g)%H)Y]^���g�
�I����⌬mcd��Y��/�b�{O�S=z�v�9��2f��M8�y�����B�P��͈m+c~5z�!_~ݣ�i#�`|�譏�l�A���W � @!yT���׎�5��g���8�Ҷ�ڜv��,�ks�cLK^O篝��߮��l���,�hOS�O��G�ϱ�q{��Hb|}_��;ʃ8�1������q��8���UD돯?>Ɔ�e��ؖW4M�u32��Ɣ�ؚ�����R	Z��I����c��	w��6��K)���r��vO��}F��۔�X.��}dS*H�	��v�K�鄗/_�~��I�S��b>a��qw~��?���t��O?�W��3ں�b��'O��c�<D��:ö*YoK����sre�Z��-?��RJ��D���.>�A��]I����qw�s�����nKf,�S4��Bd���8GT�7����FD?j����1Pqq
�{�¿9yߠ�o
W�}o��[�x�A����5��c�4��{�ޓ �,碮�����$�f�mO�2z^����2v��H��G�{�w'�}���9n���p��=z|ȯ�~��b<޲%��I����y� QW�u��X,x}qΦ44�%�y�Y�� �y�}�v���y��{��̧�� pΑ�I���,�R��=�л^yF�7�LJ)doLD�޶m�L&ܹs�5_|�ŠP�e�l6���fP��<��~:3�c�P����WQ���cx�4�*�`�{�p{>)����>TH����rI�e���s.//)�|����iL����c�>�߱�=�$Q�؏SPt)���h
9�}U�1f�fn�ι�0����G%�Tk�PS?>�@ڵ�����·��7��so-�i�?���G�����6M��א��rfZ, �B��$H��iA����b5��!�׶����4��É�̪�搢���J���ל��p����'�n��))9=���Ǒ�i�q���=��]���NJ�	I:������BpD%�B�d��j��T�""�ho�l���O��~��S�Z?�& "�'b�~��=�Wt"����r��o����?������b�:�:%ܛ͆�o߱3������l�⫯������麞�X�QB�:�~�`]H��P��ǂ�?	��x�N85���H`�BI�s��=��ԑk��g��
qyA��E�)g�ϟ�� R���\8~�����^9���>MFH�I��sU���rz�؂�O��3v�xz����.��IEo��E�?�BI}DI{�A
T8?<��'ս�w�����.��3�8��N�š��� �v��r���y��7���'�z��@-��Cn>���]'i��������$Q$��0(��?m�N]�����r��ЬV+�<������;���i��������Ls���9;;�,�V�/����}��ݎ�,g��,˒vz�Zh���|���O�B O�d��X��D���2�-�!���D���e
�;li�9??g�^S�<^�l6s����2���&O��4Z��)`N#�� v�۶�g��9��x�IϠ:u܏�c��>8V������'���쉥��j'�5�o��#����~N�}z~O�����CJ�Ji��G)���DfJT�E�����ӱ����#�%!s����% P"K�*>�Nʴ?��	\���1�!ɔ��يZD����;�$���\a?�����a�s���:��6S$a��ǊU-	�W���|C\��O.ɫ��=P�9w��jA�l>\s�����Wx�怖��"]70���ȳ�Ff�s�x���al�O�ǎ�<���Y�!�$�C�3��*(�<#\��m�ɭ�OE��5�����>�G���.�SpΧ'�43��Fi�Og9/�i.~�}��ӯ������IH���O�2� -ND����N���i�t�J��1��lN@�'mT��rj_��|l�J��e�<I��L�A���Xq9�ϟ�K��������FG=���mo(�b���˳'�C����CL��JeB�c(�rnU+m��ir:+>^?ɸ���
!UU�Զ�������f3���*h
���v�9E�O��aX��<{��?���<ۗRryy�֚�m��,�����t�y۽
k|eYf�S�����xf߀�(8;;�C�4I�vt���|6.)˒��+B�}�v?�u��xF��$L�z�	O��{�p8$)�,c�\Ο����du���S��t��e9�pֱ�=���=��������fc�u$:�1�;��c����ܻ<Ð��)��D;~L������&r�5w�z������̿}�Gw�1����9�<<���	�W��R��i�"Q*��X���k�z;vf�Q��D 
��<�Y��mǰ� �C��6(�i����}0��}.�>�����-�O�H5��2X�S\=����{�v@>��I��\�k�O>w���M�_�P�P�����"/�!&��O��}s 
1V��Z����Zqڵ9Ţc��Ѵ-F)ʼ��r�������B@T��q�Ŀ�E����0�B�/<�ҟ�D�(�.y��7� SM�D����0�͈_@��G���AH5��Y\؍��N�c��kQ�̇� �C����jVIt����= u�ҋ�MA�t�!2�Y������m���ْ�v��H9rpǌ#�OZ�5ӗ�C*1���sŒ��O��B����w�)���p<yR�8
\D'p�E�/#�������>82k񡠍e�H��Z����R4&'�U�0;V*6�w�pݐ��Mv���B�>�� <�M���b��2��s����|�xA�7�ts�dF�VB�+T��n���
1
����Ȃ`]L����g<{��~x�ᚦiX�5�h���D�c��}ǳ/^�5o߾E�����%|�Lɮ��I�ZK�=�Cݦ�r�N�☌X���)���P�k�ՒLk��#���|ɛ��|��!-�"+	.���︾�]i�Jg� �ЃLꖹ��p�d-�����_���9ϟ?G*��(]˻����|D�t��,%��"[��*&F!R�&XO��d��-��[w!�u2�Ȥ��{��g,�˲���3�6�}��f���k�s��ۤO��4�Q#�"����2��~�)8��mRd�(�(P���§����������v�n�c3bL\H]m�s��8��֦5P&�D�@ʱ�vH�[m$���Ƨ���-en8;;�m[v��ܽ�B���j���~�΍˄��%"Q���8���"d$Sc4��x��~|��-Y��`��`ً	��D� �`�Xp��>M���N���d��j���t0��>���������_�������nC����k���^����P���ʒ����D	~��=e!qR���ap���;;
$�
t�ت]�}.Ǝ �o��x�D&�*PAPfi,�<�(�>u���H�y�n�˧
��t�:�Q@���X�%B�q��'n��+b�H�p� =�O+����)�\���S��Կ�T�Զ���㛥�+�?D9��� S�<΃���q��O��s���O/:fD�0���ܛE�V��ߝ���+�=l=O��p^��o�[�kECڐa�[���8�K��[����I�%��G�\��-�������  7FiD��3�$���B����d:#��*���Y����E�gS�����7��6x��TFq�S��\TX�ڢ��$y�R}����|���x�C����?p8�,�
��*��s���l�bU��������Ȋ��(fd5��W��
���������*LQ^s���H�T���V�(J���2/(2�s�7#��1�O.��mn�mE1V�	ў,E�X��u{"����.��n�Q@�ԋ����⼣\ԔՂ]������ ��a+\]=Ee%�M�,J��}@���ZCH=�ΈD���F#$)��HI|�!r�ӫ��ENf��s�CGP����Ue�}���O�KY�c����Z2�aE���N�j�ҽ��#f�L^�"~��֜]�s����_~Ż7o9�Ͽ��?~�>|@II>2(��y���B%Q=� �N���R+5�%H�˳5����ȹ8;�*�ѧa�1��_���")�B��(�L��H���Ǝmx�D	�Y�����u����	~@�i��"�[O�>��$�*�ϵ���܂�cҦ�$pgQd�E���G���Z̬DgHm��;Umw`�Y� �>&���Iϧj���v�2��CO�E82Z&|��7
%eB�>0�r���Ӹ!�ɜ�����(�]�����0�P�-Sw�4.?�0:����c��^��[�1��\nQ�Vq�Q���g�T�z�s)���z��"�}���N�瞟�J��oy_���Dfb)���U=�����=���{�~����
�z���URE���V�/���3�^� �'_�(]P�%w�->���n�<��O�;��x!0J�E}�>3e��E�9Y���)�B��Լ�<�������-��#O�gp|����Z$��I�|��е�Li
c�#=�ﱶ#��;g�%_����;����s�EN�$�9��#y�Q��[��з�0F�� �4]��5�1�RR�ת�9�-����R%��;Ye���������?"���n���X�ov��|Hݧ Z�0
��e��zEQ�l,1b�8���RbU��X�Q�%���<��ޠ���+$����Î��߲\�d�5��1Z�(xb��i�+�Qo[�#�_(9�� �$�)�A�D�ʪ�þ'S�e��v˷�~˾9��7ߠ�} �d�#���k�X�����1x7�W%"J��'Ø�Č0BS��%�w����3^VW�Z�.U��\��k��<�������j�G����Q2� R�A����X��<�zB���i�V�WWW����{g��"79�w��Î�*zB�۱�	nD��Hԉso��2������A�� V�{��c���n����1E�I��wAҁoۖ�^��9Ǣ�0#Pu�����A�H�z�=��P�����'vO ���[ i��u}L�8�N�&"͍�'����@��J�u6w�87��(���,�,��X2��$��	#%B&n��ux�R$�^Ge<<^���ؖ.�4/�G�" ��a�� ��d��g^<i>���M���3����tf��o��q���:·� ����8���cro�ı������{�8F"�Tm��,)��u�U�ruAY��E@U��9��!D��rB\��$ӆ��3���wI�.�ԺtCZ8���cۮ4�n��6Q'ѝuQ����o(T����|���l\J���x��!�Ty���/Q���x��g��-�fCUi��1��PXk�<���
޾~C����T������ժ��n����kt^!��h��<��b��$a�麎��6�I�Bf�\�##���lt�27,W%O��s��)���|�曯�b�7�v�m;v���kr�@�z�����v��nK;�/�<��ɓTኔ�<�<C�n�|؋"��E���g��5m߰��I�    IDAT�����"����]_�t��з�ဪ\�#W$âv�2b@��G�!xB𩲕*%��2�0 ��(��>�Ň��Z����?���i���-FJ��� ;@Ŀ#�'�<����".M �<7�9�%�ԉH���19W Q(#a eF���n7�=}�n�u�*K�5"˲J�S?P�@��;Bp�{����G��Z� ��� �,߬��oZ��-��~�d���n��m93XS�zg"�����0%�$4��Y��L��n@*IY֔�s�I�*A�%:�ġ'2Ȉ��FS�X���5�sk�õ�a���T��Z��=���o�b�Iv�(IQ%
�)��,+�q����jƮ�l2�
�0&Æ�@��Gz�z���2��Z�M���5�<i��`�$i�:�ps˅�uЊ�6�(�! pb~4�)p�;�����[�'�RL�lSz0�8�uR�z�ql�ρm���)(M�����z��'> 9����4��>6�wN3���?�R��Q�����+�O*������|E����kF���O,BL��Pd���j������/��/߲m�ed��jw��4�OT0)"��$�
.�I�97"K�=�㈴�3���������j������ih��������b����O(V޽yG����ޡ�d��yzy��YX���Ԋ�j��26�_|�����Bt��۷o8����;�0��"+T�'���+l����8g�H��m��̫�
�znnn�1Τs^UUzm�勗_��_S�m�#��~�r�p�YX�H���@�-gϞ���T�)%ϟ?e�^�;���{2-9[-X�u���[�11��z�.5�'�J7t��E�Q�o(�v���2��-W��|���?��SJv���.%y
��vO��M��T��(�)$�;��Ebj�y�����/xry��W����&U�.�td���W/������#.x2��YǄ�ȵA	������tm��ȄH�S�sBHP2����'���7-*
��[��xo����_%�����s��se���Q��`�/�Q�����a��4�_y�㇁�d��5/�>��rv�-�.�L��ȍ�|��סd����HqTn�F��6N��.M�W��0e��kYM㌁A��#� ���R|��yZ(���s]ؿ�3�ׇ�2�C<�ӭ�~�sꢌk�#�Y�7�v����wdy�$���Be�3cib�L�}3*K�fѤ8ƩS��I�I�#fz|g�3�)(�"��c܈�
�Bc��NZ�	�e<�(�8Ƙ��YV+���3�1��m��럔�� iG���1�	�k:���I}�����X�>�Z��Q
��^(����a���Av:I�]��'$�Hm�f/bő��R�?IV��}8�ꐜ~��{�������Kp-j����H3#7�3SP��=ϖ+�����[l�,//��P׆X�x�8��o����e�(;z��Gn{��p O//x���;v��g�y�R)����=����%������|���N2�Y��d���Cjwe�Y�'%e]�4�e��nOp���xv�@7���+����;�ίpC���ʄv�򫯸|�"��ƛ����,�ā�h�1R"F�	�wqqA���;���o_�4˲�IY���6?���|O�\s�Af��K7�z����3����n�qK�w3-Oˤ=`���b�1�E=K	!X����d{�'��/�'�!^����f�q�#��|$*�bU�����ï���w�azq΁M�kY&���H�������:���;����jVB��Wk�����k�4*,pqq����y��W繺�$�i뎦.��i��޿e�l��(�
�>
ھ�Ϣ�)��6�E]���s�a�w��{�CG��9Ϣ���7�P������,�
��d!��m�F#��YiY����B$fJ�kv�6xV˒�o�+2���ež>0����Z���?Φ8��TKp}�p�*Ό��Agj�
��:r�y��	O�>I�~��ȝe���D�V$ oL>�����Ed�<�����O[b�$=��L�vhx��-n���X�,��6�Q�J)���%?-�$
I���H阺����Ԏ�v��J�1<����FY�<���0mi�O�E��`ι�z��f3��i�t�S�ѡtԊ��ia�tk!g�)F��n����ݯ$9y���%ʓ��H;��J*�h��v��~I7zJ���x���X`�S����~����q 1ƣ�z(yXL�idq���'A�s�{��|��}�w����Bd<�#���73��[?`�E��p�~`0P�_B�Lv�mG׶�� 7�$Z��L��L2�������ݛ������ω��_�@�yυ
8;`t�e�)�{����&������j�eM�\pyy�:D�]C�Xt�Q�5e]%�5�ڶ�r͡�����.�`��c��������R�
�{��X�+��-W�s}�a�^S/�Lݯ</��Ͼe��RU9��z��EQ�㝯O�HE����6��#�7?Q�^���7x2a�MNq~���Sz�J���_����{=i$<C]�X�=�n'+�m�p�Xs�ZST%�U��yˇw���^�\��6A�Ed����%��+��>�n�*�ɓg<���_~�:8����ٷ�u�^�)�rxϻ#��HYs��j�ex���w��޼��H���.����_���Eśwo����<1t�sc���ٳ�o��z�$͡'FA?���$׊JI���^������QV�Ҵ{P�����_s��)?��EQ�o~�b����4͑G-R�?I�GӤ��z���N���p��*~��߲�n���G6��g���%Jg\>�BJ���7�gg<{�$����]�ь��j�b�\�FMӬxU���+���ӧ\\��ز����z�Fk&���I�7�|���T�=�r�u�_��O��QR��Fѣ�d�>o�\�v�0i���z�&:�P�;%��US�ͺ#�&�>3졪��z�����u0�<���~�<
fCZ��e?���J�&��j���b����<�[OZ����OO':;B���d&Қ�?or�+��n����k!=�����^P�2�������X,�jֻ���R�cc��Iʣ3�������ɩz����G�:6Y)�Y���L�{z�'W��8�i7��st�\2���XNя�$km�
��bbH��1���q~~�y�$6-?����޼�28�`�C��z�y�B�KI�3�b�`A��sr}}���ٚfբ��:����@���E�T5��c������޿���/�5[1к��2�U�*�j��EQ��%���r����^���O�<��ũ6�1�K��`ɂ��yǫo������*D���%EV|dQ/8;?����o�������ʲDZx��a08�ɲ|v�+�+L�t��������O�?|�%0���9�,��d�S��Q�����/.@H^�z�0)iv��D��0x8�\�H�0eF@q��⃥4
�5o^��=��{�p,��8	�,0��&7�i�ϟP�lO����#�K���h�~Ƅ,�+B�#�9GɌap�Fh�"���w~����{����xvqΝ���bU��_Jq��)�V�=-�E;+���B��K�H�=�f���O����~{�`;2�����_����������~��@*�)rno�o z�?ί�k�|�x�I�@k���;�L���咾��$OJ��I~9%$z\�_��W�ݿ������{���r)~������&�G�@!Fa�������l����]�G��8� LB�Ǐ����@����B��<�!��1G��S��)��c ��}SAx�2�W�D�̔���Oz!$����1j��d��t=�h��y�Zb�Z��.nR�9n� �f0޴io2���@�����1��] ��y�>�n"9ʿ�(r!���=�d��@H}O���7Y�=��ߓ���4��w^@g�	�B�T��(�BM�c0Si��l$��w;�PR����n^G�H)t�}� |!�i�y�ƘQp�xbF�I�>E��.�OզG%�1$Џ�C�08jY���#��CE���s~���/\��=�~x:�~K�O��u7˺J���a�'x�B B$���LK$����n���l�4" c�}�\�# ��nߧ����țw�X�V:�����'Ijr���h�0@�(c�U�:�v{��f�p������D�8�:7�h��w�Wĥ��f��h�pm��M�P�e��#�/�>��緔�ݡ��%���\���w��l凞���]T#�1C�Y^�B�����	�7\��Ø42����0J MF4���G��eF�٧žu��F�=û-ݫWd��Ry��MVB�)��˺`U�4���~�P��b���}� D$x�r�B/+�N�.�I���Ŕ���IMyVSE����c�������.����T�fY,h������%��բ��r��z��Ő�v�&��#Y��H������e�Ѡ�C�;��翧{���]�k�+�}Ca���_�Ǜ-NJ�q��	eY��Ke�ú�_�G�I�iD��~ٶ=]�PJcjC�"��5K�����?������`��g\>Y��w�,oO����K�4%�v\^^"Cd�%N�p-eA_*��Fd���]�&�H��z�����-f�q���z�տ���O����f˹
mK��y���.�EDͤ�	�&c�	��4Dy�C0�_�]�8��u�m
BTD
\�z��F���]
�X5���H�s�vkq����$Z�f�|��J��J�R5*��O
z
���	Kd`8@�c�/P2'�%�.l�B*��8���P�(}�tY�aSI�iB�G'�!
�PG	\9�Tg��� =��F�G��8���������L������L��ᨵ=��O]H����c	59��S�ϩ��)�����?�M��Y�rB�q|�T��<Ip�/I�	�4�9���o)A8Fĳ<B�D9�\��2��|��7<��oEI�Vt!��n�l3ue�>e�Z���b$�#�	@i���(!��}�[T�(�~ ����*Bi腤�
'E""���a=&+'ZgĶ�	�.�U��O���~�Ѓ0+�s�
%Z+�"��M������r���cK0F?zzK�.���ؠ6}�m52BH�!8Ę0˳����w,��L��.OV�=�W�m���5r�γ���U�r�@E�W��48��n6����'gxgi6w�-n�qEN^�dv,E�	*c��s�Z^����O��ف2�i����Mߡ�$�9��	�t�88ǻ�{}���!e4·$��<C�z�^*J�!n>p��`�z����ۄ�X�hchE��9����{�X�q��v�bn?�[�=����}���������l��ʜJ�b��D?ܱyw T���*�ȃ�>PfyZ�"/R�NW�uD�~��R�+	�;�?~�v���Z��P�M�A�v���x���{��s�4�egm*�LF��m۱�5�p�q��YGPՃ��̐Z�h�6|K��p��>�r�#���"�1H܀9�P�5.rR�?5>����/uh�����A�|FDj��
�:+(u���u�CQ�8g�CwoߥL3y8j�8g���ּ|�_}�BX޼~���5�����*tÀ̊�}YV�eYf�d��<�����R�d�!��F�n��x\�>��\-z�"nc�{�ܜT�S�KU:����� ���c��'�q��1 �����N_{�B�o�c�������E��epq��N���?��L�tOM+�����R�h���(�9X�V�
M�  �zfs<MI�C$��x&�U�NZ����(ȍ���9p�I�Vl)	y�I�.JE5x�j���(?L�=vi��QL�E!e�@
2����Q� 	����<����I���Gl�!�;�,Ǚ�dZ����D�8+M9?�?р���%}�f����M�/P"�o���Gf9�u�S�d	��ԩ#��d�	����>I��1:����>$��R�];�'�"����w� -F*D�ئ���?X`�/������=`�.%>���g+@��){nH��0 �L�4��k2TY����ha�xv��129������->�\c%Fns��H��M��)��kJ%p���-Jex�#��r�jEP��}��05qta;�mO^f��ι$�;XLYQ��X,dJ��;��+��Ƿ=��ےg+4���i�޾%�{��s��`��e��|C?�L�{!�I؈I��A���1�Dl�}JB��)�ŷ��jQ ���J"H��|}u�~�s��{~�����T���*	$�f״h��)M��0�N�:�8{<���t��@��O�(�5}�ɧ^���PH�,
�В�O���YE����SA��݄�(�pD��Y�����N��aF���x:L���K<Iv_^^���6��<}v�bYqssû��]�$�6�0&9�$|�"+���_�����-M�p��~������W*@����O����Dd��������#'Ú��>�{""���I�Q���F0���|����\?3���cB�Rg��8'ѱGj��}���R�s�AN��.�����n���T��w;&���4H$J�Ols���KJZ�}#ƈ�728S!�8�(��\h�����w���ӧ\>�;���[��
ʺBGE�m�a�$Jy3�qdڻ�>�T9/�]��7=Uf�lr��c�l�BV%:ϰB��DgѡG7� H�NҠ�Y& T�$�v�
ee���J�� )�Ż��ɤ8�H�Z���bH��A;�tj7g#Z��Ĥ�d:�;-8��C(9���vD:?	���*%��'�a?��]���a 1F!�D�>\
^1K�5�#qp�h|�(����ua�T���Nx�Dy^�l�IH*b�
;*�%ݟHt��e$�\�GhŪ^��O��b��n��-e�@�K���:I`�n��%#��q.)�V'�#C�.KL��G�2��{޾zGw��H�Pg��H�$�|���J%^�H�͝�lX�%a8�D���!�Hbp�C�Qf��k�����^R�lc�4�sm�x����q8�c|�5�<�w=28��a�#[_�:���#�:�?[����(ߣ��`[D�	>�i[ľI�����`B���21��wtCK��2X�@eJ��:������8�ܐp�|H�c<���2x�~>D>�>�p�\����}P�Lq��HP�h��@� �'�[�PdB�뾐z�)4Bl��s1��I]Zk-�޽#2���R�u��~��-}{���JM�7I��;��EA��,�4x��-�zn�����.�ĭ��T�ਥ��0��3��~}߈�Է$Iת �Z�zq�_9�'xz�sw��	�@M �����CO�4N?���x�&���gH�Н�L�J��&�od�D��L�^�B��	�%"���6�+�S�jq�>N؉�=��!�y)%(K�I�L(�!ۆ7�����p�����kZ��Y,�i�v���g��ClAILV���A��SK3+R���)F�,ݡ�kZ����)@ .&\E�,�Li�32V�I�_�8��W��>[�^�1H���[�߿N"0W/8��`}~�P������i/�i�BQ�Q3FT�	�"��}��s�0���:�6��o����7 �&���B��J9����Y���,G ����� ��F����J���D�@h�}�� e$��ɲ^�EƦ 慤��G�i)�2��]��ݎ	)�D���)0��2cYVܺ�E�5����GK��*�z�T�4Jg�F���p� ����-�0Q"���mQJ��Ib���*�*���kpْ�fOU\\=	���XԈޑi=+�y!`ԑ��"�ĈC ӆ�6H-\ a��=E���^�4�Pr����혋,�u -�*7�v`�6Ib蛖**�U(����@�8�������o�w�sM�5m��}��"��DQ%-ߵ���2�ʳx���46�QBY�4�[�0�g�    IDAT3�@�>��j��Q��\�9{vž.8�6h����p@e�4<�KS3ƹ������<�[=��?�p�
e�p�	�$����ij�O�,��B<��pGzm^Į��јhZ�E+����}��^^����-W\__'/�U=v�����|��w�����g�5�g���)\;*�XԆx�+!�b��E�؁�
�8��#�?i�ǹp\��b��Kv��n��G��G����
!<ʕ�S'yZ(?�����#�b4���Ǆ��q�>�D<N�O'`��?�-B$:Z�'�C�"|?��G����5�Y�d�c>��y9-qܤ8L$�If4Y�	~H��Y��������g0��}ö0Y�,���Ǻ.U6JF�JВ $�;T�}�:@�����K�^�Kp��Y���ĔrnA1��'s!"߮��e�\�*
��)E�q;�D%.�n+�m����J�ȩ57�"H�p�$&/�C�pq��Z�29RjI�
���W��$�9�s�������e�Q
;�H�Uթ:��e�2C��cBߚz���BI��a���F�e	|iV��Ւ��6Y���EU�I���l���x/�ă�<O8��Z�9f&�&\�
@����UM^e�,r�=���(*d =&J���d�|�I�%�5�v���uQ�X)�G%��d.���˹��`ڌ`#��Ҭ��(��܀�t�M+�z�(���O��3C�B�������=�YK)��
�Ck���u�4-��F-����UF�^R,jBL������A�����.�q�`�.-�q���/��V4�E
M.�vH#q10DO�T�R�ZKZ<K��L�M(�?r�s���,���>�mZ��k��=?���mG�e�<��8x*��Y��M�lZ{��sA���>��sa(}XIP�P
i2�R&�X�e���*#�KI��1��xR�K���9�6�<)�u]�܄�+6�-���,�ɹ�<�d���������^5`H����ݖ�O��XV����@&V���gf��a�|%&[1B�@8s�?p���A&���gH��5G1
�L��Qs�>��Lx|�s3��z>�h����cHf���Ǧ*�~�`�v�i���H�����9�iw��.�C����Eʔm�󑺗�<�4��� �܇���@JʴȐ��O���*c�]ϡ�� ��� �O3HQhd�,U4n����.D�c��H�[��cbt�RYf�|�D��EGoJ����@jOm��t���p׶i������FQ��Z
���-��~p�(�$
��9�G�)F1��|q@d�aT�#�a�@4?X�Ц�p1�p�p��d��O�	��E����|N�ԝ��m1%e!Ң�(�S�5T]aQ����U�,�*d�~�cp=}����0}O�#cю?� �#F'����,Q��B����dJ�L�ƬWp�DW�͆���A NXV�O��c�SIo��5&*$*]�UAY����xK��eIV�x!�%.�;�w{D����;˻��|U��UdT�����z���<�w]�,oP�$�A4"E��ZR��{:���LD�?�41�ѭhif$5�[�@R�%�� P�d���m�a�sMV�fbNDFf�{3�ۭ����o�ʊj��U�"㐧����UQU�ppZ^')E�����GYv��,s�D"\L��!�5�8��e��g<����H)�u[���.&�E'�l�P1�V,t3 h�[�2BF/�N�q�Pq�qa8�����"q�b4��ol`+�j�$�����GY\Z�r�ݻ�TyI�Ӣ�����{;��b���G��k�z���[.��Ǵ{	F
li����ե��:x/������7��`�����h��z;�����')��j�]�eY�����eq����6F��%�2��6y��j�H=��h�G�?�����٦���^X�����+�����W�=�"���	�����Z]��Q�j���%%�Mm��>E�QW#���٤�'	��~b���	<_�B5A-y�|��4����#���?i�h����A5k�3)�)�`Z�1K���_S�7�J�>�ɹ��W�L��{��V;t�'��LSeY��1��X��e� S?$xuA�n�n����q�������V�KUz��-�k�j�j�9���� RH-�D���\�*�ZF���2	�Fh	"x��:��Y��c
�x�0*���I���]�X���16���A�e�����S����j2���D�Di��o,�,��5�JXЮ�\�7��tD:����w��b]�_��"/,JJ`E O��`DIU�y�\�I��J��D"8t��YhSjm�nD�mK�0��f+���YCUYzB����ʃ�>������L�C��ݍ}nݾFK��W?��^a������%�#<�i��?�N�l�k�8"mQ�6�ģ��*�/�h�.s��md��~�U�т��"Vt�������p���78�7@Z��	2���@hG�%v�v�P��cd�2.=�јq9�{�T�SN�-�iI�~>�K7��+�-�P�*��1�8����ҁN"��I�WZ��-E^�������,�0��WM�X�n��R8oHZ��������ۣ�=�xD/k3��Jb�Q�$m�Q#V�$C��sZiF�2��Š̩\A�vY<�B����T�{$B���������5:+���o�S6jm�$!�(�H-��)*��2�I��,��9��u��I���>g������xʎ���f������"���o����a}�7%FJ��3���xmF�qT�ϛ���i���y�#��,U���K��q���2F��lo�2�X]_��ɓt{�9q���P9�B��5�L�����q��o���F�uV[���M��[<7�އ�2tKJ��J�w!)}��80�Bq�C�i�� �������P*�51������AY!��/QR�$����ak�HM� ��6�CsI�xc��T��)�.���8wo�*��̥D͂�I�����l�ڡ[�$'����msJ�P����z}�@���k��7� )FX��v��0VR1����QM��X*��9�iD$[G;�I{�E����2ma�%FÊ��1he�o�!�cRgIDF9tdQ��Fz��Px�phZƓh�� ��}XORJd�#�����bhF����ᇻ����Ŧ-q��EF�\Tx$RH��n���K�s[�07B�+O���e�L�T	��@DF���a��evF9ى%�#!�%#�B����bm!���g��%V��3V+D�%MR
�q�N ��)AA��#�@CoM�G★V���{����5��1z+,w��w�����e���ڙ3D������sEp��
kw�8�Ne��@)O�@��� I$x�x<���_�ȓ�Q��ʋ�G��"�E��t���{<�{���3�s��7����W:;�N��YF�.��DB�I,)���/�h_���a���2�E`�c*"_Q��X_]�n>������T&�	Z�����Gh�I����6��sh�;)��X�9��&�z�ÊV'���[2N�R�Q�-���8��X��v��xwD�#���}I�UUn�j?
��TD�B���CZh�\os���tD;Ѩ�3Ғr[!UF���v��mR4�wB�hLU�(�'�<�i�Z'cW�$���n�#�����'�S �����ї��5	�&�j�g~��ڭ�'s�����j��Z(*d�ֱ�ft�k�K�qL0��N��kȴ@*(�q(�E1�JQcFň7���رc<��3��x�A�w+��<����k��X)Y\\b��qt�����x0��<���pQ���"���Cð��bLEP������N>��
R/q�B)MQ:��T;C�b�ILUxr�k���g��I�6��2�wlY�p4=9J�f^�zpj<|��;��[�����<� <8�Q+�52l�,J�:���Q�{��T��V:�����L���ｌ1!�R
Q+�5d���h�9��G q�缴��gS!��k�����Ц�
�7%N"�w���b�����s<��o��+?����B��-����E�>�0�w^���RUȎ�Wo�{�$4��4��pΫ��F�V%�?���"��apa@�I�C��ae�5�ʃp�`Y�T�M"�T��($B
S��&]�̃$�"'��ưr�3<���9�'�K�6�����Ȩ�eū?����]�q5�۪ڋo��iw_wsI%%Z*��*K����|t�6��n��"�ݸ���E����}g8��Ctϝ��#�/=�߽�ۺ����o�H��(k�T8y��$*�q�e8��=����?v�ň��ȫ!������SDKQ�l�4Y�ȉ��$�k)�� ��4����"�C� ��eA^TT.(�	�ϻ�����"G��TN2�-�HA�(Jq�T��ri��GqPī9Z��6p�0�Ag����ʁ�,,D�H�Jb�O�ΓJ�U�Mק��I��N��-�H"�blU�i���^NH��D����r��(�q֒X����8Y�FY��
OE���ȥ��%Oe��ֶ" $�!�G�y1�ٳ� L�D������r5���'{���J)��Ⱥ��Wj� �����!�~�v;@�EQ *;-�% �y�c�r�u߈�^��`�ݻw�~�:'N�@JI����i�q�]����&�N���ʂra��x0dow�*/H����*G�!�2.\���k7h��t�ݩd��C�b7q�xF��I@	P�bX	�DMI�q�I��`#���������v�L!��Η��Mpc �B8h@���[��d����>��z�u
�;��1��s)���8R:��t���{7�ɯ!&�����Y;Z�~������qk��i� x^N������|5*����q���y����������a**c�(��������ѧ�yύ�����TÄmRB��?j�_�8���h�\^�F1&��:������$�T;�&�W!��Ř�$×U@�����.�@�Ҙ�Ԇz�L6
[�X#:K<��Wy�+/�vd������&c����j�&�ԣ�����������ڈ)!�5qH	ХF���fQB��"R`��,G�����|���]���u��i.���>�W���ĉs'h���sA���6xQ;�Anb)P��z� �뱅�,J����ezkk���9�����?�H5�8�9���(�
IYI�B��c�91�!eh7k} �� q]���}U��t�q
��xDG��`��2g1��k` ZDآ�G)cgȫ�$��YJgơjxS֬;a}��"$�n��j8��!�R�2$qF����9[��T
��15+������2�X�o��U��޷��+���BĬ�Cai��a�P�v����xD�Gc)��W)5�U($V�EI�b�uӱpJK�Wz�Lg�������7�?gϡ���~��� �9#u����S �ʗ�D7z�_��lS��3h�J+h�;�T��}PG�~8�I�$	����h�`0����:����]��鰼����uN;�~S+͸2lllp��e�ܹC��bqqqb��p"��օ����4q�a�������B'FS�����65����9��ƙ&<od������vMny~�挤�e�7?�k('0���{o����)��>x=�:��򽾑�UQ�u+S�����5{�}�?�B��ש����j&I1i�1�H4���g������߃�Tã�����9���t��C��w>Tg�������
������[�E	�p��#��|��k��u�=� <�,��-娏��z�C@R�M�?������D� ����Ho�A����3�nJc�Vڦo�@���������;Ո��Iu���oާrA�p|��asi�N�uđ���c���p�_�����_�7Q��_�q�����'��,��Os!�"�!�K!��Tq-)c1am'��J2ݡ�$�b�r��ϑ��Xai[�͛���L`h�F�ȲEO� �S��ȁF�^*��vn�@�n�b(�
)b�mk�/�-w�����1B+>H/�\E��_��9�zF�����$g-�*1J�@8I�[ʲ
��D-T����Dʜ����9Iyw�b�@�N��UCk�u9nu������77�mz��i�&P��S^���g��d1�x�#G(R�mc�C���,i�:�V`"���ʖ,ʘ�;D5�iJ�t�瘟:�2�hyDh`��9RT����$!w��bLi�TU�CuJ�j�!:V8�J��P���@�yo͓�8��\�Zin��YsJ�Clƿ4�?,=�I)������	�o�D3%�ӡM����(�pv>���N������G�j���v%������.ֆs��V��Ͷ(���a������i�P�<��>�n�
x��nO�i��+u��=9x)���u���[xaR���M��m��:��u��	d�|�ɑ49� 1P�>-�����C�����������+PZ�肝ԛ�P�@3"��O)%�����><&�r���:g�'?�O]�F�9P��'e���r!���QS�јx�30�!c9{��0�[ ��f�z�m�ֻ�r�i4��t�a��)����ѯ���҇�ƒ}
�W[�F���oxkT�[�ɖzTJɔ�����q;�Z�>̃G�R5v?MJ$t[�1�4��"�{�q����>��VFH��UYҎ4��.��������k�"I�	��Q��>�%����j�uF�@�Z2p#N["Yi��q��~�c������Bۈ��/s���x��G(��
0xT�� غ�;�e<�&M�'=@�L�!�lm�p������-sَ��9q1������-�FG��>1�q�;�u�b-�"�N$�P�o\P���
����{l쎸��{��?`��-.����]"��Q�"%ZY���'<��/r���q�V�%,�ek��5N*Jk� �,Q2��\US���Bp���?�s�ݼÛ���d5,A�n !;w����8z�(~�>��U�qe@jA/!�N�q��CJ�Z�D�XI��\%ة`����N���S���y>|��<�ه��=�¸,l�w�2��-��5��;9ǌn3]w��$A0)� D�q�����)B%��~�yBE
k�Yb��J�-r�m�p�����g�l�zc�E�jU���>�g͡�����>����(��}8j�SX�:�Z!�ʔ�vV��i-۴ߝ=��(BɈNw��]�@�N�h4�/r��-��sb��jF���$�zR���c�]���۷C �LhJh�n�iy�#����(�����^*b�pDQT�Ee�-.��Qpb�)o,��K���qu>1e�`�N܈���v�������و~Ɠ<tB-���O���$��Ɠ��C+�|��R�R�0�ќ N��aq�w�>>���@K3�`6�(%5��VL6��s������}~vτ���s������ԂC��Pf`�z��Di���n�.�Q�=ZH��w�wvI�U�������ܸ�jKF����ٴu��j�	�St��gL��u�b(}`����V�@j�^<��~C/[`7Ӭ�����LU��)��ݼB�y��Z����I}�T�fc�dQj B	d��qA"5/���]��G�@e�s�r,��DUF�������1hE��D�1g-�Me�E�vj�R$Bȩ�pd�ܘW.a�,q���ֱU�!��TJ�8#Z^a��yq��͋�e��^C�GJ�*h,(�fU݃a0֪}��q�"6�i���7���O��YK3��R���m7f$*���2��![ﾅ�Pnl�����C��Aǻ,m]c| -Vc\��9O�_���>�ay?ɱW.�H�0��x���SϾ���K���:_�+���u�R�ڙ�{]��"��밭L�����I�s_�=���;>~�"�Ns��ɣ�=�ʑe�������_��+?5l^������4mE��Ht�ypU�{u��Z`��J+&Y\a�"�E�PjTo���fw�#jEZ    IDAT�V�8�$�M>ܣ��Բ5iLU��\$8�WKQ�4q{>�rΓ ����１��ʹtf���r&Ⱥ������؄K0�xCEI�iVG�9S���D�SUU7gT/�Q�,��8�����7n�@�P�_�%� 7@ȿ�x�K��"�Cka8�&$��dúo��6R�͙������j�{�R�TGEE9������ڲY�\�)� �� ��L}��NZM`�zJ���M�$ 發�a��?��_e�� ����:@���}*t��Ej|�5^�a������î�=>6{��fU��o����g������BqP����|�λ���=�-q��	��V���Ўӵ3������G$+��z]��;�P:�������K�B)�	hI^yJk*Ԟ�=B�%j���t��*���o~̛��;�}��v�ۦ��qB�<�Q�����,E��2�1�8�56`]ȿ���]��Ό��b�,i%1�0d.b_���kl,� U��PF�X9���H����H��0�<�|U��P+dDef�}N棾/'=��s��Wpm�g�~����#��n�~�+�
p7�p嵷�z�cZ|(GHI$%J� Z�@H�sWƅ!�8�FA\ԃ�T������X�u�߽Kn*�KO���,�bd���*��ǗYW�Vѩ����:��P�,Un��4�lt&�����l|�>�����?�3�~��,$�����ҥz�>���<���]��/��{�9�.K�8Վ��:!�` A�JȺy�����u���u��XLڼ���{x�_�ܳO!���_?O�����Ӝ}�i�`�wo���1���\������	�%�DctD��gx����!f0&����죅��Go���w�Ӯ�~�Y���R���܇dT��ٓn��y�~�!l��]���P�!����-��Ҩ:b��j�'t���U]m>��[r[��`�~4�؊$�a���,.��j�fZ�Navc���T]�i�Y]Me��-.��N���;&-�a0p���~*��I�%���zU��b��'�w`�$�VUh�2�N�I�%���,T3U��`���f!������S� ����r5iB�eq�Ry�Dk^(EN8;��w0��׀޻�g��f�f_�@��y�4j�N�|�>�\xp���N{�/?i���~oJe|S!����j�yB(�^��ps���O>�<��p���b\�:���q�|�%�SG�_~�ŴM!v�bX�v+!V!�T:���`���҇�mv�M~�|�)= �#��7/q��Y�d~�}�Ɣ��!���(�G$$A"G��c�*��k�{�2�t�İCZ�E����wٿ���[|�k���ˬل�)�*�|�e�%-�Ȳ $Y��׈��UB��f�R�'N@�S��l|�.o�nr��N�y��J�E��x���y����,u���o��bx!C��H� N8���r��� ��f5�����.wy�gy��_A����k�����o�	'�}�������[����F��e����Kʪ�)��T����i�mr7�g�O(C�;�EM)J.��c�S�������|�����3��x�k����|�k��x;��{R#A��9Lc|�|MUպ�cL�E�hU���.������8��s�G��%$��!KRį��{,?œ�m�{�G�E��3�D���g,KKt�1
lu�|�¹G���v[ܢ���R|�����e�jĊ���z�mZ2"���5�0�`gγ�;��8��<��O�>)��}~�{3���� �:�����zj"#���s3��~"��@�B�:/����u�]�B?���WB��������q��n�)˒��� ��5l�	scs3H�ַ��?]C�Sv}X�q�T�b��o�ck��8A��xBC�	�M�� �|~�4Z�8Ϟ�$B���c}�����ZX�z7!��=^�Щ5g@C�l�l5	���.�U+��p����`N>��SI�ۦ��Cɰ?` E�+���`��-�>�y_�wCl9��&9�z���4BW��F�>j �iޥ!����MbŽ9l�tS6Z��;,��R��� ��Xh�����!��DMJ�П�	pO'Q\>�6���>���=����N��vA�CE�*=q�M�nS���n�l�lӖ��(R-���=�8��ȇ9���شc�"�����@H��aQ���qn����o`���+�ݒ�^�m�EKf��m�q�4P{yA�3d-Ϭt�D`�z<�����`Y���.�l�X�ٺ�7��O~�9v�$�.Y,aP�D��CW�d�����%D�N�����Z��c<��B�0,�(����y�%IG�G����z�W���=bi�a,�Of,/���"�Wo0z����"V�ω#E"%��(�TJ2J���
mJI9�Qv.<QǓ$r�,��ѿ%ZiQ?��3d/<�����C��n��Ǿ�Mn��Gl�����)4��P�*l)�S
�5�8�����q�BR(O�-x��gп��_�K��N�%:z�߾�}��`���K��q�]���DI��P�D��	�g�vE�$�D�@�	��pP1�\�ӌ7�)�6ؿ}��Sg����*��#]67.����� ��.E$�s�V0�3G�-�ǎ�$Q��	IK!}NY���|���+�}�[wn��?~��k�1�����I֏��+'��'��9���0����"'�Q�
_��%�P���ǁ���CK�@�(%�&�W!%B5�k;	$!�?��Y���&ha�L�5o���.�}�(�/عu�U�`� �F����)t�����q[d���U�j�xc1U��Y�h��J�,΁��(-Y\\dЧ��`��bT�y.��V�HMȽ���Hy�-J���(BJE%�=����ߣ�͐��A� dFYT���۪D��-�@����#b��R�L9b�����TE�":x�_�7���a����&�3!�zj~*��9:�s��X{o�:�����;lll��^dJLɁ:���k&0�����{�@���ڃ�~�L�3���=��j6���(�a=�?	I��O�,A�m�7$���N%��q�4��l���_�ƫ��sf��^��lc��������l�s�|�!��|�? �̼��<�?,I�b=�	����fh޻�������B��m����k�ȅ��צ_�ĺ͎W��%�G������,+�{X�2&铙T���$��q��{�nEU�Q�0ܮx�g����=ZkK�:)%1^	����cW@���O����T$Z�Т6�����Z��i���%���±��gx�+��������E�t�'^�gϜFZO����?��������H��Am˺����3��)5N��d�
�!"n����2��;��׌v�y�[��-q��Uv/_��V�;�#>B�q�߼�.�"����e�p�Or�Ɣ�s����ƣh��}D�M|l�;���m��K�je<�䣼u�=�����G�z
ٍ��;$�@G���QxbRG$Q:ja�8���Z`e�)M�*rC����g��O�u�Dm�5#Vz-�ύ�-�k���q�E�C�38������뤴dƸ3.r��B��Jz|��.����?����=�E^r�4}�E�Y��=F���J*gC�d^g)�21k��'�#4�m�ZjP����f��)��E:'�"DE�����N�[?�>f��j[72�UB���:���@x�T�p��9�iPf�:�֚(������ ��Z!o�ki;K)�b��([s�Ҵ�qMT��Ji������*Y[[����p��vw�'�cʰV�r@c�Vb��(�1�ڛ������\���U�'v0'욨�~���:��'M�'M�$�?#�כ�'��5����.Uk��	��l��|`=7�Ygc�}l�*���o�����c3�:�ws<���P� ��*�C��S ~�5^O����C�������_=���}OwZ\�v�wG9�}M��Ak�"֊Q���^f�V�V��������%����=�I���dۖH/�X��4	���%���
�'á$<8���$��|�A���3�W�q��B��K��Ω�����ӨXq�W���kT�1�Qv���}]_��٨aV�p�В�n�QY���6�ޥ���L��,PY�%�
K\�cܝ�@
B4u\ �?�ta��_p�B١s �"���{���?�"����6����ǋ��׬��8g��QV�e+r;f����������� �Y��b�n�h*�n�,EP��DL���5�����q��(q��I���;���嗹��5���,?�7�F���������� ��A��A�}���	�	�D�pV�ȓ���7��Xj�Г��d+�,9�W��䗟C�<EY���~����Ur2�Z��ڠ�G* ���Պ�ð,)
��i)ؽ{�+�>ʹ��S�Z0���o�a1j���ϰv�8�t�o�A�mM���56�rJ�TQ*�j�p��_x�Y�v�2:R�*$q�d)�;��9�ŏ>�oG��!G,q��p�S�N�Ѐ�M���z�������P��a���YƁ���-�_����6��������A�	�|z #�D��4���׺��ژ7n�sQUeY��������EFGh)W�j�|c�[i���F?R�$I%Rjt�T�5Q9O9
mj�3H��$	�n]���� ��3ܓ}Z�*������^���p�&����I��j8�S'W���i �������_��O#��^��A�Om��RAך�hZJt�911�A�|�>L�r��dj�m�13�����3�4M��%�P����']�����pXl2�p
����
b�����;����}=^������YF��%[wn�}�4O���uw����5��>-ie	EaqR�d��Z��'����(��V��O�q���H�U��Ǟ��/}���?�M�����y���d��3�G���������`4��A��Ha��q�]�>x��!R=be���x�˿ϓ�G���{�%	��*��;�ΠZ
F#�������h�OUUd*BjT����`�B��@ �㜸��������eƕ7�g�=��S����?ύ��om��:�˜���l]�����3���{�qEY�����a���"(�#[貾�N��E�t�/�G��p��!Y��������H����Z1,��y������� .����Fdd�=� �{���KM�Z;��H�O,�:q?.2�����?����|TW���s��@B�J�"+Z�Z%�3(KF��z�R��������_��ٗ~�����+�IU�͟��k�z���x�K��/������x���>:	��򯟞-RJ���z�"EᡨRZRgQ#C���Y�qe�:�)0:��.��_�3o_�Ɖ��?�*�v�ؔt��!v�::|�0�u�U���a���~�힛�YGA��}hϞ?��3*<�����~����_!�Q��a����_Q9�h�`4��9�1�n'a��CUU$I����K��I0��S2_�$$Q�I����uEK��"���!���Gv}�����w�ܭ�%�·�R=Z*��H��&�~��Df��%�	!��Դ:�ׂ�!t�M�{)T?�r�L��榓.g��~��E�3��y��u��1A�Jb�Z�l��V*�W����D����+W�[�Y��>��)���&F�NY\�=�Þ�����Ĭ1f:n|�b����s�8[�{��ɓ1���4��[�=���K<��SE#~�ӟ0v� �V[��i��W�.GD�En���wwH��(+��tT���[�%�z�����J9���fE��c�(�\�׎����,�� �C��'JZ<��K�}�I;X*v7�8�~��/}�;|���;���n �/�s�mMnd:�I0��Q�q�ދ�ng��~�\�@7����UN������a�
[�/5�)�7�S73^������%N>�e����.���� ���/}�B���?�g�,,.���kN_��+������Vƹ!H��p0w0�Gx!b���`gYZ����:k���E�-�h�ͭ�,�;G�����1���x�$Bi��':�Ig���s�*�T�巯��0NXH,$B069��%l^���de�����x��^A�MBs"B�DI�Xz/y��|�yQ2�,�p�	!p�U���k�����͎p��9�,����{�ט�;���^����)�kwXZ^
�3�:+ڤ��x�)"�X)(��b�7��O^f��$���=���}Ȳ��]����,�X��������cL:�ٲoqZ�I᪡|_�|���)���MX����ΩY���ο�j��Hش���bA%��B� �sO��^/ �P::�Y���u��D}F<�׎_�g��	`-q4e��1ιI��$I8z�(=� �~�������
�*�Cloow���^Y��H��L$i�ی��	c?M[��^Δ!xl�Fe��j4�.�fޞ4��dCMG}�PS�٣�7��䋉1������I�;�gZO�a��r�Io��(6�)x!'�҈܄��N��B���f)X�ZJ�L��a�L�V����n��O��nλm��It/�}<h�����|�0γ�^�`�9�j�)�9������73��)DM�s�}�D<�#O>͓��X8r�ko�����He�$������k��=��jBl�?�9��-"!P���r���GF6�u�X�8C���q��y�c.�����N.�̃��_����s����<��o�����R�+Bn���'*\�d�s(��{�]'����]��������dLe!���.�>�/|�ENY��y�������K�!��oeU"���)>D�k0�FH*A)$��%Z�#��=��2V�d�侵6��|�1���7����"E��
��x'(�9�Q^|M^d,�� �37k�9A�b��❟���'Y;}��^���Čr�tȻ�>"Z_�?�W,=�z�i�����D�U��;�>���tO��Y8u�~��c����w�����,�8AT���@K�rN8�:�,�Qc�ƻ,�X����ꔠ�!��(�[8gQq���Wyaq"(
!�ƒ���$&V��m6�����'YV����Hv���-���%n�_�;�_�)G<��9�.����~�)�1<Y,��1��a�3�ttF�s����/摧��K��C?.��DG1>��?y���m�o�`1ˈ���	M�5���:O��a�'2�t͞�R�,j�ݔ����v�b;�"�,+t+��{�hҞ!X�Eq�F�����Z�J"@����]�u ��%yYM�eA6��U��v��YXZa��F�����n�0��Sw�++lUR�P��������y�8�也��3�OR��������#s���3Q�������{�@���k�'�P������l:b�����D�����;%�jt��hU�I���f��n�ܩy����ק]�@������`�7��uAvx򿅘��?�~��Ձ��'��Tpj�(k'Op��5���O_�Ji���J�Ď��[���Ox~���UN?���ߦڸM/͈�����J$Y��Z"pT��ڠ�h��ݺf����4Ӭ��P�9W/]�ʥy���#���\~�|�Y=� �/~��.+�����[��zm��f�ɉ�y����}
�H��r���wಌ�C�s��s<�ܓI��>�{����?�j{'85*�G�m�Xolc-����f�ʜjbM�k�4I�q9�jF��QDܡv~L�Q�㽥.�SY�(J���Cf�f�7��fW/�cERT��~�c~���_��(G9~Pr����o\c5�э��d�o\����GcD�	���A��Y�������X%��bW8��/���	���O��/�s�"I{)���̟������_�wq���1΅��q���D���$�u��"/U����CIO���c\ZҵUN?|���2��G���ʣOr��'�xg���}>�or��[t1H�b���7���G����!�V��b�&���[����o6    IDAT��g���%|Q�)E^�!��Y[�ڕk��w�'�^��	�O�(�,���2N�Izn��\�&���\ӹ=�|��jַ�
N�3N�������ʐe�9{�i���L_#o��Ԝ����؇��*��m��i!')���ڛ>iv\g~�\��wW/��}H� 	��"C��xd�c&b���#<�cGxdK�H�DR@�$�}i�t7z_���z��f�?��R� 4�D����.�y��s�gmm��h���"ssst�]�f��� �$���+��ш<�Ɋ>.	�6q����>��1_�1�O�S�����O�y�����vST�n����J)0`]�$�����}�g�XM&�2e��j�	t?�E�������B��F�%R+T p���ɾ^3M��NCK�Ԛ�����/�DS#�`V`F=t�w,�U=Ӟt��oN�L_cƁ��N��b����z,��N���@K��ZҬ�xTRd#n������Ivnq��1�T�$��F7o��JDai�-�8C�e1 �.
��~���ީ*�S�� o�ए苸D�ݥ.}[r��}�~�� C�Li7$͈��&.V����n��<�7qKD�S����V��t7E��#LQx�H*:�9��S|���s�)��Ko~�[?�[�/��VDhy��)yE���Rzm��ຮ�A�l�n��Ggy��&ͅ���7�珂��es��r��/����@N���&�fDi$�aB��h���2+'��Zzi��$�>�E���7�ijV�0W�.�d���ٻ�Ecn�7���X:�	��ƍ���hx���sU��Ϋ^
�E�&כ8��B6��avR���_��W~�i\z�#�/mq��A��s�6�;)���������9GWk0�}�7������3�!{��<-0��DK�)�b��e���<������Ga���[̧G8����3O2��"Q^r���&o��Oll��+�XT��a���e�,:�p��\(3�ɀ0tt:rk��3>8�)�C4È60�ޠ�i�j.p틫���m�-�EM��#��pj/������ѣQ�UE��x����tD_�Y�HG�@���H�w�)dY~�	���L�wc�Z�O�gK7��au�����;}o�li��y�ߗ��]��Cn������ѣZ^��l�0���;:��~���>��;���d#�t�19aN;�8����$I�D:�^E��Z����We�����iG�d�Es�C{8YxQQ9I�z�AU����`1���D�Q[M�0�h����yxO����h'(�t��@��q�I�r K������B`%�٦|������
"@��jkY\�(��/H=�ճ*�� ��:�F jF�:73ml��P���:��v"�Q�O�&猛vh��k�P��.[XL�EU����5�/�rճ����:�ݸΣ�G�r�4[W֐��Fl�8��T���$�>�.|v�^o�Jܤ�$Qͳ�m.,ü`X(ʊ_K[�M9����x��G��c��ɥb�k/��覊��H����e�x�����4�l��p�^�"�c��;W���T>�We��t5�a��#T�g-�㧹��9��������|���\����C-��e0J�ʂ�T4u��`@�4��(D%�d���5��D9� w)��#��״v{��wy��'$���lݼ�������y���Շ��?c�)]�hkׯsY9�5�4B)DŁo��8O�#��Rzy�V��}���{o�C�Xc��Xp7��O���/q���g��V�B�p�JtP��J�׵�Hz8�֊zO�X��=iH:DD]N<�$K�K��{����`Gܙ���"��F;|������{�nң��{�Ì�n�,��KO�[��a?'O�(d�H�h�1JI�2Ñ!÷^��^�V-���[$�e����SϿL$����/I���?��~�eO\�/ECE� C���Z�O:A����ZIB
�ҙ��?Lɒ�a;�'E=�1%6�g��E֯|�f��}Ϟ�����]����������
e����C�!m�VT������(�*2߱Q�0x����8��9S�U���l:Ҝ��M�<�&X:�,�^��� ��;�\�B�ґ+��)������cօ%-KB��"�(��PE	R#��sR�ZTHE��(}Qf�$��@�h���m���yIo��g��޺�֒N�ñcG�t[t���(y�������ۻ�����8!X�4s��4#�`�2A[I!�WH���8)��baV�\��
[�*�0֢���I;�G�H�%���n�s��q:7}L��Ɛρ�����w�(v�����������_"����*ZSW�)|�5��7�O�"�E�+|���/s&; �@<�0{MϠ6{��u�\=b�
N�q����:��U���Xߎ�K9̅5�.���+���������-�l�H�4JI��¡�?G�����¡�#OR�=��C����p���&�������׹���<�����C��}�e1d����9��I����iuڬ]�����a�{�]���3�{����F��C/�}�k���K��%ҥ.�l��R��z��7�P ]���/X�-��}���U^�4Ɲ.i���5�	N��Z��|��(c��U�~��N����Pin^������Hy��<�5:����|��_����%�֔�v�����J��Q�M�ݞI�ی�O��u�����o���G�C�)]��V�� %�;�l_�εss���)�	a��P915+YQ���UM�ITu3��dE��i�Z��h�vo�g�X쒦)y�1*���pk������<��:D�!+�e�颴$YFiT��Rx�Kc��#�[jr���w����a��g�Etcο���{��L��ǎ��j�c��͗�8_(��5H�0�(M���������~�=����f�F�$}�>���_����I�}��<��1����b��O��"�%&�R4�+� P� I Z�*=8{oBH�*�w��B���^��A�3鴩��i�K�����Y/W�$8�(�h�5LP剳1>Ǹ�yB���� �>Z�Řɮ�l��0fBe�$	E����í[7i�b���8�z��N�v����<G�e����ǰ����!�VU��;�L%�X��>p�i�	V;	����H=f:�����k� �!�3����=;1�m_�*O4��'������+�@%T��A�@4#���I��r(��y�B�J�N�����D�8�����m��y���ń{z:bE��@��\"�"����������4W���p����y�4�>��s�d�=t1R�x���oc���ϵ�s�S>��O��	(GI�H����Ƒ����z��瀡�]�pī��?��q���Oh���V̹������s��~�#�Mn���O����9њ�W&��c�y_�SG'������F��
=�.�M��}�ֆ)NG�EmNe�	�7ЙAE1�n@+��˗�՝۬�.0LF��1�pPR�g� �_Ͳ�OU�N�$H���7x������R&��=��MZ6g������d*�ܾC7/�E5�B�q���t�K9)v��0P������W��3O=F�F���s��!�����m6vw�';�#��}{�d�S��&Z5*��	�
h9��*�b\�� ��XIo�can� 
���b0�y=u�* �1�<gX:L@���IQ+�C��	if�����&;*�dA�����C���~�g��E��C66n�5�~�K��0��S�dyBZDbB����O��"����J�4�� d��Q���[��<	5�M��a�{�lc�V���sr��G|��y(((L���
����!���Eum#�8ms��_"���d�Ljzf�M�����{=9f�ă߯����T�f�?U��3�BV\�|��A���s�$G�?�<�RQ�Jt(C_H�h���~�?�o��Z^Y�������{�{�a��|�cǎ1�����G�N�$�ᐹ�ZJ���I��+U+�Nr�J	�RH�q��﷫��V_a�5���z�:��=�3�L�������??}��X�$����tE��1���C�W������v}��f8ʨ�8x���T^��1�@�,z����wE���xǹ�/�'�6����Ы/̨�´y���ل���x�~�>[!e����o����I�m࢈���\+-�~�����WA��bSR
��$��i!*��:ΐr�&��Rw8��	���ؕ���˭�]:��������f;�"�s>�-�7wnnp��9"�����X��a��M�ݸo-T�P��� S��:���u.�o��V�f	�N��'%т�Q� ���F�Ҏh�HJ�S����P��� -|J�{BL�';lap�ߌ[�����`��,�癋�5b�C�M�n��C�EA.d��^�H	_�(�Ƥ�ˎǨ�_�՛gLJԚ�o|��>���.��'\��,e ����7H������7����3|���y6v(�׮R��
S�71�B<<�G(���M��>Q�h6�)���e,.w(s�����g��-���o\�d��#� $�q�Y�(1N�U�-+�D�C
�2�Z
t���;ذ���2��6Y�I�ls���o]�S�������Cv���]ύ�6^ˤ���ˮ���	�8H�?�C�WWi
ɥ��坟�-�AJV
:�>�w����|d�߸Λ�7����v��~�g-����@q�u�RW�O`�d��*�|�Ez�\!$j|�r��$��}n�����^9޽IۊV
|�u$�8:B����
l1E�cU�����������j����o��R��O��E	G�;@i-�`�p8ds{�f�I�w���]/~#{{{�F�G���c�`d�W��T0:=�ui�W�z&rw n�������~��dx��/������I=���>�q+��2!�M��
JT�eI@�K���E|��uΓ�j��ɧ<ۃ��{D_q����Si�{u+X�x�O<�/qPꟺ����ߝ~�jQ������V�čyvnor����(֨f�*@G�	�? ��#�����ѐ��Q�Q�O�s0�j�]%�;�&��߁��F;`��ȵ��#�r湯3�F��C/|���6���/�<�v�'���o�����vv�������];���=�
��q��8B͘4-y�������C�����	sI���$B��7dny�8Rt�}z}Bx��DZG�Z��ЪM@G���� H�zX0�6J͠,:M.'6�Q�HG${CzIJca���p}}��lD��DQd>5QGf� �htK���c�_�4^'A$��ǏG�������-�;{ע_����!X�F�HF��2��"�7�ZG��G)��K&�2�8�:����;S�б�7�3\��ӏ!�H6�(��,�(E{�0�G��n� _��r3$�!y	�$'��u^�p� 
/�,Z�V�P9B-}AԠ�\�!�
�e��'X�=�O=�B����wQ�G�x����#A�
��w�����[�#Ca���#��K�ѥ����[4Q�Q���e�ʲ������w?e��yYŰ,HZݤ��a�>Ri_u.@*�FW0�w����M��r�@_�#�d��ʘ�D}�1�M�zw� ��g��;]1 �ph�T�a�(i�4����Ϡ����
��������X�ہ��P��S�[_�O��=)�2'�st�X^^�8=�"���i�a��ш1E���.�v�SE��a�!�
6Ձ���5���)�e]�>���B(_nܦ#t;c�k���>�����������E�W�EQ U@�lќ�%$)�,	-��{D�����������]��U�����Ǧ�y����9=�<�1/Ϝo��_�<�q�痤�H�q�K��cy@OğO�^�x��~đ���z�㲂�����W����\��ٟ����P��p8$3PZ��>�"��z��g����9�,�pPCd�C�h����^b�����O��G"���D������Ar�Cn��&B��\�9���ȩu�8��^)�
4^Hb�[���?�5���3���=��ӏ�&\^�Z�6I�:�w�CG!&�y�R+�/�4���<4��G��� �0ړ�h)0*`���X8~�k�?a����R���䍜�Q�`}�ha����$�h����#U�3<��"BH\M43�>��檴@ۂbw�a��d�����%kJ�X���3Mn2�#K݈h0$
C�V��x�ӝ�cA+�Á�ug�T�R�8O���s|��^��񭗿G�m�ch����]�A�������}��.��%����<#��%���^*�F1�D!�@I�D�$4�ڔ���_��l�X}�I���<����~µ��8y�$/��-�VW�]�@�v���8WLRG�U�)k��bV3h'q����PЌ0͐AV0R��6)G�E���}�w_�K��kF��>I���Жt(H�WGl(E�,����>�V���>n�*UAn0x�/g��]�]����W���!Bz�9���������"A����K)�	��,>&q��nݕT;A�����s�b�wʃ ��nG!�DA�(��WQ���L�em]i���G8g�Z�:]���۷[YK�*�W��v�N9;���3�_1=�= �1��W�^g�g }��L��N0�M�L}!%_f:�&�$�H�z��|��ѐQ�������!'�p��tt���W9 ~C����F��9����H��{�o�A��ѱBx(�X����� t8���>�FLZ��9���Y}��F�m$Y�ShA8��|���<���oY����V��` A�R��nϨh1�w�X���.�`m0�ї~��/~���<z��+_�%�}��}�љ	��������ߤ@�p�H87K<1����F\�_h�������/�o�៰�����K,��G��"'���bg��)Μ�u�����$w�h�Xc)�!��Ҭ�/���GEh��(>��9)�"�_
N���;4�g�R1�0s]N�s��-��=�>�g��0�׾���;؝MO�,Ę�n��`N��`��[��HA�|�Q�q��Y�~���c�������>�l6�Ɛ6%�@0��Dq�0�@��AUu4A�����y��6;?ӌ�Ä<ω�o�-��w���O��%;f���;�/.0���i�cG	7/}�ƭ+������-�tDs�If|$��%v����Y�:��(Bz� P(i���Ď�t���v������/���_&n���O~�ګ�s��y�{�a6�����ˬ}�k���)N�$�#����0%��h�tBD!A�k�G�-s�o���=��@�7@�9�=��|���/(�c��$؆�_����f�`F9���.,��S�ٌI��4bhMU�:]�<�k����O_�ڼ�Cp�����C���]�l�#�VR�eQ�&����8TJ�%nk��{ٽ�/L9�k����V�8vw����A��vU�+~�%�)O)_��9���  P��u��,��YJ

�<GBGcq��fF�p��:f�4�y�#f����U�����M�i?#�;v�X�\i�JaÐ��{;�lm@�0�i@v�:��}�A�3��?S�:��9���jC`<�8���?x�i�t�u�����t�~3�2ԕ���5ݯ7&ο��V_s�å�~�p��Q���#6Ҵ�+,�Y��w^b$�槌�7�4[���_�%���b˻Q 7Nf��E
FV����ϝ��_�3��}�r�F��{|��G��L��w������T��]����y��.����W��I�	5��f��Ch�峷?��_~L��IT4O2�\��S���#����?p�S�}������:a��v���y�*777�#�YXZDJ���&K=�(%Y:�l��<bi��O�XX�r����Ӈi��x�}��]QP�YWV:���n���S�B-�9�۫^:���th%P���!�(X�|�g����Gx�B��i�B:�"�
�G���A��	�����װwv���#?YF{JҬ(���e}s����i�Z��z�Cc�� Ҁ(��
�7.��O�q����)��Yh��=Za�C���&Y�&	�QJaJ�eQ �P{#[KHk�x��    IDAT)�Z!(�P�l:6w�������o�0֮���}��@q������A��}�����d�Ts�!�nV���{����vز$Id�e�d�cGO�H�aF7)%(����s��	Ոs���o���r�:aH���YZ�y���KYN�vsӠ��UQ�NC��=ʍ��1 '@ؿ��Ի2]��e��x������6���N�V��H�c��s�R�� ����w�^窟g� ���5U���o6��y>>�p8dkk��r\}�GI�h"���n��b���gq��,s���0bn�à7�EvL������U�E�ϒ!���Z9�B�ީz���� /���RZ5���:
��RL�;�~�)o��I4��z����@:�5vlt��JY{�8'3�Vc��ţ!h��	\�4)��>��=\VPV��F��cdsB'Q2e��J�@�
��ö�s�(�������<����VW6�C�PCd�bg��% k�1�$*jS�	BT��[K�A���-[��C!Q3����:���"����ϗX��t
��>x��>|[:V9I�`���Gy����Ïq����I�����w�0G@N�EU�E*QU:�^f�w�R^�FTyj����K:+���P{l|�!��g<��\�H���$�<�^l�]��?�s�.�eQ��xe��Pѿ�5寝�����%T����E���Qڋ]ַ/q��ߐ]����~�Nc��T|��|�W�.�O��{�P�H"Q4�aX�n���a��~o� ���ńHr�p��P؀���v��v�Ao���h6{tv���s|��΀�_x�G���7��PC"<��ŧR���J�s^�C\�NE�(mP�C)�9i Q���?�W�{�	Z�>�"Y��\n�҈�i�4	��/����7�]M�M�LR�LP��̯,��l3�ߣlǴ�g ���,	U@a-2�#v�ٕ���p��SdW�����ϱ�?{��<Iwa�C�v�.p�����Y��aR`e��y,ZJ�0��1K#�y"� �ΐ�
B��d7Oy�_��:z�=#h�/�g��|��zC\�!#W�� �r��ϮF>O�(���	!��� h��̯�D�*V�[[��-�p�,�i�;��HG}�ؑ7���\�$N���S�!�=�,A���g��9��=J9zv�S���_�SClC�1���-*Ii-��� SukX*��^�/*411�㨿r��L�i�:�/���o�@*DE^��9
��]�~	72��eH�֖�r���AE����Y���dC��X�#�<O)��("Ԕ��V��Bz�^��}C	(�,Kp�H�e	iR dD@��%+�j��0�z1A �Ԅ�!IS:�s,./���0f��Ė%ySP$C�+"G�;9��(+�x=�S�b<u�C��B^aP5%�C8T��~vk#5)"3S�3�66�A����q�m����=�v�l�(R�7Tz���d�ߧ�SKʴ��$�F��xy@+6��
���w:4��qYAosm� A�
��¾�=�F�Q���Z�I- ^�`<��@;����]�U(IEw��cƻ�~�ʊ��R�ѯ *'���)$RP�E�4sq��g_�z�S,4x��'�/_�������@�ʉy���i��{�"�;�ʢ��cG���27�}��sW�aL�q������
�B�nŤ&��u�����N�,�>u5�x��C�C`-E�OC������o6QY���˘�5\�mob�!I���p�L��=�+P�8k�)B�)u �,GY(󂺘�9G������	s�{��훘�7���l��q.�I6�q}'�����cl��݂�օ�7X��}��&)*�NBas���ns���|��|�����tV���r��R����Đ{n�d��Om�a~1�b��{�A��������4z;���(�����}\E5j�2�2��1U��r���}���K����s�,�8����S��d@|��C>�[��-#�T��;�cۂ�����a����,���:�;1�?p���*ݕ�X'�F�I��R����Қ���)��o���O?#pz���q�3��*�� `!Ɣ�������;v�h bO�R$�o��0�h7���ns��T����ǚկ?I��������VX�a]�q*�sY�����b��,5\�fǽ�w%'czt��4��Z#]��a<�ÐB��°�$�A��1�L��\�*fPQ�AP斲�rT)��y1FZ�HS��[A R���*ٕ�BIN�8����(7n��ڍ���<��󤫤�u���t�qT�
��.y�Q�Y��)q�t��k-�����e��|Nװ��������Fu��Uw��g�j#?>�Os�C�f-f����$x80/-����>�����U�iP�kKJ<���q���5�t��>E�����b ����
�{�F��:=�~��{f��J�E�s�1#�ϑ�(�1A4����B6Q�uT:�����g|������~;�)�@�12D�9��hF�(��!�{C�+O�fƚx��4�1� ����D�w� ��g��-���DG�0*i�P���`���tH$��S��P�DYc(�A
�{�k��i��~�PHr��V�%�<�\�!�e��5�����b����e�-r��!dC�"�!��JJ��I�(-�"�)KK�����P��F@�rZM��?`��͝뗘�
D���Rn���V�����~@o�g�*��OT�޶2�Nz�Q8�Rh�@iA J{���ܨ	��t@�!:ܥlj�nD�u�K7>��:dBPj��a�8Mi4cF6�9��~�oY>q��>�����U������1�0�`w��J���	*ʌB�+<��o�r�wn����ߢ��Ë��3'���O��W��&���r��r���$J�1�_�@	��EK��;@ʋ_e�$͍���R>��k|��7P�.sǎ�ͳ��S��'O�����ǉ�\:���A�ocsU}Ƚ޿��OR�Z�%� ��}���C�����wYZ�V�^��IҼ������V� O
dn(���d��B�bW ������U���hx���A��9��H)��wC�����8a���X�d@j����sz�P��F��&�ҿCń�A�ٴ�/j+��u�UW�K�d������R�A��ڎ?ƉӧXZ�C8�v�Ƒ%)T�xBͦ	�( �b�"#�"�2'MS�9����RE�U�S)k��X�E���ٮB{} 8�&�Aܤ0T�/(ϞV}q��:��y߲�8b��1�#��I�8���줋/5�5�K}X �@i�8@��,%�n�MlZ�mm ��{V`�@E���"�O���S��^�
A���������"���wS��/)H��*~�]
����	�IA�� HO���PVFz
s�ꉞ�4��2瓵�ӓ^rX(oh���Z�vb	�(�fdFN�YZK�x�G���g.���׹���,ʐ8��+�I�Q��g��0���A��sE�4��N��ߟ�����!�Da���}��y������|���&�J�ʚa�t�	��{�+D�:��,l}y�4����:�x��Ͽ�C�}�@�(��� �bYz�A��1�(Q@a	�	<�ve��/�r�������)J�1���+\�����c,�lw�N 9|�Y�#3��F���+kp�ס���C^�<ze}d���A@:%F�h�qJ�m�X|������=s����A��@��@�$��T�������?��� ;�������<O�I��~x����XN�w�f����:Y��)Z)�0�70t�� �ܼõw���-��佄�}��7^����d�($��4�eEXSm�JB����[DNn2��(�Iɨ�HҒ���֡�,��7��\���_Dv�<���9��)�E����w��¯���k�Xh���"��F\9YbR-�_*�ᐂ��<��.ŭM��\��]Af���c_yDb��1�eH|�0�H���Cñ4)��5p�d��ewo�������vC*IPQ�K;ٳ��z߯w�{��L�7�t���[�~���*")BJ�2g/�Aff�<P��P�u�8�PL���)��D�fզ�lL$��s�U�EQ�1�,-,�qg��`�RR����@��O!k]�^?!�cʲd���
�Q�P�-���ʣ.
(�\ �&�c:z���3�^���˽���@����`�'ol�}w��Ӭ>��5�A5�`���Փ0�F�(��݈��wq;%�A��,��(���|���LI��c[�d���K�}N�Hs\�\�T�i�FPk�:O�0�j�r=h�'��^�A��f�$�S�,��B�de��GN�ԦQ
x�9W�����:%��A� 8�#�4���j|_�8���������o
�� (J�vL��1ZaL�����~�:Q����j���!U�h�tH��P��d�N0J�n\���ϱxh�~@��t�VV�ZXD�!�R���e�{��cm�-L1빹��UZQ8������u�e�E^��Pj��� \���z����9���5�^�@8l�"c4HhG]�,�ֹ���ހ��@�6C)	*Y̲,�4����`Q���Aoș�����߱��;ۜY\FHU�F��-K�ސ��l��6��ɨ��_VYuj`,����0�Zh����"1��(-�]�����=�����m6��`��E����:n�5�&���y�"۾ƻ?���^�c���l\c���`0�Y#FROֵ��qH�hJ�:Csq��� ��t��˔�ZZ
�I��`�!c0iF#��~��/
Q�=mj5�ZH�ҞpŔdiA^��Na�F��j7<#e������K/q�kϣ���sor��7�����יo����ׁ�)$�>d��W�"֕H�kZJ)9|�qμ�-�����_?�Q���%e	"1�hd<�헉�K׉�P�e�!��F������=�C���@��X�ua|0��g}��ViÃmtUE'u�8�;R���=gz�6����p�����Ya��짾�N�9J�����hi�XL^x�nj��BNݸ�~|�¿�����Z��Z���&7��"Kr�~q���n:�i�ۨ(����@���0��k�B|�,��"�Ch/���/� Bk��V*O�%=u�qvL�%���p>-�e�����(]�O�{Ů�҇�c�~�8x�ZFLj��:�=���A<�&�����y�b0��D�"�P�\9�Q��Y�ՑI�$%��Yx2�Pi_�dథ!u)Y9&���bń�WX����P�U=��>�<R��08PU.�"'�F���4��p���J��(��i����S���tF��urI���n�tL(MBD# �����O���"���gt�A9C�ea�/֬ #!�yU�3��4Ŧ��!8��_����vi/����ɉ��ԩc���D����mFWnRd�@��!��*GWX�i��%��DT��Ջ�F�F��c�y���u�x�UT3���}�fѥ�a�d�Hpti�ls�s��o��oн�P(-�e��[	�Ä�К1���NQM,��|?����MGN��N٦Hs�\�Lی�oF��{�Y�q%��(��1�QT�3/V�|1��X͔1e}Q�Px�1���s�I�������b����]֊�w^�5�O�$s�C4҂��u������8��.a�υ7~��R�EL4p�oޢ�dE���߸�j����:��\�5�����aV�8���nLjv�!���|�E�V,�7	;]\����0R4� ��3�%���B(� )H���!H�9^*(�lؒ}�3w�i�<��<�$G}�^������_�������ե9��A���I����A���D���Q�����x�=���+�)Cd F8k(R�f�uO=�^X�3J)���utY�m69.�^`ws��#�PV���A��DJ�(xbg-Ri&�cwG����ei�z���;w�=�w�C
������9�ܒ���Le1�*V�m:��Y\�S��Lr5K�+o3��Σ:j�a��TdB��QD�s�ܔ�Β�G|���t�-��>��t:s���W�Oun)��:���cq�;��X�<G�A&v�9O2f��8��Eh��U�=�&f5�gBK�&�`Q���PW-�ιWE������^kb��{C�f����먿8��67)z�~B��a@I�$Ŗ��EVkB%�e����%u%ҁ�Uu���*�d�ԽY&�4�:������c�>'T��n��!�luj���0S��d
)}�ԥ�gy�^J���|����%,���y�/��]�QiQVҍ���HK�Z��p�}�A�����!a�AZ9W>�Q<S���Ĥ�r�_���9I�i�!��9w���8iK�(h���fȮ��F���H�a˂n�"��P�\#B�r�_5�!����$�Ԟ{?+�o�B�m�)�#O%iKHo]���/���[�E�IM����Q���&���>%p�;��y^k-�X��D8BL6���`�2��u������?��s�*��}���{��{��w��C��:�ɲ���h̏�����0��5AQ!(����%e�V���h��B�K�6�����̙�<��C|��C�����d�y��;�]b��ڗ^�n�M�=��(	�4c�g�x ���_��1�؆0I0,SC���)��{wumY�K,w9�?��YE�p �U]�q�ƽ���>�[�7�I�+���w����}@�
�M�]j���������+\.a7Ni����c>���Y̖���xᥗ����%�v�y�U$��c���ů����T�����7�b�*d�H�V �\�fI[Rx����R8K!9�Pĺa4�坻|������`�p���w�_>��� f�}%OW'��9j�����5����fqSJ\��TUܗ����C���7�����맧�X����y��l:���Gf�pX[6�O�1uӖ@n=��3mZ��A���X�9�yw�G��P�uk�e��gm��̌��x�2M$�C�|ȸ��Td�cU�Jk�RZ�Y��C$�R`?�(���r����N^�Rb��R�et�5k�>*E!9:8<�29P
|����v�B�}Du��<TR�"�b�N�j˦�.|1FB,����gL�:Y�
�]1����J#C'H�b��� ]�l.�������/6�r�<ӐK�7�y~6�{�_<����6M9����o�a�EfIT
�!'�����L���<�2c�,�+r�V����3���\���:�-��_�\�ÅP\Ô$�P*�\:���_���ܟ߉�ô��w�D���]�E�xz�����5O�����F�;���V\13FV�UƏ=�%RE��,�,�nV,q�Q�k��/d�����9)�����T	�W51�؅a�,~,f�JK��&�G�ؑOG�A�Lnk'��S��z�r&�Kâ1�T�%��oa��.Nn�H>�o&�TP	@��CV|J21n��������R0�j�@,1�)"�A	�КJ+�wϜ��EG �,f3������G�+W���O�ܗ_`���~����x�*U�%	OGbX��0
/�nv�V)e��k����!�K��я#Y�|n�%i�o�+��Jvx�����1���8�!ƄI��Y!�d.F%���+��ft�1
A������{n+�������7>�y����v�/�5������pcvċ/����1��������lD_�AH�Mj��I%�Q+��5����Gb��>!�P6�p"bo��o��}�3�p�YT|����ջ_������{?�?��o�����_Y��k\��ʒ����2!51Io�­{V�y��.��j��g(��z�/^����#֫V���;N~�6s�p��W��mj��W�� ��o#e)� O��T{N;/������7��b����|�C$A���N�#k���F+I
m$meY65���#r]
'�Q��J�����rb�[K�H�b�6��7[�KS�g�T�'Wb�S�a�MM�q�����C�9�8��1�X,����HO�2*݀B����^)�҄�BB�֍LN�,+    IDATʰR�ĉK7=�6�,�����$R�$3p��l�J���Q�"�B,"er�-qz*
�b�"e�C*c�L&R�DC��X��j9�N%k�Q��c-K�s��4#Q%г�(D�X(���cL���`E���#�h�0��Q�؝B*p.@
�ō#9E*������l��.3��X�Jw�.f�Y�<�\*8u~�&�%�rulWg�Z���P<������t1�Dh]`�I�!�(�O�ЂK�o,o��r���"�,%��(?ga(	���Y��LD��J��{̉чB.K�(�dQ�u5-$1F���$C,$D(]�3Z�Z�	1L1���S+��0�:��g�b$�@d$YMp[=3%�<�x��{�P����#}��)9*�6R�R$E�h$"%t΄�Ok^�^�Ad���n5c�3R��+C���G�i�&9_]W
 &�lJ��#;�
��L�@�@{��Yp�kj-8F:�Q��	2�h-���RD�TF`�BQ�d�.�a�Xo:���!8L��jV4�n��7��������;�����>$��Ȑ3i�3wpS6�I�Х�����A+�����!9r򄍣2!5Yj�8rm�Y��������U^��WpY���w��/����
�a��?��o�#?�������s6���2G�\�cʘ��9]o	!��FdA��3�T�F#SFY�].�]��1
9-�����R�j͓��3n�����ǚ�&D,�'J��I*��Ժt�OU&`X^��Z�d9p?%�~�?|�o��_�n�y��3���s����&$������G����)�޸���)o�����*<|z��/~2r���V Q��U�݆��^�w��F�R���;�,z)ws�I��<O�?q!�FY�@.&����&֛-�IJ-��$Q:�"s�R��*\�W�T/�B�r&dMkZD?���M��K#q!�B٪dM 
whV�Sɟׅ߮�a[Ԕ�Bu�j*|���`1!ˁ��ݴ�
k,�H6��z{��5M�$0M!(Ŀ)I�*�F����Y���舗y����	�P !���R2����dQ�{�[tM��iUJB$���)���@�	k+\��}��iK�<�`�+��B!�%�(39��4U*B	��)�(3w4}@&iA���8R�3m�e�Ѵ���k�y ��S Cq�۱@��Ib�4�&�Lӄ"	l?b�' �0m������<��\.!��J9���\�/-.HqR�ٱP��|��ՊN�Z��Fƀ�-5"�H�i�1Ő%�a��c%Z@�)$:��Ie�A�c�����D��Y��2��X$&KH��}�N�DSѧ����ƴtkE�(4Y#���3�,	1���$&��8���H�R���e���� �����J�V�����1��F+����RItdH}`;�C���ؘ03AkB@�"IC��twuŘH��z��̀-9b�CJ)�����R���E1��%�-O�a{��Ϡd;$��t�|n���7y��^��ɚ�=��T)�>_��]�R�V FX�+,ݺ�X5��0� (y�_ 
)%�:�g��u��+����>�_�"O�f�k��|���TY����w���h��;�q�o���D�܍�\B�|v�}���E���e�zX*���g<x��������5!Ó�3������8��[o�@��A;c���Z��QX�J[�q�ږ���z�iR1��#�莟�Ο��?�9XK;�}�����,�!н�!/�� �贗FM����V���ȹ2Twn��K�����'|���{�x������撧�=�z乥j<~���a5������v6�9�4?�?]qs~�A����w��q�
���C���d�*��Y��hu�B=���Q��?���B��$&_�_R�P�.f�$Yu�.��'J*�12sPW��	B�l�6Iκ-���b���!tם�qrS�]|�e� ���4o���a���B��Q\p���S�0⢘��^�ۦi�r���~���w�y����Ѷ-z�ïU͎�|�K)"o�6z�-�v�ߤh�j����B�¤"d��0�r���Y�:"����iIƑ�%��#��0A�)k�X:�=\2�ݦ��IY"�-�k)H���l5�(��JwJ��G������!9[}Z��9�P$�l���iC93�.����X�]z��)�T"���<�y�����r�Τ��&�k�K���d�"��OJ�ֈ$��c ň�g[ӏ1GF��"#� "IfP����)�C D_�T��4�'�x�5+��� 1�&e�J�
q��'���B����@���U�D�&���E�\�ݔ,�H�Ӏ�j?#T��QΤ�	>��3���*������@&O�T!�d�l�
?c̎U?�t� jŬ��ĎʔB��Rrf�	�)��M�v,d$i2����6Ƒ��h�`���*�6��(����+Z֜T�����5��D2�݌��Q���r�o���s����a�Eݹ�o�@�-}��-u#�>�����w��g�*%�� �VȢɎ�at8W�7Z�b�{���/�̗��:��!=�_����U:��D�g���D�������Ot?����+���0hm�1�c@�Dm��|Q�.����j���1C���@5��]G<M�`(ZfQ�\?:d�=F��(
�zt�U爱��r��_2�k-�mW<�ɏ���c��3�0�u�ȴ�$-Aeb���F��ظP�Q;���w����s�^��w�w_��u�����{\'���p���e�(ҵ/FN>`��k��{os��S��!0;\��5ܚY6ܾu������ ��㆖x�s6�1on~��"��Ŕ��g��x�c���+�����EW��������a�.�.r�{|R��&��w���,mME��DE���s�:�b	.."����`�]�/ͯ/�B\~�6�ݿ�^7Ʋ�H�+$:)UY3��FXirY���pyDƃ]Y���#�r�LR9!vc�B ��r��/L�'����$E��Q�~]��"!�HXk,�jB#�����ad�>�'!e�i�p��QMU� �rp!N�6ʅ��Bb5��1:Gm%�*3���H�@MUzv�4�mΊ�p�E�#!eJђ3y�̈́d'�(���}�0�֠2Xa�DM��d���!E�CT;G�#"���)�l�K(t.@J��]�w5A���qt@�6�$��s��9<Zr��N�7�i3-֌JJL;é6g��(�0B�e�0�%Y�)� �w�q$	m,��"���l��ӵ�L���i��0�Heĥ�$**S����d��C��552�s(!�m5Y'VcI���V,[��l�Gf��9bU�w %J)�S��ԍa�
�R$��&u�T8	A+R�H�0HEv$���i3���O�1�����/��UVX;��r�(K	>�����!� ����9�/q�������>�s;������"�#m���H����?&��ES�����h����pB|ʄ�
�I������
Fǣ����7s�}�u̬��ZTS�$$A��[�køb��C�.=c����*D'���T�PTZPk�׊m�V��g�(-88��\A��%�����B
�uU�ʔ�bB�;O?�1�6�=	���A9g6
tH�9lʼ5��UE�qB�ʚ�bm��*ֱ8#���1�;Fe���h_h���ȏOm��,k�,�b
�^�9=a���Wy��U��9�ɊP+�چ�T�zɲ�����Cf����B��ß3��U�z?r��M���Y����I)?�:}�h��f������r)���g)�(8��K�{�im�����$ŕFshC�*͙����랡ZpX7�	]SU�Ǜ�Sc'��}���ra�SqĤ���䫪8ؕ�gI��k��jG�fUU)�P���#;T�|�����\=:�s��'�KN�/P���wW$��D��������_6��+E��B��$^�=O�S��54����$��=>��t�*H��~'-���9�=��%�4%L)��R��d!I9��7��B��t-
\��FP�%&$R߳uO�Y�'��L5m�i��KF)�,?��r�t6&H9�Șv�y���f���.�ː����Eۮ�.�߬Jk*�A��rNE�#1l-qc ��( J���kܸu�7n�9ߒ�Sw]��t�(��6�K
;k���� �,�C'#����4 D.�gJB�|�~
RH$B.L�������q��PC$�}����d��h1�ms&�ȿ��L�:����>1�7,�Ī�q�F���i,Ѯ��_��2N{GҒ�G�5-7ma�Z_����Aj��֢�Gb�Xk/ �1�黛�9G������l1g��t]G����1�|�G���i�3�c�$mPB�住����r��X ��;�Œx�XՄ(qkǙL�9�>ꩣ�+���I��EI��!�;?9�	�4����99�������ӿ�O����Bl����	j���R� 5M�I#��	r�FTG�@��y�t���rH)h*�5%"���3�J8M�D9Q�B���(3��
�ue���G��U�d�)f+�H?f����1�����Iu5#��$"q*���@j��auE�d)޳�dm86,�9��ҁQf�M�R�[�֌f�qC<?es�Ó�Q�S��s;�ɒ#٢r����/��i��`I�4(:��� g���F�Rs��-���:7p�s���Y1] K�Q�	��Tߝ����sųd�39�-Z2�I�񙭃m]�dc����G�:�����H�=�}`��-�aZ�;�B��n=U6zb�_�/[c�못P������ϸv�MӔ�����~�(�u�_OUUM�
� <�)k�r�`ִ�����1�ْ�þALb�#T��|hU�K�=u���R)ĆM�"�y3#V5J%Dn��)C4�b��^m��'F�/�8]1\T[1F�tTA��V
���|�sl�-1�@�VJr�I	lm��n�8F"��uJAul��Y��t�K6h��FԚ!�bèT���q��ΰFJ��^��QP��2�9�r�,! ��o��yKʸp3�2��,��3�v�u���cNO?E�@%�� Lq�ZH{��,��֨T*�S�;��	��(G���4�P�!oe�j���v<+Y
̔g��q�͍ �d�:�ڵk��P�jj��5�s1��l6���72E�"���"/�Q���s�޹�ʂͣGD�P7�c�d�� 6mN�bq2:²�.�ē3�_�EB��;�'��`̑ӳ5#����ɔ��R�K�.7����k�!1m�RQ������RbM�kH)��
I�g}`�(�pU޿��~��p`�or�:V�S\gT�����t����b9�p��/ŉ48��HH�81���r�w9L�RND�T� �����kt���s�{��,2&g�C�p9�t�y�mUII
��V�̍Q�u������� 2$���vל*c�JMHKd6�h�A�T��ڶ؇��gt��'��=�e=xYH��9g�X>��"A�T�XP$D(ֵ��!H�ڴ�n,�U�.�k�9G����)�
%�ZAآE�X�r�!�O�+A�`���YC�$�8��Q`{�L��,T�D���3kg*3��b�0[.����s$/H�����.V�=�jw>��Iw��gI��T�_z�3�r�����1r�kC(^fʋo�����k�4t�1�mE��X�<e�G����&	�s����½�t]�8��D��X���=}�G|JS�[�5km����,�m[n߾͛��oQi��Dh.�E{Bد!������q%�秤hj���yy>;kd��]*�C�/�/`�]g��H�.mq�!�27��«;xz����Uڗ_��7��_A�	�@$ -E2�\B �R5�.�a�%��3E��#���ZT�1�����Y���T��ҚU��w�����b�]aMN��>z��,X�MS�pJ��� 
.�]w�I���BT�0n`�$M�N1 7D�/̀�V	f�|G&AV�v#���r��7����l�,�3�4�����خ;�����;E�#9E�H��0Rq��)n zȁ!x���W%6�����Q��w��Z�ιj$Q��^dd]��'O=N�����y��I�Њ�V(=E~�r㮤d;����gl����Gв�N]w�V�6=�T,>�
/��7��_Ɵ������c^������Mݿχ?�'�|�ELܹq��醃/�ʵ;w8}��O�G�4��Ј	��}`��{bdI^H�vs�]�=�q�%��Md���'!�X����\���1I�s:���զ��#s[#���mB���m%�<E��Q����cR����H&��R����.���8�M~�,�i��N�B
�FI*�ʼy�����HzguZ��G/���p����D6�(Q:�:+Ѧ̋��8��H̉,�d�H)�c,$:����
I�V[B����R�#���SĥL�˽��ĥ����ج`'�M�!�DX	"�ܚ)�%���b($ڔ	�����S����I�>B����hd�0R�Ǟ�w�2AV��!�J$0ɼj0�19�K�uG?th�WB�]���}��n\���
�GO���͝�(9���r�	Ռ�U]B7�=��r1�+���M�^��w3����WB2���V.��H���0Ҙ̕�%�3��nq]h�T8�C�O	i+�1E������n�a����n�'i�L�XxMJ���i̴I۩h6����	Z*�nSb��!N�2�w��wE)���am��ӳ�Qԕ���1�M�V5~�elx�����\鹱�xv��x|�� L�)R�r� ��V�n���^��W��=�Ijd��"BLH�Ѧ�	Η=nGR(Z�#�c��緖�����g�>Ĉ���|��o���_cn��d�E��ҙ��1�Ƒ0�N%�.��N)ML�¢,6�%�n�o���6�U���O��o������H֗�C�4���
�̇�\��wZ�b�CU��P�#N�]��)Y���o�&��~�=<����]n��7Xg�uCV��T:ʄ0kkH�quL�0v��ʆ���*��'lWk*��)s��	9�~�|���[%�1K�rFu�:/�E�:��Wzr{J)�=�����y�>��:�Y�l6��l7=OOO�x5��79::�]�hD�4���ܻw�`Ŧ8��K��G��;�+���5_�r��G����~���SGWy���w��m�������(C]K$�a[e��9�:�>�Aj��`0�&�Qd�Z\�'���'eEYԔ�h[Ў��ϸv����0l��"jS�5l�rݥK����9�n�G�=w����P�b.���6G�	2��5K���ȶ�%���q��q}�H���L��KeY�{V��.��11�B�U
�Vl��3V��W�J3��_�.�6���O�X����ՠ�4/�jN҆s�(wQhlJ���
���j�KTg����Uj�VDJE�iKll%�g�41��1N&TI`��y2���Q�H!��c	���V�J�v�{�Y�5�J+r�$H	�.��uVEI3sU��>�F61zre
�d$Zj��l�������,�F�ud��k�L�B�7GR�jK�,f�n���!C,꩔��P��\8Q��w��gm�ϣP��y��w�%/͐�D���!D��l�.
�*��J'��̬ 7ҭWhӠm�j3�8l|.2�I�L��$�����:�S뤔��*��;����햜�>�&��R9_��t[>x�C����I��zOГR�B>Fb�{d 
ϣmfHi���Ɓ�����^���vI�e���cB���_*��M�	c��[dR$�A���(����z��5�rN��=~�[�:��.i+�r���RJt��9�tԪ��v�z6x�aK��)iK�]@�!�z/ٮ7��rG�sU����Ր0���B��w�+���,g��5!G�UX��T�ȍ�����,�$`C�z.���/��q��1~�X$�Fa&�$�Hm$ەG�~��K����QÀ���%����5��K<��1s� �'9F�,&E*&|�c�͐B���֫_g��װ����ػN��,��Y�Vl��.f�W��>;�`>�	{3j    IDATu=���-�ӳ�Sq���g�l|���>����i������D�(YKE��+�����zq��M8�n2���1R��d,Qk��
��9䬦>\r��po���m����7,ԂF^}�?�����|������淹�[��6���_������������[�����;��ᣏ8��� ?@�����O��ֵ��n���[��t���s�$�J�r.�-�e�e��Š@�p;�ZAJ��״�X�63=:q��;��F�9_!UF���O�1�/
���愄4�y��ggkfU�t$�b��\!�.�����ŵ��b	�ul� Aa��/��C'�E�!'i�B�D��u�0����f�P9��2 ���9�	1`?�SSr�,��4�����������Ĭ n�IJ!+���1�Q"��׆$uA�6�$�C �J��!�Dt����I����J#��䨓Eg��.%z�s�6�-]ױHg���A�|��IV�kŕ�0�9�COp�#e�!2��O�bŪ5+J��D�@3gq�$S��d��s�1t�����Ҋ6xfVё����iD�D5�|O���/Q����#3�cS d���('u���)&�q�\�v]..����/m>;�%`KH˘"[?��TJ�r($e+�Yk�>'�^�t�e���@�f||J�\Gd�P���(�J�P��$�� ":M�_	R�)����S,Ȝs�����0a�Fr̴�Ň��V(,$�@��G�ĬV*�h�G�
�M!�*�͉@��D&�h֚���Ź��@����c!渉�DBN
,+T1�J�U�����ů$%�\��v��=�2Id���F��W�7o�Cw�>���_2~���蒠��R��܀n[��+b�v�8tH]_�0�}bfk\��j��DK�=zx���	� a8�<�?�1���zA�[����*xNW��#��!"��].sDǢ�����b���u]s.&7�F��_|��撴)�H�%L�9ѐ���	����o}�7���<��}������ܞ�$�����y�Y��X-q�-"F�)��,A�c���8߮�砮���������c|_��BU��,���g+��1>����h�y"]v�1��w&��+>�tTʰ��@c$�c���1��mѪ�_�'Oy�O�8";�3[��Fr¹�����dF�LU��'��UQs�7o���|Ƽ���`I�P�V+������w燜�c^~�s�Ê��S�{�|��G�=z_������Ïx�ͯ�	ϡ�4�o����h]b*�pR���Ѥ,َYL>�J�t����k���~��W�L�Dܮ��L�� Ǳ���ٚ���Fi���P�K��՚\����HQ��s�gH���R �X��:��Ĝ�)�%��s^��wA��?�Nk/��5��ۋ���L�ϥ�^��`;��9�d�[�Q'�Ɯȹ�EW�9O���C0�e>I!i-�z�rV�&Dp>�B�I)�ρ��)RUئfk�*��2�<�[zi+��@u�T&$���Z��d��q�$���'��l�ӫ�J�7�����@����R+j�0����>
9����H��t�X�$#�d�HH����	vV!��۞8*N��9s9��#��UE�e�L�|$ň��ܘU\�tl�"E�L���Kc^q�A��_g~�z�M�]�z���j�H�

��ē�B�#�s8����i�2�hjB۔�KD�uM�z?6���ER�u�G����w	7��/����E.J��޲v�䭡�2Jc9
B��#�i��%	�8x�s�J����1[�k}G��#�)�З,zw�G.�~�µ���)�u�S|-��B����.z�(�&�p�f>Uw������ӷ�°��Ǎ��}�m,і�[Ӈ����~�1��ᦃ�(�����=�py�q�ѻs꘩��27�H��Ǭ?��1fr�X[#�l�2���,YU��+���<����CLž0zje��Zd���h [^��?��[_Ǫb�`E�BJ>y��ǿ�W���Hcd�$��+p���|�7dbX.��ڗx����ݿ�s6����o����������޻�	F��|^���0`�5���{|���t�lm�051$ڶeq�f9���W�~�JI��9�|�Ï?��V�q���V�fp#^dbؐa;��Bk���G6�|��{Ȧ���L*\$J̧�E�PU�łs�Y�@����`qȫ7op�d�$��	"�r���m8��y�2�C!�F��bk�z��w~�S���~�s��)���7��_��'��+�G�plj=J�$p#�T�R"U��#c���w^��m^��3A�Or���w/���;�g)��CrvcǑ��đ���d#�Lte���,x7�R��!�RX�����Lz�P�(��녌!�ˉ���x7�)K�\��i�ķ��ȧM{�'�K��#SC /���ʜї���؏δV�� #���1��,RNS�Qr&3uJ��W�������1��zU���l4�Wq��YY������Q1�GW�m���lV[�.���p뎏��c�ˆ���r��U�rI�,k!	�-�4�ꖁ5q,�BNs��LC-�o�|���1�(n�1�p��{Ϩ$1�x;����D�B/��䜘�Fk�.⇁Y���>�2#�J���%�VT��n�kE'4>+�������}'~	ʿ���&����30�t%q��#�1)3!�$ˍ�t.һD���H���,+C5�t��L%�d���F&�}���]8Q�q?Y��F�~��#_H�
���94��H1"rħ�)�jhꚣ�#NNNǱ��TQ[��j���r��'!!(Q#%���9sي�W���/�1����fF�NMR*)J�i�	�JU-Dhg5�L4:�֊�ʒ���'���?�I�x�a{rJ)��z�p���c�zÒ_9� :���9}��m+����v��I�y�5g�����T�B�l��s��xGGב�`��"q��;�s���4C��o7$%p��w��GO����)��jMΉ�m���9��"�|�wH͌q���7�{�X�o�.�(�_��o~��?<���ÿ瓿�?C�H�JB[ʩ��tqĈҭlG�:�\1�{��x�I�-]�S�}�����Ɨ��9�z���oNs*��v�k���ǟ�����#�*�O�Q��Я7�l�NL���!{Ҡbf<[!��<�l��G6>@�"l�I
�{���k/��/�t�������R�@{�7�2Z8�#��?���x�+�GK�\�C�*y *K☹z�*Fh�jA[-y��	��>cv�>�Φ����vRv�"_=HS\�|!-�L��c�=�$��3��1צ�,�վ{� 3 $�Kr� �JZ-d?P+�k�FE�\)$-�� wC4 8���fڕɪt���fVus@�FtTwVvE�5���>�Ͼ�L���R
ш���J��9N��#� cQ�C��
΢u�������q�h8�`�]!nd��n"<���s��Ń+Q2ڋ�څ���ĸ��eL,��v^�b N\p}��N�ݴ������b��_6���	���?h����}�2�\�ȔGnd~�zR��|tY"B�RƴI����$��z�j�s�u�P5!S����4����o���r�C��ߵ䉦�W<{�9��AIӵ�C���Y�Vŀz]��]W�4tfŝ����C�
�^c��8�����IQbV��h���1L
�?{L+��]9@%,��������G�߾� J	g�m[㼡ԊNKt>�A6��G�9����@o6*�	I���4�K�iPX��FL�¯��f3����"7�K��f�|���k|�\��=q���}�%R"h% x��X!h4>`�(��6J�Ge��������|��Q�ŘWKoL���_�
�!b�|3�B����2���x�RI�:8���^{���1O�<�����lF]UQ�#{K^I��8�5EQ@�1Q����qz�/\�����%o��s}�A��_��q�p��z^� ��zZVJ|E�R4����ѝ�ҩ���!xڮ$�*Y�N�>g��	'GG�J�导˭W^#Ï��?���O9�9��;$ݚU[c��{��g��R亟')�uגܸʯ��%�䣏9}~������ W�87T�D�1�щ����T���s�����1�
%-��0��1��3�G�޸M�!�Y�@L��C���y8?������'<�!�%��h�w&j��B8O**ҵ+�s�EJ:��Z"�������ȹz�+L��u���Erp@K:����Q*#�	*����ϗ���;��G�f3l��Y�Y6k�D�B�it�V��Re�=�TT��rB��W�s�>�Yv-]p���_��NGȤ ����x�p������������s�v���\�ݺ���D��9�+��y����YB+w��5�'Oy����_?�L�mI��EI`�����s�2��лH摒�D�mR�0�7�ظ��O�%�\~��9�P:Jl��b!�D p��"Kw3��ć�I��,�<�H@ے{�,�L�|�x�LN�>S��� 	p!����P���_f�<������yM���D�o�)8�良����l�J��ד�-�z�����]g,��t6:v
.d�҃;��u(GHP!&�)��r�Z���$N��Q�#����5u��Δ�ٌ��?��_'�D�v�6�;Au��Jlԕa�{�ns��-vG{������}�߼A�j��A+���9çG�M���}�?�-�	eȋL,>Q�F����r��������PZ��>	sk�I�s����?��K�2��g���)� ���j���!}�Ø�/��_��������H�7�7�Q�}��X!�|�nB^��Q����0��ES#eN�4ț!Bډ��:�H�TѡS��JFk���U*�:O�)�z5Mך-9/I���k�,Q I�fgg�7n %\	W988��쌧OSU]��z�$��qk" �ĸ@�6��ۘ��1��2ʴ��I!�C�o6v��\:�[��Z�n��Й�1t>@��*��f���"(E��,��DY,+��9*bXG��|H�V���,y��\�'�wVqr~�mb����#>:��_�U�r�C�^
�"�i��&�@j�>J�m#��[_!;x�jx�5'�+�F������Zd^\&��&�Q�-�<x�]�U�2?;�^W�i�c�k>������w����wX�/�[K�ȇ���������;�Ja�w����4��:�	��x�N���Y���4m�J%$J����p��78�}�����:g;���	-��:�yN|�P,w��>�<<;&�v�_��_�5k�<�G;�1{����)	AK�w2n�s�T�*�Dz�]�c����[_�ؽ��|����9��iN�,g�#EJ���m�x:f��jw���e}~FW&�V1���Q���Ԓ�t<���o����Mn�T"M��2g��k�-��b��y������⤉�(�!��a�'H��.:d�ύ��H��&.�}���Z�F_ؚ�Џb#*B@8�z\!i�a���lI�Kj��e\�;s�l@�~sF��l���:�q-4R��;�N��o���4��7�7v	�MN��MYnX��E3�/�Q���ݼ���'����g��7�@��;���v��.�ERB"c�d����q�fX�uCg<R%dRж-�R[��(� GS*~��!V'$YB�Dr���j�lv��mjX-��Rq~t��ǟs0��Vu�����)�����������Th�u�����>�D�*�Vh�1G'��+���l���>�2-',f�q�o;�4M
�rH���I2`/�`-�Z��d��)IZ���&�Eu���>lkg8����������r����?�?��X?����@tf��˗���g�>�/��C�|��`}qIw'����zƿ�D?N	�=�(������DH���K�������ڦ�PJ!]$=ot�I�`���K�����7���	Zm�sƘ~~N϶��`�e�\����Z�8�?�Ν;�?=������ӈHh���
A]x�8���u[m�R
aE��
�:����Z똴���އ^�i���9������e��!��Y�	2$�*�q�h:a�ޣZ��gOi~�#���.���06��ڞ�(t�������dq��|���bQU<y������ck��h-Awk�B�=�k�T�H�������Op�0LS��wx��	O�c��1i&�&G�g��4�u�UC�4��"��\�D��R�#�U��{?F%%iPdw���㪔ݝ���<����Bjj�L�����R��j�Z�$�$H�m֜�����\�Myp���Ag�匽vɧ���v깶��b%(��'M��L@��2͙�����6��)�����o�`�7L�u�>�H�B7*��g+K)��W��1��l!0m��zE�v,�KƋ=D�1~�.�ȳ�3fu����:*a2؋��5���Gh2��˿��ׯ�g����ԍ+�7� ������2��G��ZoC�w���8&���E����!HN	��C%q� 8�w�BA/;��Q�__�h�k���IS��-r��0_H���X	��]�t�6x�W�K�H���yߛ� tw��:�7� z�zm{�����*ba���B�9�p�f�,���b>E��_�) �����k!{���*:�O��$Z�kA�dϥptR��s4���zo})e��p�/�+7ؽq�$�<��S���݇�ՂNAe;�uC�Rvvv�C�X@Ӓ��9J4��ȳ�u2�4����N�5W�c��u���NEJW-9��C>8>�^��+%���%Uע�F�42��[�'W)I���!Zkf͐+�!�A�\��׹�����3��g�񧱋Mt��Mz���<��|�ߣo��/ �KFb�C���$J��J�К�L��,O�Yp��p)c��>>�����1NZ����m��q]�T̵���D\�ɣT4D��e���罘H63��/>O�Gn�Cq�u=Y�C�Nb�!UC�:>�JEr�G�8??���۔e��ի��Y^����;�<�I����E���g��m�5R��&�x
�������ySh�K���ͣ�e?�cDd��PY�h�ɕ+8�X�V�EFX4Py�Z|��C��a�%���{�*0���t\2ݟ�^W<�����jv����'��B��ќ�2'tgH�!����F*v$m�a�CY��\ �;n����$���Cr�C]�4����Yt��!|`<S�n988@�ğ���B���K*5cze�z~��?�#H;^�����S8m��Ss����8[u$*�Z���� *ʋ\��
MJӮq�f������hĪȮ���FS��{̳�ⷿ�M2鑢$�u�@����'<=9C.,�K��w��OO ȤC���(�3KBg�u�@*)�S�I��h���J��y�����{�'�y�s}���T��%6OH�� |Բv�Qâd�q���љ���d��J9�|�w�O��)�[S�Y���1���u�Wnѵ����!˟���L1*�6Z��ޫ����:j����,��BćT Y�����s�&Э���9��3�7{ }���8`�p�ek?/W:A�1�FR���_��h����!f�[�0NF�B$H��QMa�ޜHm��7���#b�BiR2�±��P�L����φܞ�-��Ҋ����.��������Y���è�b��1�YkA�h%�D�U���b��P�hM�-i�g\�V5hER(�̱?��LN�Y���7n3y�&��ǋ*ːR��)�o�J5������#Ui4�)$W_���;7y��'�?���u,��/���n���(��"�g\� !�3C�(|�b���+��e�J4*O@@kMX������)��gώp*et�&A��/Rv����o�6v���v]��V�T*�4e��*�]�����?@�#vPL'ט?�ϤxqS�x��"�����"��k���
%���E�؏���
�Hb�k�<^꺢��
Gۓ���$a���[ �m�s��8��^����D    IDAT<Z_w]!Jg��1������I}�3��k�iI��?}���lF�4�F#^y����%;�1�����Ni�(U�H�Խ�C��A�>�9t���홭��>l+�
�m���""���@{,�jT��8�\��
�������Ue,�BVd�!_Xt:�њ$(�����W8]4��ɧ\�q�~��������sV�*�"I!I x�<Ek���s,`�@zS��T4��Q��E���ZB�5N8n��f]�H\���S֝��[orvt��dēG)�����6J���R��OF�'��6`�@*��Q��3��4W�1�B�|��J$�ŷ'L_{������R�"t���xM�Ƥ�M�(~N���W�']���K?�ӂ�׈<�-W<9~��w�B-+~�!x~�׾���Fl	�}��혟����{�<�pk�%p֜�IE^0]�k|�1^�H��@�%K�6�iC@.AS�v����$'/}�i$�|�5LW1�"0?�!�G����S)|�gKλ�GWC4+�i�$�<C��yb��4���C���O��}��q`�Λ���/r�;�x�h]�Ĕ<�P�����!�K�Ҥ�iޓ�oݸś�hG�Ο�((��0������s,�N U�W�<V�(��u��Z`�� ����"����tV2��m�y�����{�E��P���@�e���C�%��:J�����)�M4A�ƣ=4�S�;� |�N#�������jG,� ��-t��#O7���"�na�`QA�!'�����á�G
C!��������!�<^V�&0��g%Z��&m@�ڮ%ђa����$����N4K
��:��ٯ�x�����&t�Q.�4������������K��tM���h��S��V��4C4�� x��<�*�2��d�!+B)��7ܼ�MS��C#(��:tq�)Q*�u��m@i�ܹ��B������l���>�tz���p�$k�҄� �7"�zvB' �,��_fpm�:�zE^���/qgC]2�`nVv��
=L1vM)���\�HR�/�~� ����D�
��5�C���!*:���!P��Ĵt�P�ܽ�.��8P��'�	��ĸj�m�a�,�ƒh���a��\V4֒H$�j��&JY5*Mi{���cm]2�P/*\0��HLcX-+�fs�=?��իL�SƓ]����NO�9;�Q��x�����T�:�#�4��ȕ �i;4���������Y�	m3#I<�4v#} ��|��� -4���Xw5V+�.���)������u���O����3l9 �vI\��G��Nȕg<�����',�(Ah[l�-"�2&�)u]ӵ�[���M�Bo*@/�Р$2�	�l�:�s�ܽ�����ë7��qr���O�ҭ�@ݵ��ϘUG$*0؟@����pB��H�f��ŊG�T'y�k�����>���Z�w2!�����[ "�(�KV�(	������LG|:�C��h-q��K9(XW�������;ܽ{�����8��d9M[a��q6��ak0�oCZ�$C��x�'hm�~�&�zU�5$YF9Ȑ:���HR��MI�d]W�=}Ơ0�)�y����"�
��� ������[����͝/��;S����w���xx����H���+���_z�����9Wv�N}#��6݇�X����+N� �������x�W�%��9v݀XcHC\�6�ᣳd@nO�!I��HilΒ��~V�l�H�q��K�r�����%$B[�A��h+��y���؁Y@�:3| ��D������^�xf��y92v��Z�V(�P�m�{#���j�=�l�g��_�d����p�U"��$��R	�KV՚R%Ԧ�s��()z�CL�4MC�&H�1m�m;������k&R����|v�cN��o���i���j:����|�i�AA�(����쌏�本�Z�zY��N(�<�۽�Y�5�}N\':�*IM�Ԋ�y>~ĸ,���T�+$�NH��qY�9Kk:oP�i> �c���bZ��DC���!�#��o�k�r���{�իW����ɭW���WHL���gsv�.�E��C� �`�m��w%5��lV��$�	����؅��Op��$*c<(cA�"��X�Nu�+���R	���:�{�[�	i�7�yJ�jY�V�et���v1a4r?�Ϡ$Jh���y�p8D�����^�㈸�᫪�Z�r�d�\�3�pxx���>��c;�?�Ç�����v6�Y�BX�p���#�e1���8��$�xHr]M,���
�bH����r�<g�`��tB��lPp��6��m��Wx}����L�|���4MC�bPF�����,�� ������H���p��".΃�4��Od�fy�b����g�Z�d�|<�zy� ����,%�4#(�-<�(�r�.�eA]� ��+�2��E�j}���{���O	:#_/ѹ�4(��!�Yb��9,��}�HM/�G�0.P5Y�F�#Q����[�mi�<�v'����tFq2��:��rȬȑR0ݟ�')ղE H˒`]�KC��[a#SW��]!��U �-2Dݴ�,�q6���p��`�%EQ�&9Y����G���*a�"�f�É�/K�m����_�w�[�rr�'�m���`��e�W��8�����ۈ���k轝��)��ܐӢn;��;vX�����Rj�v��Ϙ�S+���������C<�,(Hl/%ęwo��g��'�G(>�$Bh2������k��#(A4�JP2j��,[��qT�M�m�!E&D�i;�ÎB"c�҄��u���E�s�k��/�۔L����Y�J�&���وa$}"��Aq�8�\l�ó����D9IdW� *���tԝ'�:�Ka��n�B��9BI�T�)�qqq.��2����ږ\	�"�ZЬ�H�6B����ppm�������:���m�|>'Is�"g_g�r���S��<O�Y�>�h�RI�p+D�pـu�^��+��r�K|W�U+�<y�d4&�� �`�T4�.º�r���v�l�D���(�@�F��	L���dt�u���{�w��_�*n�9��G4�?��w������ii�X�~���;���A��	���-q6��m�/��[�9�6������^����������2�Q"���c\~�
��d��gC?��s*��ۥ�V�����<�zm}L��@����M����|��d��:���`Jp��U����7���YC]הeI���)�x`vzF���9l�<10MIM��c����ی.?c?��v���	�P�^G��x΍'sųc��Ox��Mʲ���Y�hgʻ�⛜�%v��k�zI�^Rd1	�|�`�Zm?�Jc�+:�N�������O���P!{�"�ˌ��[},I�D��4M)�u���'+
����z����W�`�&�e����*k;��I�ȋ7o�`~�OxrN��<{[���!W�=)�o֜��4u�4��;�����9�?����5���h+7���E��.�#:�
	��
L$t�$�Q��kki��;�y�z�f�ZB�OL�`P��X�bA%�$���^ܨx�->J�D����8��¼��!(t��e��:��^����Di��1�s��o�����g�`1�cl�1m$_%	j�0����W��dz�������;�o����[�@����:���t�`ox�k7_�Y��6�qz1\�OzW��r��Y�"�PK��dL�HZ�P��>?��l�@I��z��LIZ�bh����{���'B��W5i����h��Ŕ
���Q*��u�h���T'tkKY��U��Ԥ� D���C���� ��H6M�:�s/�H��i�'��(�3����и6Ʈ�˲��������c������&pi��f�B �En�N$�[��ZH���(MT"��-]�3�(Q�6й*��f%kgX5�f�C5_�����/h�%�U��
3	Hߑ�Y�\o�hR�鐻����kWIR�����3;>a6;AȄ�������[??�ѽ�y�яiϟ�3�XS���EJ͆��B 5^�]���/q���iۚ����Yq��+���;�`����?a�\P�KYT�,OLx���Q�H%"�xi�R"�scuG~p��o�a�r���r�?�	����W�ڷ�߾ŕ�ަ��UN<!	�L-&��C�^"�]�z��/?���lP��؇B�g���Jҵ_0����-k]k�^,���V�o��~kV#D��n�)�"z��D�Bl8˲dg�GQd�U����#/�����/D\/�K�1�y���?;;����>��sNOO��[y��{�� /־X���~M�'8�r��|4��B`��n,���d�V�p������w��1����̺����zMk�ۀm$�T+�g5E�Uuۂ1gY��۪g�Z��R(����՜���RZo�dD�)z!lC&;;XkYUK���������`4���ո�v�9l��9�(dd�e�n�Ÿ��d�lF$>f��$�x�c��s�A��\`����S�_���~��X��!cS��.�"�%p�8�W�F%	i9 )rd�P�'���u�#
���n�"t��l�^�����1����s���f��]8/���Zd}QY�P�\�#)G���l���9k)1MK�W����`��]@L��&v�>�g��$h�l��O?���?}��<�{�|��֛_Cc��
)2J��?�G䊰��������g�{lX��OA)ɺmHx�p�X2� 9Z6Ь���4A��i+B� ~���Y�|o|#R��	��>��u�P;G+%�mHw;;�D�L�lU!&|�R79A�Ԛ�YSe9���
��[K�Z�M���x=����vX�X��P(��`��ٌ�����Q#�
�2}��8��4 �l�v)Pb����r��d_�sq�\dOG$&.΂��Uc�=i���{#n\٥�,ճgԵa7��L �	"� ��]5%�E��,�w=�E�RJ��ƨa�`8���[y�j���?��Œ����k�{?�)��?d�:�Ie���D�%����F��X9�j:��{���8>>fP���/�"w޺E�eL�%q�r|��3�j����J�{9� �^���aݮh��U�a��A�K�g����r����YÇ�����Ox#mx���`o�w^���SOE����MDs�'�Q��E�����gm�/y��z6D��{6�r�H|c	ΐ���!��G�/��ݿ<J�q�Eg-"�8f,
�T4��vf�sق��8����{!DDv�$�8�%o���ɐǏ�8::b�\n	u����}D� /RlgX�V��Ӛ$�1��D�2�3&�߉����y���%qV�X}��;�p�5��w��LR�)�y���S	���WI���iJ(Lې�9�h⟈t;��TW�����ѥ�� r#��"���O��FU7����\.��PP-%M�!d�zݱԊ$Q�t@��U�0�ƴ��X��x�#	�k�.���Li�崪8%R)�ŀ6hN�����`XH��G2����Mٚ����}�v�P�$�4C����:��c�\ѭd�rr�i���x�p�aю�%���J阬����!ײ7��	������$�	�o�M�����3T�
�-i���j�D���zIR���	4M�
��yB�?k<z�ӵ�nI��,�8�{�������\��?����x�f]���dO��ѩ��ᇍ��Yx��b�'ѐ*��:���T��E��b#�����P�ؼG
�dw�:rwJ�4����i�E'�����B,�tuG��h���#�,i���G<yxJ����;��������Y/�`p�r:dqzF��	u��8��c���K�by|Dw��D�d���d<�:���+
�uMB:�!��舼�>���)o�|�-�v1����*�-y;�ܠ"���O�u�}�� �΍�\������sD��D�e׹n�H�T�Q���9��>E��5R�(ٕQ�`]�jY�M�2�L���e2�X�w�����������0$TmEil��]�����Ga��w���j�u<{v��~��ځA�@��4ֱ\��sf�3��h�S���1]�f)~2d�3��4�W9���h���O��Wػz;��ךE��n;�͇�A��#�]�RA�X�n�V���~�,������/+A�xhl�K�n��|�bց�ӭ�MՓ���:�yOJ��2f@!(�r�_�p��^*���]�HӴ�e ����|F�i�N�Y.����C��E���s�ޜ.�s�e� -b�\R����J$�$Jh�[Y���8��C� �!DH�uH�$��aB6(�yA�{�wnRO:,H����z9@MƜ��d�\�v5E=��ΐf�$�����i����~�Ρu�s9�6!��(u]#��:�"�(�s)mס���h�u�Ã+Y��$Mh���i"�kP`�����j���=����1+�Q�x�D�ܪ���ءKI�=2��i�����$���1�,'���Mן������*KQY�N�{�,��q3\W�m�Z�e�q�I�L<�y��YJ���}B�F�!���K:��H��ΐ(M*3�v@,�$�EM��v�Ld�U�D�E$G6uM�
���4uͰ(�4��ij��A��긳�p"8O�S�ֳ��Eҋ
��5�l�ɽ��-���_}�ӣ'��O���)&�7~������r�:3��!Y:"�+\t	�"v�P�|l^}ǟ$��TX��rT�ڎA���(�s�"4ޛ����z�H���f�:O9oi�
/]�u���&,e�Y�@'���,�4�Fh�����������c�@'Nq��C��?���/�����_�=?��?�N��ʷ���;�+?���|�ŧ��?s��٭�|���/�W�����Ͽ�w�>��r�����0�{�œ����4��l�yeO�j�rٷ;B��i�l}�`kB⹰�*�{�>:0���
�A���5pr�b>�bػ�O�3V�s�b�eֵe���i6�J�p�t0�Y�,j��E$��Z$gE�0;9a6;E)ō7x��W�Ӕ��G|���<y�������Rx�L�*	�G����}��b�I��%����p�3(����霣�#v�v0m��{�x��)��dY�i%���������;����|��cZNOOqy�h�Õw�r�={�������9�z�����w�̵_�E�8�-?G��1x�^�(ʵx�t.�³�ʵѦ�,?v슋B�t�/u�AQ��cR��{Z�Q�hd4P�"�],e���!EQ�e\�<�p�d0ܡ��mm��2;�HUA�b!����V�!���>�޽O�m,
��wFJ|6��Ey��G<��y�XgAl��m�v����v!K��$!O_��pQ�}���#�~0 �Mn��
m�����ت��> ym@&S�y���L�&%W�S�%�j�s�p"B�i��El)��a���#B�yI����ߗ*?�L�A�`X�Z.��$!O3���KJJ��"�H��:"I��iEG1�H2Mk�xL(��hT���bΎ��G���4���[�咦vtG5I��K��U�F�T����l�9���8K�a}����M�e�h�r
��H]���P-�;���i��U�ຘ	�:vL�Q�j����Fk��\�b�+6�R��뭌�E��U�|���AY��	�jIS�Y���1��w^}�,O�{}g�%*ф���脺��Ì�����y��Z�޾���0�P[�����0�~���\�J�e���(��B��񅈶��<����}��@W7LG�5���%j4`�j��1�6��6���gg���E(}(��k������1�a?nxY���SU�"%I�t��u`*Ǫ��p	�;;/9=�SgC�P�J�G9R�\ϟӵ-��I��p�lM�3���Kt���o2��O�0�y���ŷxt^���ɏ��ݻRa�>���z�����^�.�*x�l�c�xw�v����|��}$ynf��uG�i�m�R*-���    IDAT{ҔC�茗)Ks򜵐�`i���Ɍ����H%)�d:e�3aմT�p�W���;|��=�� k<E�3o#�!�2l��Tk궥5��'$I�3���Pu�3LG#R)PBR$��#��
.>32nZ[�x�R�4u�F�w������b�`4,�R��9�þ��f;��ѵ��s��oY�S�#���������C���~��+����0���7���� B@��;_�����+�?�!g'G(�(���t���:��R��#3����qo�����!�� �!�yV�5�<!M���6�2>�UU!G�A����t�BD{��[�V�C����q&_�5�݆P�YG����:�4���qHiHM��Q��?�e�y�oM{<�N�w�=R�H��dE�!˶e0	� ��H>8Fd#";�%Krlk )��.E�xo�y��ԙ����a�:U�E*�
�]Cש}�^��>��i�q^I���5�{��4V6�B�ի�=.�/Qd[XN�����
ʬL�Ʊ*���H..-c��=Ťµk����ԆMۂL�����gX2��ȺȪ�3�Ń�y������goo������L�k����͛�]'���	{��|�j��912���)2��M�"�
m�T�^�X{�z��YJ��#���n]SLj�ܹ�Q���C�2,�O�R��lLMUT�g��<�l��'��	�!t�vM���#��$K70T9N�m��S�X�x�'�tYG=�RG~�D�>�?��6)�gs�)���D��h�1�L�-�Ƣ:G.
����� ��&�<�L|�bݬ���QZ�o�H>��jB���[�|��PM�(
2�K��Tw���*
�e��0���e�����K�\�60�p�����u��KG���2�i<�4��E�1%j��Ww�o>�����_&?>���QE�.b�1�{��,��?�u�ny���8?�r���
�ir��nޤ�6!/BJd�R�IMJ�*�	�T�GzK�0�(�(Ц��Z�d
�. � �a�:�&mF�%J��
�����1ٯՂ!K�!�X'���G�"8lV0�T:m��B0;��d{S�NN�IQ2[bO�kyr�>���;��7Xv��ӊ{����>f������⣢;k�������2��:�#,l��x��us���O[V�Պ]=���{&h��C��8��u��6"�5��ľG������L(\\�D@�B;�0�D�DI�t���y��<�0�nN��W)DDjâYSL��c�Z�������w��Ff0t�L����9e�"�`R�T������MO�IA^�T�Qd4ޑ������m('j�yI��pѸIɉ���w=m�Aeh�6�v݌48�2)�!3%FGz�!���[t�]�AM�8|�m�pO�P�kd��h�X.�qP�(YQ_+�5�!��<�|mJ�k�TÂ�w�����C�O�1��c�w��c�$uq$�/	Z�.��uuQ|t����Hb�@x��S%�/��J#� WeM߰s��S�C0���2���=AE��D,q���k�dDt���;c�i�7Ivq�ϲlk��.�����w@
��~��1R���䥃����Lf��*c�^�)M�դN�q:��	�ƚH)Y+�M�N��q�@\8���2�������9�6���i����,]�z��oi�`'���K���ZI|$�o{K��������ՒfhXtK���/����R����WS�n����dǆg�眮׼��_ i���1���œ�,�)�$��G�u��t�"=�m��ﱽÕ��/>R�%ӲB��^3-Kt�aI��,����s�!&�fc{�gǄa�߬	�����4��G��Lx�n������-|���L���0,s^y�6/�	y��w�up�n��ɣ��L���/�
^R�F��˗S˼�8��e�ڢ�&�\f��t���Uhx������3��6-������Yb�@
���"���Р���v$�D�\d�G�v���YF%5�'HI�����c��w�H�
={��S�r-��2G�!��B^��ag��Pƈ�7�����ԯ�����*c-&�v��>���������;�Lp��T��!�/UI�O�٫���;NGcύi�R�d�9��D��YK�Z\�	x& ���*��X$6J���&%@�ٹ~���=V��o��!0��\���99>���)�����$��z�⫚�|���YY3�4Z���h[����r�&SvgS��|���v���0(S�xG0+k��������?�G������<;���-�����/s���,�c��(����H~S�|ÖQ��h����S5�X���V���F!"B�ӳ�m�~�pCOߵH]�Gf@Ha.1���IE�5|�����$�.u�#KM�X�S�O8���#��3��AF��������d'��b�~�c���X�B��u!��.�d�*��k��H��}�b��N�Ʉ2x�Ѷ�,�[Oy^�Y�c�!^x�xL1�����~����������r�����G�O�`������z�͇w��O���h��a(��'J��?�Y����ߤ�qQu#��I7�/��_�S��\3/�̶�TmRW�zI�!U(�Պe�o�#��7*�A��f;W!(�r�#�Akl�$�̒`t�)�F�݆�4]��bZS�u��}{!�����Lx%
��}9��+��c��'j���A�w��6rm��~yJh&�y�(*]�T�s8�EAYO�A���Yl��޻�ү��U���r�!@�<ē�=����ٔ/�k���������t���f��g�g�x��k�n2X�0h�3ݝ��(!�����ί�g�_�9��9�s�S3�kz!F�'zO�3vg3d�Q�i�l�<��_�:e^r2?�]���"��h&���7����Ӟw,?�ڭCz1`]I�_1?}Aa4EY�|q��Nx����b���"��h�q�Ft!A(ʪba-O�>bg�o�r�g�������گr��5vg��&���y�����?��gl?�n6�eAY�؂�d�b�BĐv��!�d�,������kJ�h$� ��|������;ܸu���Xm���C�Q�F�����&!����P��4�+��!%���g���{�'焇ϸ]L0yB���/�T��リ`��q��6g~����y�OcR��YXY�]B�J1��SM�TM��I���� � HI� E�"~gbJ�&ܺq��{&Qќ���K\�S��RC6_�؆
y=e��2�Xi�P� f2�ֵ�L
�r�p�ļ�������,J�.7�M�����wv�59������))ʚ���~���^Ń�	vZ��"Z�ě��Q�#U��Ĕ% H�K�[!cRz%q�(.Q"d�w/	���`LF"D�V�*�LsIa�1��"���@Ӭ��ۭY�N�����r6��$ �Appp���<H��[�[<���{���ut�&��1�Yh
-�F.!���Z�m����80z�S��ڞ;n&kp����5Ӣ�u���O�]/�J��{����ԇ��H�h1C��%�����Ï���z��\rͻ*�;��Ξp����Ϟ����ď9�	�tM{���Y��t�O�9.�$��)���W�W[��O�=B"l�G�9�Z$1hf4:�8>9c�܀Љ����� ����D<IUM�1��l��eB�g9����}鵥�{�<geҟ���,K6#/Fz�2:9x�����}�����=!�\�L�!x�L+ m�#����;���q���o�	/>�!b��(��TEŒ�A"��L+���ȫ��YQ�;Y������)��%;�)�+���&z�Q%�b��<?���R�;��Kv�g\[�v�9^ L�~ߠ�8?z���o�����y�z:���ݺ����(��1�x�b�t4T�����<ϩ��^�iہ����v��{wy�m��9������d�e���������s�<�=�i�5%3^�U����G?����[����S�\�f��oZBHT�0�DS�����{BjL^b��I�J���t}CU��������O�^��vc/H$>�R���[7K�~�1��|�w��y6���8?}D�9��%�^b�J�MtK���-R	|}du���m�Ӷ=�,YmVi1u�i��^�O��(]�{��ɠpk�;3�,C:΢ځ�������o��������������2���㕷������JK^��>�������IiOQn�+#���6�(ï���#�}H�t�Pɘ#+�臄1R���2���
���#�C�h�#���~��1Dr�Æ��?���>�^.�uF�Zqgg��޹Ba��B(b�1|z���̐-�����}3�a:�Ȝ�ŦG���Q���"�Y�s��6���C��9����������C�� ���5:g��_�ᳶ�Nk&2U�%�2�6I޲�n�)EF�y$�b�X��t�h}����_	�N}�	n\�U*'q��R���d�M)�fwZB�ċ�0���ݬ�%Ae��v�v3֋%��f�!�������ã�U���5��|�;����1��J�6�Y���(q�G�1�g\��
�B� �a a��CĈdW�n $&S�e�lR�Uo��	Mp�spp�B����|A�\"CR�w�',A�!S�Ar�����_�:��:d�������.{�N�T|������/s��_��w���)U������48���T�ٿ�x���'���
G�Z�ܥｴ�~�G/�X����a`%����/C�S1"�\0/���zg�~8ݾ�$O���,v=�G��[������8;9���%s�K�R���1�����MI��u ����yJ2t.-��2(Gl�9_���e��E� �8V ����9u]��&�+���B@�nX1lZ��5���ۯӜ�"�ݠ�|��ѶL���g����x�UZ"��B18O^(�� �v<~����g��w�w��	��	�����2�2Ec��-+
"��o���?f��KӵU���޿������!F�(v��)�Cg7@�7tbY�$�e��'���r��to�|R���Y�����5O��ǜ�W�ˆ�j}DK�:����"��9c��]�(��a��VoUېN>Rʔ'>���J��B�d)l� [�i�%��f;|��_`����Ɋ	��$��*�*�+��b���vx��@
�'��>�����Y.N(&Ez�L�����J߶;{����g��7�y���a�\���p�^S��?�2�����Y��.� �eFU�ɲ����'_�ѷHF������_�#^����)�nI�7L���H19�蕯rx�:s���s��?�s�^r1$�ڸ)Vr����I�� Qe�цH5a����;�P���Ǉ�B&��PVȼ�q�� ��dJ�bD{h��wh/�rMT���j����6kr�F�M�.Z������%�~ ���dy�e�@I���8���y񂈤�sJ#	~ G�>F��9�����4/8;=c���q�G}B�zJ�|��_�߿�9a�,Mߠ�H=�q"�ΦЍx+F��*JdRI_����ޏ��N�/Lb!��H��Ȗ�w1���C+�S%؝$k��'M�3O	�<�j�ݚ��Y=��y�c0%��8�vD�3e�{HQ&��jq��y�q���>rvv�u~��1-�C���X�_w�#�d�Sc_UȔ�1V�"-x�X���6!��	��d�~��cĐb�sm�u��Đp�1#��J��C����c^��_b��|��;v��3:JѪ��W�絷>��Y�������BŐ���g���zI=�㶴�f�+���O�Ŷ����{ReH]�޷	���	Wl�ɕ0l[G���>G�n"����|�y��&��8_�B��/��&�|�-b�|��s��9���@�'�|5��w����k�m�r���r�����"Q�V+�L�4���n��
- A�dD�H�`�\>0��b����pyA����9�����b����IB��Fbc���s�O�r�?�^Bۑ��#yl|˴�0�TY��0�+r��í6��s>?�����|G6�$����`WKT�RgY�]��zT�>)"�=�0��;iY�=GJ�ُ������yA9�Q�S��������$+rLU`����x���H�AW�*�m�}�3�z��r��4��{z�������lzס��[+�|N��赛�z�z0C�i�����d��:ym)R �8����DF@��'d��w��{��i�Ⱌ"�B��d2b��������=�uv�ݴ��'�~�b�6+l��TEH����8�������a3�����[��󓧘B��y=a����5*o�ۆ��ǜ.>g���<e��9�9��f���S���q�Un�N��	O���g���
6��:���{wy���k���߽Ϗ����	Z%?���M���v����xk����jֶi*�BC�yE���W�0�>�
d�)	��;O��>��%?~�!��1��.'�AѮ��eF`c ���FIC���;K��8M%���e�v��=�v�z[v�!�2֍m��n9�m7XAj�d����w�.��� !6xĦaz�h]�4>P��K�a�S�ܱ��yDs�L'X$�$�Ks��j�>�vf�W*.�_�21:��0�h)e�R��BUS�uPt�"�H1ý����=��P�SZ'�J���}�bR3��FU����(��,���_��_�9w�ܡ?�������~�&�sb�m]%��0�.ӆ@ �  ����C��f��x
,Y�]r���0ptx���h�pI 0Z�KM^z6��(�{�U>��o2�ȣ�}��������fj`>�������k����x�k�?|L��Q���BIu���ӯ���i�)����9� .�$��������4����z��@���ߎ��G��h\,�&=�V�-M4Ƹ���� �����[7X,<~x�G��`��(
�z��(���Jz��On�i]��?�U��x��>�͂�C���v1_quч ���{kS�Q�ԇ�EK��V=��1�9b�d2��Mƺo�H��*/�OszL�)���YRhA9)C�Q�b��?����{�<c�^"�����д���Ү�xg�Z��g����2�&(�&���N`�� q���>8ʲd6ݡ�Z:�R���G�(�Δ�u�|�Lj<ѝ�E���Δ�`�[�����i�������+2)D���ap�#W�A�
%�7�F�]���U���4��/�I���𨻋r:�C=ۀ�@�c�IY�,-.�%�`�A����4L���}��%�9�!6���F*��)$e��	���OO؜s�\0�n��ۆiY�E��$V�a;1���C����x��o���z��)m�0����]v����g{j��@W�e���MA�˔ 5��f����|��|��}��P��ǜ}�G|���5o��z� ����1O��m^y��W��}�7�k�x��$!"b@Ȉb��M���,�. 1=F1$R��0�!����1�:���h��]��(1¤��T��@�R�F��#��eC,!�YZc��rS�S�sl��p��܀k�8S�<74]:���dfP&�]-S�A���\f�iA�uئM��i�Ԛ��QH'�r�1�͆���
^�,5�&�4f -��1%���~�ڂBd��eL�2��P�C�����2�}��� A������H����>�Mj�4�3���'�j�9�YF�肣���v�6�iͺmȲij=�l6���#����x���y��1���{���ہ�����<l��i2���6�)�S#3
!c���d��Δ<���	�ł�|���	{{{�Y��SǺ�Y7��%�i��p֝r�k��AnPeΤ2����������4LKA�:���9�7��'��)s���>~.KK�߸��,
���\^����-G�5޸�]܏�ﺲL)AQ�����B�qc��ڂ�6��g�5��^b��+=v!�n���͛87��~���I�)�j��&������OS!X�V<}x���d�7�|b<^�~BL�<uы�����R�2F���6���3    IDAT�#���Cg�F� ��CM3\�Xl��(��5�Rc̟<�9���y��=6�������X����f��0��Ɇ�E=���Ɍ�����BLo1�e��F�(��hi(��]�X��s�IL�~�IB�r��;>���VƄ��*��I�+gZQLk^��3�a��sN1>rk��:/�C �K�<��]�퀨���B:�`[BY����Ct6H(&��f�yp�!�!���+�u�p)P$���������@�c��m��gd�_�񽻼��c����Q_?"�Mq�a��X>z�G�->�ַ��9ZD���kT���A�*%�� c"L
���Qz�S��'6��̐*�7��2?>ey�1�� �nY��lo�<�u��Kt����L1E���ܾNQK�ر��{g�i�>g�|�kŌ��U�����}L3�p�×9q�W�T~�T��1��Z�e�GP9���\8�{����nI�5cFI���B��
0�g�2'�K����ʓ�ӶM�$�r�&���#>F�LH�`��`��(\J�
)�Ʊ��s8g��"7��~[�̔�.׃��:�U~���&��}rAL&6�%�A�(�w�L#Є~`�l����r��b�@�!&d����=1K 1&s\�������V��N���~m| �H!�*R0���,Ӭ��n���(�(�}ץx�iμ똾2cg��w������_�9M���2�v�����M��w��,V�m�R�2�)�,�q#[��VWpebB�BGQ�e�}�6�@UN��rrrB��5�xⷴ��n`�4Bk����'h�A�t�=���S�32�9YoX(�ΐ�%*��Pm��y�`~~�6#���jtk���'�[�����r�'��'���B D�O�2�>pl�0۹���EW6�Gy�@�ud�F��!=��g��\�8�gY��q/Z�α��������z�6J�����`�u<}������}b��x��M�Ҵ=�t���>��v)%��pA��ap�o��R�6@/;��O��d�ߎC�F�&4�$�U���C���\lo�e��8��4/���~�s�G}$/+��#ߛ���U��Xω��7k�~`�]"����6H'�^b���4�ki�h��=>J<2�������Za�	ߵ���|0�pAx��N4kix,U*�
ϑ�aS���y���#B#�k�f2�8t!�B ��@ָl�xn-1Eq�Ǐ�q�QU(�ru����6��@�%ꝓ�b��UF1�C��{�kYFK?U{�}:�̠���'�������c�h]f4��z��l��t����@��k:��Z08�Dlm0���)l�%�L4�(p�a�r۱~t��8���%+d0t����8���yF^�Bc��w��c2�����k���-Η'�K���!�����\U���[��	��y&#���u����4�9������@@(A�;FE�On-eb�K���c�9(�Cn 7q����a��)��Uo��f�jT֑�7���.2�H���SBH,ta@���S�9JA6n�Z�R�.��LJ�"O��n��20&c��ɕU�G��#$����:|!p�"�@��JR��B���>_q�h|"��QZ3��5�w�9��<MfpDv���%�~Mɔ�;L���Ð��(�`dD+��)PIF���d���8nk�+F+\������4��6]lh��t�k�>�ϧ�o�^��7!/����ES��凞�v'�]��೻H�y�wY���Y�.05)<;��vD���u^$ؗ<�+PYI����CP�6px���}����y^�ٖh�dQ�2Td��I����!��JCA�\�֣ª'���	յw9�6,�d�3��v��֫Մ��:m�����d&CF6�ֆ+�?�
�R�~)���S1(|�XzO�� �$���V���e�2�����`AI����1t=.�ZbmG��1L&q*R���>S�0йm4.X2	RE���a����$�sαi��6�2o�Q`�K��Yr�)��v��ιq��Ɍ�dB?LgYQ�Y��l�j~�b~N����!�j��B���H�L���r״4C�D�uF�NE��i\&01q�e�# �7�Q%�C��s�@�sG�?%�}��������s~r�t���Mn�.1������]�:Yд�x���J����F�r�֢tgΟS�Ȕ"�`�5�`���o���RH��c��wc���{Lo�s!5�t�jgFV��� ۖ���
��+|{��K����8��%��ͳ�3���r��>Eb�a�)$A�4n	���%�2�K��Q޺Mp����Q�LQ"�m6���{�|艡��[�w��P_?�>����1��:<����C�]m8�ڀ�փ�0��BM��Ve���E�HB]`�@4�Tl\K]�{�X,�s�Қ�[�מ�/�^�'3VN���<�Q�+&N�G����d�1e�λ�V����u���-��2ٙr~���{��j�����\�k-%��T q�y%>~"Z$�e�2�,�A&UL��(5�[$�AF�V�ٽ��
���5&�(.���s�<������9�yՊ ��Z,�N^�Zڈ�yN���\�����>�T�W��?�7�'�2JfBQ1��.&/֖�v�F�d�s�`�Z�>��ӱ�8�I��R�kݹ��aB��Cj(�JH���E�ϳT�������2���|u�G�OYv;���b�Xr���b��Ԥ�,�"~����}�s,s>���9~�9Z�dF�t�^�Nc�zCn��EfG�va�{��������l��s��&�7��n<�z #ŗ-��c�ko�F���Z��'�ke�,��Q��������?��_�&����7�y��<?Eَ�{*Uq��� �g���3l�%�MHσ�����?��ie��cn���0w~�RJ����۹չ�>�/^��w~A��1��r��D����R%/���8���)B�2�t:�Mi# C
�j���H��z��V���4]�67Ҋ,�*�m��w�\B$H�*ac+!:K��S2��)sd[�T���K�c�wb�H@���0$O��W�x#1;·Hy�Unߺō N�L�g��?�Y����}3��,S�}p��o;��5�b��c��ꌙTt�\7�uK���l��+�߼��)������͔"�@��>cdR�R�V��d�w�tg]��>?�'��,(���-T��������D���l���rC!�Nf9�h�>q���m��������j
ȯ���7��������Đr£�2��Y���e$��V����)�[��R��֊>X��7+�}�!/���"| ��Q����x��� �L�F�|��k�L-�(��C�H�w̐|���<}���^c9?gRܼy��zɭ�7�d���ٯ��\��W���������y>���a��6���an����v"Ju�lw��������w�ѿ��'�(w��BI��x�R�3��}ZąN�-.^���#S)�B-������w�L>�����ľG������TR 5R��!Dr�GL3�ͼކ9��U�^�%�K}ő-��\mk�dϺu�t��_�d������qǲsν�3���F����mQRSg5vpa����2ٍ��؛��%��r��^��F��O�X�������!D�����s����NM�I�!�"S�ϟ��{����9�����'4��ǧ���Ą�
e&�h˚pp�p>�9=���\z����b��v�!�+��-�ږ�K��l��e�3�<�	5i$�L�w����@����-U��s_~��y�X�4-J%T�r-�v�Bv3���������x헿N�7��sjc������9���=����I�ٔ�/]?��ű�Ӿv� ]� ȗ��/�̾8/7�i�_�]_�T\����yڴMײ�;O��֊�s���򒮳)Q5��d{`���M�Mn-s� R�hR֊sE�t:��:��iZt^Hڡ�X\%4�z��j}�Փ����5F�)j|.��㽸̙��ߗ���*�������E����u��L
B��|���!QDB���qH�M? �B!�Ҡ�&xI�gk)2��5�`i↮W����`q�K)��N���:Kc����J�H���!��*U����(�
�d�&�UUSO�(�	*S�l?�ڭ�O�A�:E%v� ���K����d��})+��$����(�u�%�unX=y�p���'l�|^������$2|0�q�$�x�,,ro�+�]��Yl�!�JV�9Y.Pr (��O����k-m������?�M���d���%u]3�ԳG�$�)rڶ��(6��:|�_��or����_�~�!�o����.��9�bF^LYt��|�'�g��	����O������i��ʗ�A����dX��f|�������؇�q4�2�����M��?[)�N���')��5F��v�̍J"rC��	�[oQ^���k�4FR*A��"zv~����,Yԉ�68\tTe1Z�Ҹ���b{Z������m�,��%��&�ר$�k����z�:f_�B��M����c�0��BH
�/
����y�_6�[v���o�q���q.J6���'�u�������	�*Z*�wcO����Ag�:r�s�(v�	�4dY���&���p=|������E��g�x��1S7��@-t~��p�#��Ͽ�_�%��kt�d mǦo�MK���0�FѴ-&�b޼�ɳQ�h�����04Ӕ�=M�p���f�lFx|���Ӈ(I��ABg�G��LX�M�~���?k���?r��ց���"��d4�c��~��w~������ѓ%�rL\�����'��_�U��j���gT�s�QU�ґq�c�a�/�ɤ�%�M�ӗN�UU�`�<!������Id:�R��ݶ��\eY����\���#R+���inݸ�믾F�4,�K<۶�(��-�z���9���J�6�52E$�b���\`�H��xA�]ZA\0�K"}Ak�Hz�ȴ@IM�K��r��ЊvqF~������9��۔u���؛�H��g~��|{Dd�VY�U���R����DR���� ��m�ط�����a`�پ��a,�D-�Dm��ޫ�k_�r������դ }@�2�2#3#�w��>�ؾ���������f*ӷ���Y\��'ۺƶ�m�����	y����	��3����$�)MUMs���cuG�.Dq��a#��2�PqB�dE�hg�>t���r�pL��,"J�ާ��T���3�s3������E��:(X��,U�dH�IL��/��W׊�5I�[��%���?su|�ۿ��s�i�ȭ���4�z�EŢj�s�R����9��{�qrp�m-Y�й�4SD����m���wd:�5������?�K3.�E!PBFj͔-������Ǉ��3�+_"�Z6�"mz������=����N�G�e�|��`s�2ɻ����'du� �?���������"�F�Ve�bo��<y��?y��*�lЙ�]��w�:�.djGJ����bm02�xܲBw��/����B� JE��ȥf3�qY������OnS{����V8)轡�-i���5!������M_�rXе��$�^8'��l�p i���	f]A�����������^�e�g�9�u g|�_����W���FGpt�C�~�'���f�P�g���e�IU�9�/���G�0w���P�n���j)���0^ctD�:��8�!U.�6=��8���������Gwyx�4�IT5��[������ЩY��J�<~F]�am�P��uI)���ҀN2�����TΒ�6�k�<]������R�Qh|JIPxK@���i898���a���ZGHI��,�A�<�����r���?��Q\��@$gG�f
�i��Nf��);�-n�����\h��u�a�bm]\waf�U������������U!�!4+���$/\]FgY���q�[�$��kt�q������<mFq��������Is�� &��.fz�֭�oǣ���QJ���SI��C�cw�ܡ�*���;�ƽ
���{�+S!�@إ|��
���xͳ�����!�`.ZR<Q��p�R���I҈��'�D�}~��oB�e�4%�.�k��P_��=ASk]O���1��إ�����\`M�="��uG!5�$���4�:�j�X�#"�W����RR�'GE��2�8J��`H��b0&JB4�P���1�����Ɏ��ef��I��t�%;[\x�gn��Ӌ��B,���bI)���$}W3�9�����c���V)f�&��(�IV8�r��F� 9�JH:�S�-��f�(9:xN9]�����9��"UT�)�p��S��5<��{<�s��K�|H��������&��ᵝ����-ʶ��h�O~0�����l��Ï�t���;��y>?�:;���������jF}p�~0 ��=�5<�%9��h+�֚�FFU�x�M�2t ��^I���D��j�=oBjb0��n���5����C�/�-��0"���I:�c5F��<eQ7(-ѱ��z���!�"���dY���MU3����l)�{�������D`j�i���۱��.���,�/�X\��C���re�)V��b���֢�!����Cڮ�Z���w��?]�'	2N�:��8Y�$ŀ������b�l���Br��=��Ha��Bi�TEc{z�q�b1�D��j<=|����K���|�uT�QWU��ZKo��^��(B �b2��`N��Kv�!�	}F��q�HSM��e�9���gDZ��K���CQ��Ӵ4�'+r[� %�ix�ZD�b��l8b�d�����7�dQ�"�3"�Q�Ϩ���х^Oˀ����I9g{0����O�&ǴiƖ���n�AJr>ST"Xa�%A�������&�}��������?���>��r�B���w\��cZ�?.���SEx�XT����7ߠ�~���B�D���麞�d£G��z�
{�;D:aP���Ή�E�P�w/2s�r��]���)5JH���YY!�g<�TD���s�J1��Bb/M��LP��$���J��E��K1�E��ۖ�jЛ����7ٺq�����>c1��E$��{�&��:"Orfu8ꮽ�g���,�ԧ��o�������TmMUUP�,f��!��$��ic�h����#���jM۵!)HzV�R(���t�4!]�G��8�Rc1Xa�	H��;�tZҹ�.H�׎͗�z��B�r�^l���5f����c�|�;t�a@7Ӝ���)Fjy ilX���Itt�1��8
~u��v���YT3�yAd����Cu�V��6�/�:�Ђ8Rt}Eߴ�Ռ��FG�,��.8Zkܒ��Iw��߿�����s�i��,�������]f�=������1y������mIi6��r��qJ#�Ɍ�ȸ�r���8�ġH���!A-����A'��IQ��X"�QB�}X��y�r&���/�:��j�F��qV�$C�ӜQ^໎�y��������s�R顣(t����A�h4��w���ի<z�w�2�L�s����dc����a��뗃�.�͋���y��"����/\J��Љ�|8�P����{<9:����8�˯��JՒƛ����pV�`o<b���{!II�e̒'�9�,K�℈�Ak���8�'�%�wt�	�W�s���Ř�HK\�S��E�Ԋ�`#�b�C�)��3�3�<	��3T�s��sԶ�k�gg�<����+��(I���._���3�v���`<j� -�!D
��-+��3"W��g9q�Ӷ-'��̧ST�)�o$��9�Ɍ��^��5�29~�u}ٱ��S�̦h��(�!
<���"���	Yˎp5�Y��fG�"�]��/���
*��C��!K_�����V^$�����W��n~P���R��
�)g@8`    IDAT��!�g���m���23~������ӎh9
H����W���b��֊s�����<���cL�A6���i�<����h��dB����^,��VϽ��Kr�U�BJV�����Ձ�A���G�-�,缮i+���?��;dv�S?�7~��]���O��������^g�4$I�0G��s�*K�tD�br~���>�I���U
g�=i7?���+�����m���C�Ƣ������wo��w	g%Y�#��F8v�I��X�ϵ�D �@y�QB��р(�ıy�q��bd$�M�-�LI⍐fT����O��O)|ƪk��&�Vϊ&B�����{ּ4��a`r}LOĹ�q�������@�G�FG<��T`�fqf��cL�!�$��m�#�3���1�(�,fT�)բ��e�%R�'y�"���cA�O#�1y� ]�%�z�"��ֆ�Ju���W^�8;;c8�dw��A�9F"���%�����+������p�����,]S��5�Pf2C��/�Nx���������-=�����uS3�EJb�m��ՁLh���Tdd���1ny�Ǵ���,��P�nSu�4%�Qňv�`� ������X(v7��(
��¬�7dJ�/=��,[V��k׮���G?��K��Aü��l@~��KҞ�iB���v-+zis^���~��/wT/sL�x]\�>�&T��Y��_��M�����pew�G����'��!Y�C,��윃ɔ�(�q�*ۉ��s���$��Fx�]GgA����Zp=�� Kc�y�1i1���i��/�S�UG��1��>��}���.�i��&Kr"�d�@d
��C[��q�#�C�LאHM�Z�v��p��í���È�y(�c��x}��I�8Q�W
!B����-lo����i5���'�늫W�p��WZס��wX�5�Rxkq��)��hu��5��[t�5�Â�VhȲ.���$�.�g�L(҄B�X��c#!~Ev�箏��������Ϯ�/~Ϫ��鋦��[��\ �	�����v��c�!�\�;i��̦ܿ{��ȉ���i����)�-�G'$I������$���Uų�O8=>!Z���qLoJED*�/Fˤ��l�`0 �(�*WM�p?��Y~�ug�P����_`ݯ�{�[��@{lS��5qs��`�%��tP0`A��w������$W6�5:����Xe�M�(���x��4������"e���"�L�8�MϐQJ+s�s9͹��Q����C�L��&�	��:�a*Vi�R@6��$Kb��Ʀ7�(��A�(+P(�,#m TLEha�C������F��o������h���p�ӵШe��c��'׭6�ē�HC.m�ಁ��$�1�`m���������_�"2D��|Ge�ӊ<+XT%Ÿ`Q��Zp>9FyP��l��x�p��t�SNϘM�0�g�L�'g�E���s����ɂ��Ì���y���^�w`'5j�����G��"[��{y�ݯ2m2����f�T<{��˗�y��kLΦ���3��DOK�>B��Ӗ�?�O�݄��~̞P��;��d��;�~�������#������J�~�P�г&Ġv��A�LN��U���&2�@�hk
<i*8�:j#����餅��8�!�CHŢkH�?�>9�ѤDF)���53$~0di^{�u�����T�4�(��*�(��:��9�ٌk׮�X,88|��
-�Rfx�[���m�ش��{A�#��)��Y�Hc��3=EQ�4MH��EA]פIN�5(��25� 0���إd�X���|�y�����fƲ�[BߑҜ>{���1�x�?��;���=�~��rN����9"�y��e��qzD�D�M�gX�Q��Ӳ'�2G�iq�g��S�1s��KC}2��=٠�v5�������G�v��kWI�!'���|Uc5A��A4*ȣ����j1�;���4���㽧�mբ�.�}��m�|rJu|N���Q�c����O���tޒ'���`csLg����渦�3���G<��Sn~�U����x��_�AD1Z��`�B]:!S�t��G1��pI��N4��Et�(Np��Mc��O�DEA�v蚆>����_��CH�Z���1�&��Z�}��n�%r1�9���`�GE	�W����QBg+��(�C⥫QV��m�A[�0�}D�z��`Lp�Cy��AJPĔ�!pض!��~rvww�2x�;<G�D4]�B!�BA�ft]�J���ْ/#��ix߇��8�֙J�~>����`kg�ݽ=�OO)����i�'���*�0֓�;"�KU�s�#�[�8G�Fsu�/����nB�Y�R�X�o{�KrWm��a[�>{����_�F5�Эe�5},)���j������Ӈ��ߥQ 6�8��YQ�x�2����S���3-��0;|�sg�v6i�������z�5��Ǜ�(��:b��0�ZDA�8H#F:"�"!8t	��E
�����&^
ـ,I1⌤w�k�I�^Af1�i�\`4�	�����g$��C�A\U�A��r�}��_�އ8YeY���-=j�Q`�)�5t�p�e�4&
�D�g�:��􎪪hzK�&������qO���U[����&��6(?y���4m�m!1WǗ��y����=��bF���]{��K�Yɐ�K����[4�A��+d�\g��I4�@]�IҜ���bv	����go�{��g�2i{���m����0�r�EE<���o"�7�տ���_�)��=���}�{ޠ���o}k(�Y�����Zǰȑ�cR�)tF��kz�	Lw��ޡ���$g�ګ�"c0*���������	����ɽ��<I�����b�u]ǣG�ְ���y 8"ְ��`5�_,!�e����W��r}ȯf�EQ��z�]��4M��

�p8�,�˟-0�ǹ`��PUޫ@Ҳ���+�~6����wvȠ��\�s�Jp�.��
_��*�o�?��Y�H�(�(1��xƢm�*&I�S���|��K���!�Y��UOU�0�D�!��T���Nx��}T����]E��DH26�G'*ڠ\,� Gu��JQU��/�&��vđd#�puE?,���)ܴ����C0J�;6�!��qI���4	{j� ���%r�T%<��!��~��-��6���d2��� �b����7,>�˕������a�%BA�	��ȦGws��4��dE�Z2���B�l} ��pK��������_J�݅P6�0�'�
���Y?���`�������c�c�AX�}�$���Cv��خ�����J��c�$C�u0;�
�(<�4+t�P��f孻���nܹ@�K�du��foo��bA9_���{��M&,�����	�ąl�����9O�wƗ/�R���z¡/B��2���f�>�s���?�{cҔyճ�w�^'<�gă�"J�yN���ޑw���x��{���R�l�x���������u�<��	?�������U��t��tv���%����Y����QR�୯�"��q�����矑N�l+ʹ7Hy�r6Һ�ES�ƚH*6�)�	���;���1q�Ru8OJD��^���T�e@� D.�?��g��*d�@�&xc�
��tN`��i�����x����!�K	�AY����{ϏPQ����U]S�5Zk666pU�oڪ
3ʺ&I2\�s��]N���`@�Y�?�����(�q�Ķ-�|�`���لj^�s�2�c��G�yp�t4୯����.��v^��5�E�x���$gZ����N���<J����>׾�_P-J
#�]��&�g���\��WQ������������>v��
*�0Xu��6���XcKI�RbZ��;����t�J0"��q��w �l���<b��>ͼ$�
��ڷqՔ�yͣ�Sd��P!��kZ:�/;����cf� ���>�Zn����`:�2��և��,˖d����{�<�C�X,.hw�uW�eYx�����j��u�I��^ҵ�:0e���配y�!�b]DHB��`k�o��o��7 �A�b�'��c����`�bs��miNQ��AZ ��E�r���"���{$=�,"Q)���	B#}B����e��ۢ���z��/q��/C1��Rbi�Y'�	>R�2>��tm��=m[3��� ��eE��8���
�o�gz):X����
��t'���12M�3����>m]���9V9��<�)�0�*�il!u�iE7k��%��)CZOId�QI��з�`.�
�F	:�1��$�	`�k_@����ř���K������r�z���� ��y�j�V8'�횕��A��9�"m�29ӡ�aT�L�����[ ��$���{���Y(��EmX�t�ǩ�I��a�w�E�h�7�7K٪8_�+��{�N�{����4����ρ@�K�)4��PK��i�
���vĊ`��`��ř��0Z(�P6@�\���w�7tI��u�2�+;���\���&U9�_��W���_A:A[�|z�3�ݧ�W\��d^�o�3�!���X���[||�.����}���#b�(�����2�R��!V	��=���L��Ԧ�"a��k�_{���6�u'��B:~�V��6LS:� gP�bzFy�iʎ�u�8�lk��ش�����2�_�刋�*/kHY�}���ª�UG��7xQQ�!=��s~��D��)*>���1j8���>ۛ��}�+��c�����q~x�Y�q��	�O?���sd�#���nQ�^]7��.�s�D7T�)�>���
���<��k&���|�A0���ާqgyz��(K9��=66�RE�hGhz��cE���������׮���_ď���j�"�˘N̑��v��M�ʑgr�u-�qt>b,b&ˍ�8:��^;�'����{�9q���ۣ\�Ֆ���L���t]�O�{�J}���ì����\�0�9x���#�.xr|B���j�ozi�����8^�蛦akk�W^y��^y5��ʒ{������������(��׾FE�eIYιu��ł�ׯ�ꫯE	>��������_�����LǼ��;\�|���S�<y����ឧ���k(q���e�(_PN�ˤ�U'p��>���L�g�I�ޥ=�gO9��6f��̬G��D{Hbf�s�5ԵD��D�� %���-ie�PF�4�aV���R���'h� u�\x.�W����#z�	F^+Rb״a^�Ĩ(�7�ଈ�k*��B)��=m�PNgt]�d6�3��,�?y������B`���w6���7�w��'��x-I�<͠3t��d9��>���ͯ�ŵ�{���Q��
M���ofO�a���6&��G���?���6�<gR7TQ�V
�͉∲�8�%�J)d���o���qň���;�/fϯ�����!֭�J!��D� ����/�X�ڱru)�R���� '�*�nc�RYk�[��	��JGԆ��QJ���8����:����VgHBs)U��Yv���0�@�]�?V����ڶ����R��s"-��!~�R�����2�2b5�>ح��a�Dg�/^�U �*=j}#/I�^���_z�����?<��	�р�\����Ư�
U�o��f�SNΘb����+=�͹��;�C��̪#,�Υ=�-%�ł�tZ0�#u�Q\x{
��і��	?��Cڪ%W_!��f{X`�	�-ޓ�r�.�p��>�<�s����+ڇ�I�Q2"�k��x� ۉ�-E�!�\/��-	O�
�/dNn�)g	M-;��+TRd1�����o�{�7��]�Wo��ƈ���������ѝ;TbH�3ؠ�O�OO0�=�W�T8k�G���}���`�gx%�z��YΑ3��ڑ\�c�������Zs��]<��ٌ��Cv�v�ڲX��N�t>��l5ἱ���_B߸�1[����~�#n|��l��T'�]O$<Z+�����?�	�G�����L�= Q"T�^^�J$R��p��-��f$S���7�mQJ�=J�*�ғ����.��Y�l{���=��a<�1)Q��d���x��ã�܍�xz�q��]��+�����pȍ7�N�y��)��7n\�޽;(%��uM����\�z��w�2�M�y�&����u�w~��!hۖo}�tM��˗y�Ɨ�u�V��o*�j�[o�ŗ��6M�0\g�2�g? MS���o�����W�\ᣏ>���0H��Z���n�ݛ>������\���D���>���)�iD�E(E'���8�'!A)��5dw� ��6acS1�K�ְ�MkPR���ǒ;&������.�����Dv�yD9_�� Or�,�>G[ͱq�� T�w��[���Ԏ�x��8�c\��=Y6�ҕWp���g�ќE�C���*�^y�eTƠ��*l�2ր	I���ls��e�._#�7���#f�D#��:��4�aB�s�5��}Zbz����3t��l�\�s�W���f��ϵ�}��xm��E-�����j	[�BE!�j�/�2���
�_�?C�_�f��	�� �5Z$ĊH�T�x�v�b�8ia�߄,
�%B*LGŀ����]F�C���^�PYQ�> �K
g{��K>�'�
#�������@�̝����AdKc���B��^��\k)˒tsL����y�B��/!|)�R"](:�R�%|x�׀�� ���_�.��X>��;����x4�J\��:�GC�����/)�D�7!$&%����SlP����d³�3���PZ��c-7�^�*99>�VJ,���Q�Z+t��kI����4O��w����d*����(fsc��
�t���ټ����6����l��~���)M�gZ�2&�z���@_JP��xo���K���8���p_k�C9�S��AKɈS��`�(�t}G״4MC���8��-#d6b�����M�׿DO�R�!�^(ꦦ�{��M6߸���M�'�9t�	·$QB=��u-�C��(���ΣED�3"���X�S�K7��o���}�g���%������%{;�H*�T��c�'�Ov4��k2� �Έ݌������ ��|��ڗ趷��	���O�r�o����-=��)�=ZxD�p�R��-�Y�$�m۱���[D���f+�����Lx.E"@�|�[�?{@�#�yI����I$ׇ�s���g��Mn�ʄU��Z#q�Ya�������3�F��_}���� I����ߧ,Kn޼���v���o��ohۖ�}�{�q�����������Z���ש뚿�˿�������lmmS�8��?�	]����~�$ɰև�~�PXmf~I<��`���������R��O����3�'O�7���
�D;h��6���"�Q:V�Y��0#��nBN8:FE)�aQwX�t<�
���T��}���"�qDt��O�iN#�y	�Q�����R@g0�29��u=��o-I�)�E�:o+lﰋ������@6%��Cb!P"�"خg���y	*e��ʠ��%!��1��'癏�$�$M�bL~<Ab�`k��x��l����G�$�&n��OS�������nL2'o����~�*����#�����7���&�����n2���8��?��O����������!B�����Y6���/Pϋ��*�8�o	YDw��E2��[�W���RQ��5.�5�#�|�R.4US�M��1B(�5�}�$��fQִ��	g�A/�(��|��P�%�jm�s�#�U+4a�����L��(XK��4Ib�%I�p.D,��^�����/sb9�]�bi�*�������C�CH�"d[{�r�l%
ml���%G�O8:;g�����aQW�e��
�(�t;,�����c�����svvƢ�3�q8��g8�0F`��B���=����B���I�$A��$M3�����hw���xw�l�з��������������'��1�Y� �Rt�@VxT<��nkA�*Q�2Q�Y����Þ��:>8o	@� �#�%Q�yU3�d���Tc�.�s�שN��D���z�t:a�ꕀ�8W�0y    IDAT�R��xr-Ȋa5��h8<j���ls�f���çtUKLJ���H�b�VE�v��ބ|j/�2b����2����_�
��������e��"�2E�dzF[-8p��waN�,*QX-2b#�� ղx~����8��#�������U:��h��ʲ����E�@���H2�MJ(P A�P@� %�tV��2D�#b�y�%1i#M�7A�7��Y���'·�LK�ۻ�l�yv|�ｇ_L8>>f�&�ˬ��o����3H���_]+B݊�����v��y����cm�y��Mz�қ����u'�X,�N�|��G='�I���|���8??�֭[ܹs'��f�yNUU$��O?��Ç��_[{{��$��f�D�_���+S�����R�"���1�3KV&TJ�'���k�:�^ ��h����q��LK5�`MO�){CWꦧv%����H�(�b��&J�$[CT�����_����{�:��=�a��(4�жd:[ར��P�qDWUH�v�4`� a�� �@�0;=a����	]���!Ӄ�Tu�$/PJa���!d%�}�!PF#I����)q$q]K�S.m��#�N��ܽ�w~��g�[_G���-�$e^b�#d6F��� �=_��o1ڸ���U��(�1٫o�|{�v���_�'�&^q2.�����b5B���?��z	����.�^Y��/��O�<l-8��m��V
�u���T5y���wx�d�G)REk�t�5Q�eKS�(F�(�<��<\�>�����й{kם�Jκz[k�
�	!�J���EJ�'�X� �'Q����9:
ܪ�HB��_�3��i�!�@�݉���ǯ֚$������3\�}���Y�Fk�f���]f�s>��}���խ/A�s��~��OPڳ��t]�p0�H�,�@'1��خC-_�^��%�"�#Z�SwmH��Ӣ�"J3�Ԉʺ��=g���gT���k�JyRO�R���!�g{P�k�\���e����u�a:�����X�o%��d�JN�Y/��闻��'^�=��BI�� ��GxG3!8ím��gS�@�G��/Qv-eS�%�XÄ1��hb�ED��`N��@����U�L>��&(B_R���%q�A8�f���8M��dL-$.���ӳ)���g,f5��)��Rv.mr���<����h�=ۛW��g��k�뢘ڍ��m��6�A�n6`q�c>��"����W~��='
g��y =�	����ˊ[��k�D��J��*�Z��ٌ���\�as{����'HT�b�t�F�w2gZ='�rIV�g���ܸɍk������@�t�|Q�N�zK�Y�ڬ�2V�b�u|�W�]�QU��(������sNOO�y�&��۷�u�7n� $[[[�u��L�%�m����QJ����`0����<~�!o��6�����u]���ŧ�~���_��9;;����8N_������:�1	:�����_�W���?q)S�mO��ˆ�8�M9)��kZ�8Afe��qu{�,����w=�I�Lq(��g2��#f��aMPY��B���kQF�:�3	B�����>��ݿ���}���y���/�9��c�y#OE�Ej|Gm��a�<���]��Z��Qu5������D�a�Z6�`#����nLQ�2���&]C�5�����=��(�>���C�}vH'2�ؓ8O�c�k�t��M�FC6ӌ&$��
�0�r��IC$3揎��/�#��-�d��]���1�t���kT����5��!���e�~UH^6sy�KR����Uz�[bE([*�.����D "!>�g�$J�:ޕ,4�2����ײ�<���a�g�Sխ�E�HI��(Q�ܶ�löwí�F'@>���� p���	�;��r���IY�"YE�����L��i���=U�$;��B��{��}�Z�����lӴH2U��h�΄ �X��a����:3)!���L����!Qk��{Oc���)�4���M���e/�"l���=�`����e<.�Ic�c^,x��_ H/:��GX֗�ۊ��hW��02�[=�A?c���:�bY1�cʡÍ<n�K2ܦx������b�i+�U����d�"��&=��$!��T�"�@Ɉ^2"�N�C��T�"��H/�D�zZ���n�iCP�����~�ǌ�mN�#����b��ސ�(��Ǌ�+�EA"bF�	M&R<
���-RH[	H%�HJ���,!oXCٴT�4� c=�Y�����;�-!@�*#HU��mc��貦&�N#d�1�4*M1�s��g<<<�~�7qq̰��m�^k��=&�	˦aq*�Js�bʝ�(��f^������|�m%�R��2�+��9+k��7�1/�3]-y��O`^3��Ͽ�"y�tV�\���"d��-���mvtN�&�l�87�5Kz^����{z�&������ĭJF[��w�|;Gf#���>�B ��ۮ��Rb:�+�q,i�2�p�܈�Za���i[�sH%ɢ��ȓ�&.=ES�
As���9�~�5�f��p��R���C�s��G��GQ�5����T�E�8�ʕ��c�ɐ���zs�N�x������cΝ;�V��1/�c��ժ�ʕ�NOx��!'�GL�S�������dcģG�x�7xᅫܿ���7o��hC���Z��_�~�q�v�Q�RuBh�B�;�My�k�}b�pN��=Oyr����s��2�݌s[7h����aD�8e5;�b��>���.<U��Ti���=�p[��GD%6�0hh�lp�!P�s.���}d�7������}�ִ�������e�i[\k���rxx�1បMA�"2)9���'waUcIF#�o���ֆ<IY���*��ZL�8^���o�;��>���ʒ��n}�9q�<�Ӷ�~w�˩�_]�E�*�و֔�|�!���qN�@-Y�YE�O(W5y>DM&�._�|����	�/��ŕǷ����l|�1ʠl�5��ZH�� ����5�}-3��Ya�n�EH<+
"#(�
G�:!�
[�o�N�]��
�'#&����hi,m$�מ(��DE_[�˂Ţ��#�8�)IMKѴT�E�%�ڶd2e��H-q�ߒ��`���@CHS��0w�[�4f�\�d���H��ŶUHb�����4�\ʲ�VCk�gU��*ƹn<ꂒk82�G�>a%k�b��H��Q���e&tW���'�a����Eh<5+A���Cϳ�u�4�w,C)�u4��"�1���Lz�v69��1��l��	E��8G�8hGۖ�x��h@��,��� ۚ�y�Pw��c̺�:�܂m� ��H麹��<��Ͳ֒�������~��d2 �Q .J��R�c<��JM�B�`qĽ$�(J1��C�Q��"@u����Z8��:X���L�hmS���b�i&�;���8)C1�;d@�.�����UI��zy�;�Y�5��|������]��Q�$��k�F+I����c拂�|�0O���]�߽�4����۠��$u�h�
�^X|[3hI����8x�ʋ�����K������8f����*/+V��ܚ�c:��Rۍ.���QN%�,�K�|z̤ק)n�_>�D}��T%}���"�=�,�ـ�J.Rx��&�s���-!����ZK�B8�z�/)jK��DB�ZK�c�o?��bI�fx�X���$I(��sX�X���UQ�X,������yvwwё����uܹs��l�����^{�5<�GQ�����c��V+vwwIӔ_|���!/��駟2�L���`�s�=�1�{�)E�@J�+���`0�Ν;�L�iJ>3Ce=��w$�~�w~���^f5_�)k� h�~�����ξ�{"%���ST�����wBc˦de-a&�� �.�����Z#TL*S�R���US#����l�>����N�����:͙��t��j2��z�e^՚�tʽ����6�x��U���<���9�{�8�X-Y�4z����ܘ���ӌ�,�W��[ˍ�Oxn0 �c�4Cnl���i:�k�A	��/��y�0��b>;&�;`�d�)s��u5�|J~�<NKʲ!��ap�ɠ���7y��ߢ��l�(Mp}��	��⩌�Y���.��L/���,OI)����;�sxgqH�:Kme��%���,z�+ޕBz���Dz�N0R����7d9�:�غ��E4�
L0�Qu���yz#��QU+�HS�V�mM�d�2dD(RM�D�eEY�H)��$��ۆ,	�W��i��6%քF�i��ӏ�L&c��<Ii�E@��G�;w�ꊕ�t Ƌ������7��7���2x�O�A��Ҝ��>������a��ģ]�E��WX�E�A�dI�,�$Rk�y�!mZK��:���N�p�!��!��Ux�*�Y)u���VV˂�Ɉͭ	! Ó�}z�q��II%h��(@�y��5y?�gJ2O�n�t["p�:%�b���FD1�ɘb�R͏H�����A*b͒<Kj��1%%�٠-��L����8<�$�LN��
g,���~|�������MF�1��,���p||�1��X���1M��l�aY�E���K�e9������e�
4Dk)σ�9'��ĉ c���`>�����)���TOu�HO���:�^��H����C�+�l�1�#�g�ZK?�Qm��#��Ru�����A�G
�R��.�TE�ư,g,���T���!��Q-o�H#�/��&�4H��G=��|]��Ж���]R]�6aD�(��
�*t�.]�����{�����o�,\�~=�9>|����C>|��0�9>>�W�^E� �;::"MSv��f�;8�����`��~�����I�,�K>��3NOO���bkk��������s��}z���m�g6��9���#��߽��tΥф���osq�"'�s�vm%���RH���$��i�A�`�RT+uC�Ċ`~/�rw"�%ZJ,�ILݶ�MH��c���Y,��Ï��\�p�X�P(5�{l]������=����t�M���SKY�I�r����2�Ͱ����$��z%Qa�Q�h-9jVԍ�ɝ|x�g0��7����&�>�\�g<�������laM�����3����,R�p�)I���$b�I�I����Ɨ�r�Wj<${a������4O
���*�,#Cߦ$Z�`��FaI!�ru���-���?��}
��0�gk�~��i-C�CX�ݿ�.�5��� �%��z"S��h�%�#ʢ�*��4�\H���p0fZ5���z��v�=����F[�HGC��P��U�E����8$N:CkjBք��cj��DQD�k�
��&��f ��&Ob�4�&��$�'�Qۢ��M,QU�9��1�3��'���	��\c�#�:�Y��ERx�-����W��=��[�&���w(668],1.���q��؈MS�jV��K�W%ug����X	�i�%Z�X�q�D�;�y�Zi�Ԡ5u]�*�MI]E�\��5�,"�2�1E�j��Z���=�<�z��-��!�ш��1�b�E����^9Ϫ��������C/��iB���F E����^�!�^]�O�%�BRUa�@k�28V�~EAmy���0��N�|�;������������q��M��(W+f���)e�eyG�mKdI�9�k=mՒ&	
�I���q��#n���b�$�6�&lll����IW��`$$��K;#Qё--�h�R�lD��xGٴ�X!�����ɈӢ����P��mT��y�s��d��.Vθ��(�QB��ka@��
/d�0����<�x�JR��8Oy�����Ƀ��=~���,�Q�%eٹ�����:¹Ё���}��G��gv�Ʉ�,�����u�V06r�H�y�&J������F,>��#��7�N�쳱����c��>RJ<x@]����럲���s���։_���_�Ī�Z>��K��� t�0��ؾ���x��-Y�O����V�4�8K�"�T��T�A*M6�3�����>��%m�(J0N�c��>tC�cr?��H�w�=�9J[A_��S�� BE� uL�+N����~����o��H�0IG�^h����t���X�YLg�'%��$D��dQ�ko\���+�OBp��m��,Ky��1m�ppz���6
Iq�`+�`+�;�	[�[\���.����8=>d9/8],9�?�xz���-�l RR�*�1!�\�<�����V��A	M�u����4}�������3�[^���!;����߃Yt��g$d�)y�{���f`���Iޙ|�,p��B	�Y��#���pጲ#!��Z��ha������k�3-���������(�<�Q,K�G���m0)Z��ٌ���{�u���o���n3�CB�b4$����Z�BQ�!9��2����{�z���y�ˠ�HX�$�� P�c��`5]�%�c��<O0������L�p��z�^��i�vv}%�N	Ak-:(-�������S�S�ɂ���3���+n�x4�Nb&�J"�����okQk��a��U�~�8�R~����� ���'y�[�`ƭ��9�9�&c�+&����bE�4��a4`�`9[�#��60�>˓z��#��!�/^$�Y������iy\��,HJ�D��hK�ޓjM���f�>'��oVz�V �?�RBvz�4�F⼣?Pac�����ѣL��	��.2��\��ʡ�*kH���l�1-u�P%�V�͂T����j5�C�qUI��a���*T�
՜���ϱ�:�Hǘ�YKs�Q�RJ��9�Q��oQQF�9Q��h��N`��2�"�J
�������w~�����7��*�X�O��34��y�[���T���힋s�@I��AS�٬x��{�7n��Cd�I��<��V&���m`���Qｧ�k��#�9hE���l��w�w�z�*��c~��q�����P�9KQ,Bbc������%���jɃ+�*����<�֭[�9�)�HӜժ�ƍ�9�e]���/��֭[�n�m[��x�pzVk�����k����f�x��̖<޻�d��n���bDc�8T��̪����\�x#��F)����Q�����;wʯ(b�&T�2�8Ꚏ��j�dI:ء?q�����>����a3.^���4m�5%��ٖ��}�����f��kX	�I���kW����mZېnL��������ҕ�NO������C�ſ�C�<xğ�?����x4`����	H��Xq��Ü�t���'�S��t��h=Ҭˊb��k�1-��%M�ơ3����>i�3G۴��l�#�/�Ls���_�gV�?��aǆ���N��Z������Fl���j�m�u���t~,B���<[����-=y]���ޘ�Zp��b�ֹ�]����bM8�55�ф��	�q�qLY�=!������������?���q�c�m���c�:E�	ԍŶ�҈8�%��&y�sx�O]��ߪ
t�fض�b�C���)�Q�s��lN6H���p�k��ʥ��TIY-��A4��Xk��t��O|������\>2�0����VHW�˚'����y��e2�d���X���mN{[�uI����1X�q�ଡ�Z\�>�YD'��6茭3Xg�5A� kI�'���5��}���Y��4��b<����(��ff���`��2��{A?�^G9Y�R��o/#�)*�)��]������qRSC9/Q�)/���'���5e�]�G��,a��x��=K���C���0n5Q#�"Nc�eY�0�uG���m�i��{���w�����is6�[H)y��1�X0)&����"ȰNN�����!<ԗ5I�YV�4V��(뒺���mQB�9yϘf-?�Z�zdL.�
W8�MK;������|�H��f�,O�`��p���!��/��M2Ss��X���u�����g��g�JF��l��B�"��� �3�!$!֦F��aQ�ˇDQ��4�E�%E��JS6�,«�!8�PTU���>�CK�<e<�)�n���    IDATݢ55[[[���f�w� 	Z:�(��}l[��O���N4Q�%EQ2h�p�:W���3��?I����n��3M����
g`]4��$�����ѿ�g��$�'�[���[��P����]5XcH����������9ݧ���F����p��5R��A�u�i>�vΣ�
��>�7k�(A���� MJi��&�u�����8�/�3Ff��j���9�{§�~��/oaL�bU�(WHeS�Z��bVM͟��rtt�����(���f���'���7H�W߾Ƶ��Ai[�0%�"	ӓ=���a�Z�%\}�2Rx�'�G$Q��P��Z1����J�YN�(�#7-���oȏ�H�J�9��Е���K�|J��� @����G��%�{?��?A�C,�{�a!��g�O;��t�?z�����H��Q�8K��]1�Tձ�]>��#�>̺���ޑEnMU0����&��!<j0��=���ONH���V,N�FCP���}.x���KW�������������7��"�-��$IB�F,�C�g��j*L�t�G���u��L��9΅�&�b�6'��gkc����)�|�)Nkvϝ'.O8�O���H��H�����1�_�o�����=
� �����xo���K�	q1z����U���_���������	�ɐ��VM��	j�072HӔ�l��t���m[2�O)�%�����k\� E��.��L#�E	����VJ�	�Ci#�/�e9�	�8&RQ��V5mݰꒊ�ց@�Jj�i��;�� ���Kb���-RE�ۜkHz�Η�"���`����K�C���I�����1-���zc��8T��&�s�1�8�;,��h�h�&t�³���1��tJ���5͞�������kWy�ګ8�8<<��͛�~��κVppp�'��`4S?�G(\�tD�F�!JȮ �PB�%�A�|��&���ހ�P��KlkH�D�S-�l?w�w��=����'��R�6�~�|�"W�K�R*�|ِz�n�](��cE�ȿ*���`|��H�����z�:t�Jw邖X��xD�}�W_}7� ���Z�Ҙ�}�m>���|���|q���	uc�m0eI"��d�m�Ui�k����_���mNN���H���[o���o����<ǜ�Z���$��PI�d-�)���i:��(dY����"�y�w�D8 �<�m[�~j��6��f�u��ٿ��y*��!��7��'�L�\FKM�k,�s�T���(h��	��@c-Nz4a�����Y���c��b�ν.��|�0�EQ�"��do���mSq��(%x����6eU���#?~L]�`qt�n[�a�)�-�L���'S��$h6�}�O�Svww)�{��I��{���!�à��)N
�����:>LY�#�6��CڦĴ5�4��&4�P����Y�3���{�'���_a�fQ,�sMJ���T3z�6_�o3�?bh+v����\��������z��]����Y����(Uw���S�$�t�;���w"x�t�<�ΓMf��]�z):��������eK��)�X��B�Z�޾���e���;�޿����[��o�+�nA�,XU��Ucp^Q���љ[�i���H�|h��84\��.p��E6���L�S����F�)��/0����uĽ�z�t�4�ݳ�{��G��S�^�@K��Ax�V �G�l�1������$��w�6ΑE9��Gϧ$IĪ�x�4
���/�D<ass���'Oq��F�1��;�N�|�����p� ��i��DJ�f�aS
a���#]��+)���F2�L�{q�ţH�gB�gyp���jCGT��IM2�1�t�$IX=�G%�Ha���3���p��4b����'1ҁ�k��sf��U��px)0�b��u��hD���Ѣ$az<#�^��®PŒ�j H�x�y�Z�7�3#S7�A���(�5��T��|������/��ZK'�,�'H/Ϲz�*�^��W����!G�,�K���jU�>���}j
#���i"�aJ#/:���-=��U�@(���s��}^��2I�/�Ll���)�	�T�Sܨ�T1Ac��&$eYyv�B��Aj���lHrG�3�$J�ذ�t0p�[��eBop��J1�MqB�\�ʋWi�`4�)�q��iI��Hil[�d8��D�]0��{&�	/�pu=뭷�{)J).]��l6�'?��z���/�ꫡ({��>��k.^��ʕ+x/�}�6GGGDQļ˼�������{O��cww��h���^�.�loo�����8�B���e`���Z�u��9�����7_�7]�Z��g�+Z��R��zD���V��&���u�eEU�鱀	�U�{;_
)�z��i����ۅ�8s�s4�~�pT��O��MB]W�4��-ٿ������QT��S�L��~�t0`���"T֣2��7���o�Xl��p����h��_�����i889�?����V�9�������,�S�X �f��f�,��4���1��Iv&�8o�ɒ4�u�"��bE�ִ��El#��1ތP���aж�C��y�P��x�xf�%:�˳����ڟ]_����U���*��~M��;C�TǾ�;�X����Qk,�e=Ԏv�$��$S���K������7���m��p@?K�����s��y���ӟ��o�������׿ɕ�_��O>�����/n�fUդi����"Nr���xՍUگ�`�qD��g0̘�Ɯ?w��`�1�����C�'ǜ�ݤ�si���=�|t��U����/�إ#���"���ր�h�4I�yMS�]�b0�D��4UA�D�~��7H�\3?�K��E���UK.���x�
�=�b�"���d�ŗ�;���8w��'�i���y�bUc��H8|d>���X�A� hp�lL��w��xs�������%$i��=���x'-�~S��i�Uͩ)��t�G#[r$M�g62�{\�5n�1s�k�Z�i�dЧ�����Y��
ǩ2Tq�o�'sJ9%�,�H0.8z!5Ά�6�JZD�Yo�AG��.DD��![�}C��4F������.q�ʥK$Y��{�i�AD
�Y��j���w?���c�Tq����p��s���6��p���X	�����@��`��ޠ��"�ؖ�*zy��h��KxpD.43q����s�������q�[����?����J�d��p���U^��ߧH,�pA�5�����u�Сx�0gH�;K���Kuc� -z���p�u�:�4ZR5K�"�̠2GQ̹y�s��%e��Ĵ�~z�3�n�E��8 Q�(˂�>�)�N:c� ��x�">�a�D@0y�W�Z�����}�5��9�4����e�X��o��{��t:%���ı�x�s{ss��տ�G}ă�Ȳ�7�x���-��b<r��-QQ�q-�Z�
�vSJn�2���<:e0�����]��!BK����^ �YO�i��x�(��0��8o�Xİ������h���	��YU����c*�vI�)�Gl�����_���\�%���A��I�mjlQ��hH�899A+A�T��8R��>�|й.�l�����?�{ϻﾋiK��~�~?�O������V�u��A� �d������a��ł�bF�n�����틤*	Y�CZ�H��?<dUW�Ȣ���(�T%���HKo���i�A� �xn�<�Y�z��RƯ�
[������ub�����mAk��φ���`_#;&�0�2���=�%YY��3D�b��9
',�������
�$�R�s�����h0h�ZO�kT�����u&�o�}�*Kq�a^#�g�۠��Ű����*����e�x�d���}.��pxP����5o����:�Kݴ$��W��u���nݼ�g��Gwo1;=bY.)}E���QFaBc�ǶQ1���svv��<��,*��Sݿ�3-[[cr}��M�������'잿��t�<�8�`Ψ�B��6�^����""�!<6�rnS�!��I�S��C�x���#�Sc��I��K� &�&�d�ڛ_g�KDYΪu�H����Σ����sxx�������0ZΠ���Q�`F9�L����BG�$�G)��x��p�b��s
g��(I�BZ��(�
�$xf�E�7-2�G�$;����o~�C�r9��>J4ȶ���������%�4�h�Γ����i}Ki�x�! -d�>���"���x��F@mY�!�9�g�I��(J����F�-Jb�����	/^B��Gǡ�Lb櫂Y�"�S��ηy��KE�ݻw���g�e�iEX��8ʲ"MS�7���ZY*i0q�J߄Y��Ғ�1��&ۆ�!ᡗ��Ä�K�G�w��?�_9�CړS�?|�Z�99=B�.I�7��,y���=�2T�g3óMI�O�w??��E	]���g_sNf�mŕK}��>����YLKz�^x����_�%<@J�+��z����tg�a�t����/�ļ8��v��ڎ����.YQ�w����/�$I"vww���`�
��~�3�1�ʻﰽ�����[��g��hĵk����Y�}��ty�s��V�׮]c2	9�B��!���'ؚ��3������&��K���� �J o��E$:���(��T{	�$z>��5�p(����(T�%�e�bX���/�,e��`��h}�P �Ƕ5����E�1M��t�Ҷm@�@�y�B�R=�%[�ʆ�l�䓏���px�K�/0���ύ��E��d�m/:d�������^��uX�g��Q?���'�b��D��m�����c6����3VZ3�kN�!i<a�RJ5F��Gf������T�Nr^z�U�_{��O?������Y�h��:��v��K����9U>d�x�B��r@�6a:��U�ܜ�>�P�3�{x*-;�p����_�,��� |�4�\Ŕ�9�K���7��+�u����=���ͭ�?�����l������8:<�׾��\y��.g%�J�K_{��^{�f9eo�	����GOOY��óu�,���0�������ĉ�1��{�<�s���#"!������K�qz��'���4��w�r����������h6|8��
���)��It/'��ՠ�Kb욍�����`;I�I��x̋W^���W �4�^R��4�H�۴ԫ����'����=�?�!��)YSд+h�.A)�5
�C��:[kt�#���ŏ����"vFی��I�g��Y�qR���Y̧�M�����1}/X,K拂����*q�y�1�"�L�J2]-q�b'�T~��Fi|�R�JVeMދi�f6��;������]��ntg�`/�k�^"��6��$��/I����E���Ƅ���m�2�5u��>��s�y�w�4M��Ѵ5����f�eY0��*���	pf����lBam�~
��� ]����Ja��4JqV�\�X��4�#J%'�f�[Lےf	��	����?�}\�I��y���}���IO�����{�<���K��_�Y�3��k��c���Ō��/�[;X`1� �9�P\_�����=�]�]��M�JIʲ��@��tDk���(
666x��w�L&|��'ܾ}�8�R�|�u�B�y������\.���y��!/���Up��tC��)˒,��㰪��}�6����b�6�9�����1�(���ϲ���_�F�� �;�8w�������c�K����>�/b��|4
���5	K9�F��$���Ղ�\�kG�Dy�_V8٠u��Sƛ[��e6?�µx2��
�!J���\pkt&�AX���iI��4ɂYS��R�e�`1��e�1Н��؆8�0qL�̷�Ϳ��z>[���S.]�lP;Wu������7R��8gܘ���h%0>D��y�k����[T,�%�y���ﲽ�2�|�%T~�i{Don�ӄ�����o�C��zQ :�;/%V�.�H���Yq����S��/~�3"��gy��L]*�DT �:'�*�^�2X,�����z��Ĳwz���f|�"��i�aV�X�������c�|�-^�,fS�vw�1��'pr�Ϡ?�-N����'\�w�������K�(
v��'\~e��^ycCfD;=�B��$a����Wq��gkދ�3q6���8兗.��ք�~��߻��,e�Z%q��W���\������P��ŀ��<�m�$ �Y���^K��$�R)���C%�MG/]z��<��˂^�'�4��xƵW�Kԗ���(9��KR�o�lE_�X�ǹ:���/�^#�F�'D���7�dg�"�Ҙ�2`,B�;c��S�OY,g���lGV5��);�F6�F��F�؂��xԶ,��9�X%�D��j��VJN���W8"D��:M�z�v�I���wn]��SBwDg��\,
��jQF˺`�Z���׿�2�_��d�N�����ɓ'ܻ}�4��{=z,a�a>���a�_�%����/?��ͬv(����4N�R�V4mI]-�B�&���)�U��[O;]Һ���Y �D2"��.PZ3MPu��Ƅ|8舆-V��4�TD|�;������L����=�]�2s�Hy��o����]<�+��]����[_0��?%�m.�Tn�s;����Yv�y(�&<'�2�4��7�0Ԅ��%�/?�T�T?�C����h���t΍Bj������t-eY"�d{{�o~��c�_��g�}�M����1��Or]���,wɽ�P � .�(J��m�ew��ݫ�=33�|�鉙qD�������l˲H����J,�^��]�2��D�1�(���y�y��>����N�C��\�z����%)�sf����M�]�������T@tFɯ(����ѣGE�,��ɄW_}��/.O�q8��s{������=��S�Z���N�< ��Y-��dq�A�����s��-6����1=�c6�$��Y3+,�La��#/*�+�}M7]ź�aY��'$�q�"MS�H/�ҘR���:�����6�MGO��b���)r2�����:O&غFᩫ������&��\@Jɝ;�B�Q����6�/�ȇ~��ppp�x4BIIEX���b��K�C��E���|:E8PRb8,�RH�*�5Q�غ�+ͅWnp���tё��P��ѐ4QĽ�� !;�C��s�,!DCr�K����������nQp�o1�v�Yÿ���b��D2�8�|���|S�7��V][r�������M��9�v�|Zpr����X��d�y���^���(�#^y�m�/�ȧ���'����⫛r��1[�/r��+����]�i�k��T�V�CUQEx�L������Ib�j���1�%��\��˗�)�>bv�}I��-Q�Pec��k���a�F��Ra9��}묣�̘%>RD&�M�.���b榢%,q"�,$��.\B )ʒV��D⫚n���r�S��QIJm���-�����Tu�}G8�zr[�:߈�NQ 0gX�[�|�.\�������"���u��J�"f�n�մb>9C,�{3.薚pFQׂ���"��Ŝ��ڔt}�����E�5VF ���6�z���d�����\.�_���zޟ��ߋ7��52�t�-�8bg��_���/���%J�(^�����F`�ct6^&��yN]�R�ISz���zm�|>H���ok�N5緷�qrv�� �oБ���'DiB�ա7�t��1�j/@y�EAUIV����B�M�J��b���I��˯�[�?"��@6�I&%nrL���Z�������jJ�f�w�~��lQ�6������ڌ_�16,O��M1p �I�&	���t�:�Mɪ�k�n����6�_x�?��?�>`6���Ӳ\���,ј���Z��3�]��[o��֚�>���?��(���z��	^�8M8���������Wo���	�v��|�;h��}�6��n�����
#��|�!�v:�.�����cn߾����~�~?��Ӵ(��b�s"-Rt�����������	���8�R�V�E�E�1�� x�?=��밹��6�    IDATF/!i��X�l�h<�w/p8������}�lĎ��V*�����M'ċ�Ӥy6I(�F'1�� �tK��ݭ.I����Ez�.Y�1��{����!�,c������G8k�$1��c�����q���,�(˒[7o�}���yI;|��_�ּt��|���++kıF���N�G���	d?Q�F�����Alh}��.g�����/|�[T�S?���_~�y<�*A�oQ������ti���)���ry/�C����g#_����Ιl���Ͳ w�z�����mF�W����0�ɜ%E��`�)�צ�m�֚���#f��w�{���ֿO�� �S�[W7�������3�ߧ��9==�l�t���[��ӄV�Og�O��&V��fU \���>urDUUlllp��"I8z����>�A����}��+��}��.zxF7����G�^�i@Շt̠�|vU�]����}h�J�D(�8ąC֒��_���c֯��::F�1��Q��#V���E�덠�4�P�v��1:G��tYU{;��TEN]D�Zi��AtЀ���/��xO�,u�l^���)���^[d�4��*�$�-���|6��,C:C5�¼ħ^J�N�Y��k����
Ó;���q�$������o���Gԋ)g#��������}:��b���L���AΉ`)���|<P �8jkh��ٌ|t��k�����U
a@i0u��5�(�����Sf�)Q���0^X]]��UC��8:9�s�l�����u�g'CΝ��ښ'O�P�:i�3Z*�^�@�ߢ25.�T�X@�(�G(���ZA1��wx�xfy���#�����rV&\|�:��&S7E�v���w�wo�^x�K����\�DQgĭ�ސ{?~�G�JK)�sZ)$�d%��->��V���\d� r����.���m�.�X���|��ʀv��N�%/@��yN����1&jR�:(-������+��\�����m����,�BMk<x���1�{�\��R���C��͆�������z��g?`gg���a�X�(�~,�:��^��`Bo��θq��Ʉ�d�J�5���V �����.��ߤ67�F�~�t>G�t�r�TZ�f�Z�F@Ƿ��x||ʤ3hEt5$*A!���FR�u��V�Vf�eY`eC$kDJUU��x����!V$�6��c�UiXY�r��K�x�4n�Q�����իW����?��ʹ�-����#��t�x$�<'�����F	+���X�^���ʓ��R�Z-���7��Y Y�T�4j�(�JG���)�$h=�$"m'�Z��ǿ�?�nt��2>�O�����r9Z!�5��`l����/"C��6b:/�Vx����O����떟�9Q^�c�����8B�ָ��~3�4Im`k�W�W�h�7�s�4����������7��\&��R�錼4H���;�`k��~F�I����A{�׾�[\�u=dxvB�g�m1������p�N�bO�53/(Ua��\�ܹs�Zm���۷(f�I���ֱ��ʫ�/Ү����o8��3��P��q;���n,�a���K��)���~w���|h��E;_)4�X������}6�A��S�8A疸.&���2>;����֊���xvJ>��LE�IH;1Q+�����㓧�.G��	:��j�S�F�ݬ.�|1%�D�XPU9�d�|�016/1��/!j��Mw$[]��ed�c��QL�S��:�w���v������O^��{��/]������8�V)*TI���-�|8�2�w��vD,e�T�:Ո
�ٲ��(Tk��	JFA��=Z
����Ni�&\Z[o�2G�1J�N��,o��I�CyCڊ��'�QJ���$�qqL�D|y�.�����T�f:����Q���G���8;�Q���v�urS�p�����O6m+k��m��0�O&ت��.u;�(bD�K4���n��!q5e���Ӛ>%���x���_��9{?{����a���7+�.�/`by*����s�E���k!�M�K/��}�p0�H���~ ���.������=:�.�^/�[��CG�YteP������(��,6�8\�ũ�7��fee�W^y%�!�<|��=�ϟ�ܹs���+c888b8�R����I[A����+D�8.Z�.\�ʕ+lllP����"��]'Z��QBЉb�o���]ǘ�7��=�5<��OhiI�k�k��V*]�q&'MI+%�. �#�Z�C��0�{J�9+3"WK�$�#����챵1�֡�d<�~�s)q�B�{$*eug������_$J�l��&I"�Xb�EHI�j�Mg\��lop�����p�i"����_���㝥�b�iG�4�<��rVz}�����(;�t��.e��)JK��	D"h���AVfD1���:���>���ɐ�j]��.в��d�*���ß���&��]zZa�u�-��5�/�v�#�[�v�<�w�ܜ
W8�I^"�G�����C��J�\�(�n��`P��I��NQ!?��ZA�\��\���spp����%~�Ο���]���o��.��
�� A�׸p}�g��c�_���wɲ��,�*���0��"bI�������jwy��1}�	���\��0�k6ϯ�����
���_��ݿ�5�It���D� �5���2� ��8���|uo���
�%t� '| "96XA�)e9�[�N�(��ziHkC��>���[��ھL�t�e�k�O��v^��DQ|�z^����ㇴkCG̽#�Ԙ�B�
g"��i7�?)QJ����ݿ�Õ6���6�ZF�G�+�z�<u���Z�ݔ��D���8�PM��l��f���HDGSaӍ��%B��s�m^�7��ڕ̾����Ԁ��ר67���7��{����È����w�@ٴ-��LJ�s��o$2,҃NR�҈J��"�c�ZR!��p�O�Q�s_`8�3�8��c>:%�F�V��ʀ�~���\�|�V�"�cV���}:�M踠Vq� �E��!T�|7N0��n���ft�.� ��G"�9<<${�ǩ1ȭ9���i55W/_acVr�������d��.u��QYA�GDV`2�f����"��1i\P���d�{m���_�#��Gl���gAh�P5��!�{�W$�=^����/��l2��}�U�"��.3�v�?�����98<���n�Ե
��\
0Ue�ȣ��`m͝�����`X�K��bc��D@���?�ɓ'�9::Z���ݻ�d2Z*����=Opm28�<�C�p#��N����)�|�	���!��>Y������O/��xvm����?}�/����G���������F1�٘��kyO���F=�tM�Ą$B�[���R0�ft��*�О���I��`�DkI� ���C�-��g,V8�|��k�Q¹sy㻿�΋�1����Q��Ca����f���\�>����������hXy ��u�QE�s��#U���I��BxAmJ�<��Jɲ`�L���`@�nQ��F8Q5��`e�)F8|�B��X�NU@��3s5炈���[ﲙ���Cq�.z���`�![/�C]=G�f���,߸����������m�k��}b�\3W�E@��.PDU��C��y���oZ��>�>�J
YPVSV���1�Ͽ���A��`��F7�ŃG)�	�o}����y�������-u���4i�Fv�VƔYI>ͩ��퐊%t,n�/Q~�ã>��6Ov���3���)��x��W_筷�`��9~�>��,c�#�P�+�ܐ&�,R�&�N.�/_-~�D���iSI��!�7�	mn%��eR�X��A*��E!�"��g�5� vw9�.�}8�1�`��CYS���^%`+�O&G*4$r! r,�:��%�bL��$dy��p�����@h��t��0�B�#�
�%���oI����y�p9�ռ����SqVK6�>y2�x�eV��H6q�o�����T	ꥷx���|�m��� �����#�eN-"�5JX�@�7��^����o�-��"�Q؂4��V3���t�k-��]�û7��j��铯Ȋ)E5�#@Ǵ��_����}^��2UQbˊk���%�̫��x�fܡ��R��#���t(���L:}��YM��T�2ܽC5�qy�}z�;:bVV�n��V���w�w�vS��\ȧ��s��L/N)m�j4B�eȍ���^x�J��l>a��"��z�/�*�����c��>��$�Z@�P�LAKkj���=���m� �fY�����gI玳�Y]]gG{5�s��b�ּp�����_RW*ҍ�F��ڄv�1U��P5�JG�R�� eY� �&���8��`y�O����ï��~�芪i�*���K�\�,2 Z�'''|*lJu��u�撠罥,���l�pL-�6˲d��ÿ����+9��N��I��;L~/��.Z�A��I��%4Rh��0��D:\lY�c�*cs�Ɍ���}E�E�,������^�d-Q'
Ib+�y���4���Uνx��Ή�B�t$d��2fv6���c�����^#�������C~�����*�
�r���l]1�GTU�4_X��JqF��6R�β��2�:�pUQ�DDxRDK�W���NW�J#l��1��l�)+�q���_�;������I�q��������Or��C^z�{+]�o}�R��J0P/��" Լ���l��I�|�X�����{�Q�[Ե0��
�S��b�a R�:���&��zK-!�����J
4o>�DF�����HA5�~�.[{����Ѝ�>�� ���.�{�L�>��1�?���W^���7��؂HC�ѢZ�rA����(��V�E;iR��L�9�}���._�?a4���Z'e4��Em�z�U���������w~����n��Z���O-�l�atx<ZI�gJEH��$1�����zQ5��L��<W��Fh��$vN=>AۂY1'k'���ߢ��p�v6D
I"BEl�[W$�c��2��5�_�ehwyI^[�*�D�I"b[���T�A���9�l��zCe@[0��BE8���
�=ڋB��)FD8g�J��]�кa�W1y��R}����tDLy6��sV7�`
�)YG�GUԔE���.�o���o�6;�����^�"�m ����T�J,����	��F��V2��q��4uT�1:q�6χ�
�W9��>
W�*Pi�JUT�a�
Y�̊������v��7��������!�x�Q�1��9h�+I��(�"8�󌕕D�����2/p���`�YD^��
�4M)Ƨ�\h��� =J���
qg�{]�"�Ԕ��m�(�E	ǶF�6����q�7�5U^a;)�|�Њ�����\!��1��������#��xe�-?��IIU�υA��.d( �8
\g��#$^:�>���>�CZE��`S��$��߼�8���[d��P�h����� f-�_��\6�/	�a�"�QJI�g�}+d7�*0��B;�H��yh-��z�`�ѡ#��[ڸ��~���K��9�z�4^�[�Y� C,���pH����쀸��I����W��޺ER�`J����7"�pZt��^d�8防r�EM��gh��v��|<�ٚn��R1���GST�4�ט�f��Ǖ5�Z]�T)�.^�_â���{A���.��O��'�p||�J5��
��g���a2AՆ��;Y�P{Ls�A#���A&�.���FM״?X�;M��H���n����:i#�Y�H-�Nk���jK�=�5hk�8�D��fT�\��|���(<`��Y��^�q��^����s2!N���2�S�ʠ� FAGa��)t�>Ѹ�\325� / �Y�b�=�E��� s/���L��8xu�	�q7��2U8�+�h���K@��:�,���Ŷ��������/�����Xc��A���p��h��������p�/_}���sHS{K'M����<GzOn
���~:��}��S�s����$�8��Dq~p��s\�q�����or���b��mV�hyo�X�D�7y>�p�l:`�Y�DJ�TϮկ{h�,B��k�˓Sxfi�A9���@�1饫��?]"Mc*]����k��6(<S3�.+�"���`��,�[u]#+KQd8U#&��?��٣���b:y�1��(��/�nn "��L�?�#z�:�>���-�6B�3��(���Gk͠nQ�6��!:k�Ce%����(�)��^�������+��~��>~5��\z���-2��g^�O�ᔢ}kӜ$��zRV��I;��Ւ��k�}�ll��4�
+j|�q|i�t̅g^���1.��󊲘q6qZ���㏨����qe��SVP���&����t��JǼ-i]�d^��f��� +��,�H�iQ�������t��!C��!tD9������N�,2ј~�du.�c��������G��o���w�v�!�@:��Y�s#bUQG�Wt������A���c�H������p�CVx��<�5�H��a�g�H77�{딓��d��qL%-�����
S�h%��O�!d�s�rc��/���Ο?�]YP�(�(
�,k6�`WI[A���Y�>dY(ƪ�
�p6�N�CY���EX�r߯���o#B<���Dc��Cq�����������V,�;�vUr�ע��G��6��baF�H'UP TDQfL�a0�`�b��Q�t�&JS��1�|Q��)��P:!U)Z��^K��%3����|F;�AFH�(ꊙ�X��`Vdqt���![J��v����l�l��G��8D�:��̐q�5[״dh�[!�J�k�A�������6/^�N��ӣ!O�w)�"t=�6��k���M��sw��l�ۭt����i�F8G�_e����u�����y�_�+��O�ՖK��}���}��9�x��s�?b���Z-����%D��F>�QW����<W��w7�ş�րC(���L������R�w1B�����MU��o0�!����HD���(LA9;c5��[-��V�물��h>���Gd�G��2���S����iwt�=�&+0y	�१rɫ�"Q1v:#^��"�l�Ղ��&��Z��;/s�K�������ݟ�qp��;b!)l�� �Dx����-�k*=�&��/Fi���F/Ă���B���#H����bQ�O"cDY���$i�j%T��B;��r%5
��M(&��x� �0�&�n!��*��C"To����Ls��!�Y���I�`�+?��l��7�6�����/x��;/^&w5Mc<�:=�����G�&�Q4�+B
'pVQ%�K��e�I��`���6��ul�6��e�~�0��9��3�����o�������{�^�����ҳB��-�Dj*f�q��V)�o����5A3	�T�@mI�F�KX|M^�f��3��9:9��V�Q�k��
��e�������ұ	����6�ֿ��$��<�I�(���I����
�Ut��&4fck�V�EYې���M�H��V�v�K�,�	;L���?� ���5Z�Z���U|�Ú�֤�:>�0��ɌhU7��!nїi6��9ВkԼ�l>
��2��`a�>��s�n|��W�cV֙�*���pt}:q����v�R���x�)�����MY��b-�>��]�v����0ư���͛7��/�tUUp�����dgg�Mloo�������0�����K���fs6loo����R���� �t�q��2�{���.+++���/�[Y��A %�A�B��f�Z-�T���뼴s�2���?!�ߧ�O�kK�����,�~�`�-��2<�Ե`^X�.l�	��;�QJ�Ɉ��	REH<�)�����C*�X�E̫	�)��W̟�']['7��dL��E��?�g��$;=����������5j:!��x6��,U*�V����M�5i��H��}AA��$ed-����ǿ�i1E>y��<?�Z�    IDAT���Ǐ�L���a���`���ee}�����?|L~�.b:#��`3�����R�lm�����g�f 5��	�R���c�����UA]���5!3n��RJ#�Yf�{�LDLCF�����u.������E����&1��'��\c��_I�
-$Z�M~�a�B"�����!��d	=m9��}��#6^���6cѠ�7_{�Qg��Ov��1�v������R��%1g��V�8��!u�9��ϱ��
gk�$�V�o�s�E6��ď�p���'�;ڣ�I�I���e��y�>�ǑF����%��H���"�"���e��'�JM8OUL0�w��'�Z�@����D��(�@/Z�@r5�EK�wH4?H�(��ģk�1�|�cGg�U�Ob�Tho�i�D�I#q���ј��������ID$��)m�ùMG`ms�#T�J"tJ��Q�೚~+B` a@���3�ftv����cz�?�W���JG���/^�������R
ur���C�t��N���]�Q<W�.��3x�)�)�W����g��B�Y�b�@h٠���&��NB��S+���6:v��$ni�`Z�UNm-^x���HJr⽔(��}6�/��<�t4%5�8A	IU[���8�25���J�����>�~%XI�[�C˄����!7[V����0's����GFm<QK"��:�p�d$�Dג�@�#�'��e"��@o\��:�D�SQ�E#�i�]�| �GX�� �PB6�"�p
mzTU̓aάv$�U�V��gr�+L��Oǔ�R���)�>`+B�|v��y�Ç�M�\�r��t���)Y�q��y�^����	�n��^{�,+V�~�U?~�o�����l��F����K���ܿ�G����x�7�9����8gȲ���{._�L���޽{ ������쐦)O�����#�����@Ol�BGtW�y�M���D�3�����]v�cZI�Œ>(�D�!aA`��6�`7U*�K8��}�@Q�0�%�tFUT8ch�9y@��g�|N5�0���r�O@�he��=e���n�J����CQTV9�����rt�n P�A����(E-���jd-�|Q(ڭ��:\�b����luf����Ͼ���TG�R��
%b�(!?N�nm�:B�hR'�5�C�ʣځiR���e�v���tksa�i]1.N��%����O~��û ��Ԡ��Ϝ������&k�A#���������" ��"|������i�����Mؓ���(�ä�xg;�[vKY�����l4��K��2�NI������̰��Cg��)�N�����&cF����v�w��$'�+T��emѽ>�+:i���;�/����z��j+b|�#��>�wF:>a�ۥВYz�
!�D.�@Q��xg����/��y��֌�սpx,�.B?'�EK3@1�R������/|�����T�Z�¡��&�SiP[��qCB
m����QXW�O�X��ZC=����XY�1%���3������Aq|p¹�y�����[�(�v�(Ex���=e=gby����?� �S��XK�l���OI��R���{\�r��/"�e]A-(��1��<e�~����/h�3T��LN�ty=�1B�E�HW�b��G<��9��6���4�(�� e�6���$�I1U�ȳ���J-,EQP�%�"'�𘼤�Ͱ���K�0��q���;�2Ҵ�+�rij��B��gԽ.$1�f�e��@D1Q+E�z��o=^EH������,S�'����"���:�p�)f����*$��Eb+&՜
�0I1�AH��XᰮFzq0��3e*M��<�C�6��~�Bv�HT�p��HEh������I���3�ϱ6�c��)E�Ĳ=����un��޽{������ΣG��s� ��� |��g�u��˗����,��O������˗/��_P7^}�._l���3����s�?���,y�7����Ν;ܺu��l�7��M�qp�G��r��6~���W�\��ŋdY��و$������O����'���gl\��|�[l\��?@�WdH����٩D4Q�B�E
t+�5]�y���3>�b�C����k��iԬ7J��^;B`�Js���O���|�����%�jZ�6=�G�O�0�L����+���3N����э}jV�H�XM�.�iM�uUQE)
gpUA,=>�%u�ΐ�DxCV�TJ0�	*邮(&�P�E���F-*E;���A�o�-��XR����r��x������ē{��2�(�6��z�5��tHup�\p�i��8Y��.�]c�t��ryz_�������'e�G���d��&q�J��F����/��퐍���8A�ăgU�F���v<#btm�#���Ɔ�=N��A����W�{���UIn
�ќ��(�2�[�C	OL��mZ(�\����s���.ٽ����O�}���0������%����|��҃�L(����kE�!{⡽�H�N�p��.�C�?��e�LJl����fԜ:�o��-�d�z����p�)|�B�]h�.�������/�΅
�����k�R�Z"�N�P��a���):vHW�?���K_d��R��<�P8C�l�h.�P5���R��"J2MQN"�b^N�*V��b�{�������{ȁF9G:���<; >�������o1>=c>��j+	�����.I��4�uTyF�QB+�2�T�'��ƴ-j*�i(����F�Q�X#����U�lb �|e�pTe��+"�	�[�"���u�U��R�N���O:��dg	�e�{����;�8������� ��M���th�)"�qq@�
kpe��:ziB$�$��0�2:Q��RL�}Z+mF�1�f7�[���`���"l��X�� <$J"����{�y�s!	�{��qS蚠^��Mw2)��i��MHj�n���+F�5�7�u��c*��<�����0o:�A#���v����߸q�/�����}&�I�H4���x�$ͭ1�Y�X��ի�y�t:�n��p�{����)o��fj�L���I���C��1���8o8<���㇁���kh�)��n������e�+�^��d� ��'9=����Y8�.:��:/	���F�KX����N �;-TQڊ���u��H<e���*�L��,:�qᵷ�;b����s0��R*@,�9|>��|aCH�ɉ�l2���ۜk��[]|�pRQ���V��~��耞R���j�Y}훰�FQ�h���i�I���V�VB�N(�b6Ǩ�n7��ߴ͵�P�J�2�4�r�et��
�+�qBb�g������-ֿ�J\h
�9�(�!X{�m�/s�;�����?�*$�@x6��u�8aD`h,X+�a��7�}�����(/�������y����"r�峬��0d����e�(:�mB��xv���B8M�,�s8�Qi�h��kC_u)�g�|tL|�>��&��$/�t4S�[�j�,��Aw@�
x�C�Y$=]��UE�z�+�x�2�����;����m����A�QH��1���9J):�����o��i�;�q"�-
���y���8x�-�_���M�F����=�s����%콞-��;��
;�ts�F�@ 	RRbP�biF#�������p��/~��eW�l�eY5���#iH��Dj�x���O�q?���=@��b�}y�>������o@'c-U]�3j�-O�+����	@<�5F��J�◴&�n�ua&�TbMYWh���[j�H"�%R{t�P$�i��cmC�H�@����x��l�~���x�����²X,P2�1�as���f�P��"cFN�=���,~P 3˻wߤ���[o��]��?��h�0HzTT�,v�A]��4�,�T�A��K��?�F7/��M�����i%������5����`���,h\�m�"��j&���1eE�/(�����Z�3��]*m��C�[kz�:�ID��@:��
-��-�$��Q"���(+"�HX,f8fؐz	�A*���a���r:e�װqN3/���C�,a7�qA�`��\{�*O~����;<FR��`*FI���@Eqh��5�[����U��Ȑ t����e7K�9�Be,z���~M�ST��90�%���E�LR�i(G�Z����� y���8���&Ukx�Q�>��#����g�������c2�`�Y"����B ������^������oq��%�6wZZ_h�_�v��~��A5n��U��n�1���c�՟��:,��ri��	��y���;����/��y��������~�z|B_;�Ё����!�l�	-`K�'Ako�ʚHxJaLM1�B:L��»p������'lZ���ϿB�8fqx��W^DF1��d=�(�Ai���W�ݒܔ8%�Ƨ��W�y��`��lX`p�c�z̓]�՘�T"Fo^��7���W_c��؊X9��B*�������D-;I"-�"M�%Dm2��B�Ľcf�Sd���1��u1T��ɔ��.Y��."2!I�z5� "��P&fg�"�l����	��=ִR��V�T�|��ڇ�z8�[B��{��O�D��I���Z�[�~H�����O׶��?�O#<K#$u7�n}��X��*AyIe���I~J,cT�0k,�VӠ����>��	������=�o�D�?��ŋd�}�$e8ᅧ�
�k&���w���oQ]����t6g|�>��#�U� �Hk���D��׋��� �g�-�-���H�:pʣ�X��t�9]��L��`�Æ���.�%���8뉥Wcꠓ)�/J���G��{k@
d�p�)�n.y�B��k���oB��x�ZR��=H�TH�if3"!�mg &p`���������F)�'T��Z��]�����5!(�9���G�J���hOO+\��yI�k�ї#^�ʷy�_�	����#�ه���i�+" V��P�9+�1w���G�ǳ�/�
�ϧ�(C��?�6�K�Q��7�n��⌣*J�E�������تF���OiLE����sv��/(N��%ɵ�����KeL�%q�9$�H3�C{)N�Ak8ֽ�$IH��ʪB7	C�%��dsD,*���G<��;D~�����g���p�`���?�c.<w����ܽ�����!�8z���b�/�@_�B�bQ6OK~,�H�l�3�-߶�KCӷ9Qi9YT�6v�T��7�����Q���:�T}-����9�T���c�r^/�������2�ei/��?��>s�W_}��>���b�|>�Z�h4�(
�1�D�A�s7_�ҥK�D�ѣ��d�?�)�?�<W�^�'?�	�Ν���kL&v��Y0�i\`�Mo�'N�%��r��.�RN���������\�2~t��H��$Ⱥ��IR���6t�TΉ����ޑ��bt�P�s�/��UH-@I�lB�6H�β����'��WΠ���P��'{��{���-�҈�^�᭣�'����t�</�![�����~��c�	:��W��W�xR�Ò��dD�gv�j�>�KW��A+�U5�Lh�U�8�	G#k�������&���{��b9��I����q��U���vFZ&w����b���pz�'����;�׷��^v�,��)~1Gi�O���r'$~��H_�8O��D=�LZ��=ۖ������Ԕ*b�,R%B`�tH|�RaX,r��Z�n�9�ЧXQI,4ySSS���Xd$�>Ʃ�볱�!�Ţ �����D)h��2�Qk�������f[�OP�l��|L�{@��H)�i���y懛<Q����!�N��bM���C��K��cN��&�n�����	eQc]�$�
mԀ�����jKj�ѓ\&�DI��E�$�B�Z5������g���UK����2�C�?wgH�p�=M�X��Xi���%m��������zAK�o���r�� R ��(O��m�v��>o�L��+�:�B��Z�sr%�3Xk-��LH���P5Q)��	IoH�OP�-���F|n�+F�/s���M� ީ���*�,t챥'�g�H����ף,�A%�X@<_J�&q��EM�T!(T���|����;G]7%7o�5��,Ǹ�5�C�kj��܏�4Qɬ�TB�D"�g���p��mE8Oc;Nv\Քd Gkk$I����� �8�rA�)R-���H�)��5���W��/�ė��_1��A�0ϏI�u*s��/r��W����9e|����w���o�*�׶�<��>襎���'�R���#n>���k��Dq��,��W_G6����>�|�joI��UJTOg�{н�R���\�|��z�����y��W�t�u�\[kɲ�������������dY����rk�ϲ~)�t�������������+W�E���[&6կ���c0m��b�L���}�0�5i��{p@T�F�S�
GT9*�!�Ŋ}p��UMԪFJ)����R�pZa4��P:$5�#��� �	E^���L�~ȿ���[D/C���`^�Y��T�)B�s�ơ�
�a�3|�OgL�){�f$QJ�B��D?����ˀ1-�t1���w���o�#hG"F�h�g�D��ek���ـ8�A�s,N�A0O�c,	Q���i-����8ez�}�j<�b�!�%����T�£f���J2H��cQ�H�/�@G�$ђ���s�b��P������n�'�����G	�0!j����a��9JFK�� !z�*�^RIH�_W��#ED�em$�2�I��n:����,�V$��9�Q��EO����H��n���-��cd�z�in:�|r���=��e�iS4�ƒhM��l�h8�#�QL?JX�Pk`���!$��pf��×�u�sp��/)��!t��9�f�q5��eWr�5�Cm\DuZ��D��SZ�������	��k��	� !�KdG� ���n=x�G��nV.&?���*j���,_��/�*���u����=�l��_�L��G_�h+��9BXFCM�u��6%��$qB6Z��Fk��N�F��]�q�-H-i��
����zt�Fo�O�D�Ǽ���0{p��6H�R��[74Qн.�S�x�`���C� �d�/h��B��75nV�Ɉ��P����g?c��^A�PZ��2�F�(H�갱�!��5�����#��H��O��rU�}D�̦%��
Elnm�J��9�*�L(�s4�)�'����>N���뛛̏y����)���-�������Z�g��{N~j��w蟿���8�$��G?�qZF��b���k;��(�q�rS���rE>d>������w�}�o�������c�^����_���i�f�y��9w��eoo��`���}��1J)._���/�LY���c>|�R�,˘L&K��b�b���W^��ի��{��tID��������n>���飏��������9�W����A��cCt<*[���8��A*G�#Q��[���X�xKmkb�Ph��	f>G�Fz�V���5�z��Rn0l[�U]S��!%d�>&�Li��!�9�|LiJXkȧc�����ЅcV�ڡ�cS)|_3�Jz�B(8<>��"d������K/Ǣg�N�}����.WJB(�i�Y�Q9%�ˊ�t�}q�r�!,u�ceB�DA�s�Q�����R�i�x�&g�� ��G7��45��
U��H%�և�؂჈�Q��9�%�ʊ6�[6O����9�c2�
��
�u%V�7�ĜK�1��^4���u�M��:�	�����(#�i����V����Y�q�ʔA�I�g mӠ�g]+����qJ�֋)1� 
_-�a/�*(h��r>c|p�����G���ĮVǹ��I���샱�w"�o9C]U�uپ^!��;��.�u�z�J���X��qf#H
;E=�fƾ��u�d[�)aY�J�(N������y�_��Y�ᓔ�O�{ed�T�=��ʵ���wRh-u$���1<Lf|    IDAT�������hې�}���<��b+�V����JѵeM�̭	�B��'꾤%pNPUu ��k<��d����~��?$ٸt�<0�sD,��d<9!���l���H!�����◒��0xL�7]9��iuM/M�"M"<N&�c�<�$�0��/C��
�t��� �8i�܃�NR�,%�S�d"!���g��׷��������+��1��#�f��/?��׾���Oz�`��#���d���������n�^�j~Ł���O�m-��+x�O����z���L�j�ͧ4q�X�ܩ�Ǔ'x�ɢh�X�������jba���*>|�+MI���|�[o�պ�����szz�;������bY�w�n����;,?�ܸq!������������Cf��R'�L�������'�c�{�=��f�d�����Zé��w�}�����|�gx�/�ѽ��ctԃ%�3xtv���)-�b�Q|hg'4�X�]�t��TDQ��]��,��=�s���y4���/�?�Okk����TDJ�4Ͳ�px�4!��=!?9��J��qq�g-��ɔyY�x�n�:�T���On�=���[N
��ָ���]��
eUgq�ķ�>hj�	t��VqD��ڃ=xc�qL�@�A�8r�d)��������=vC�;��r�x=�aP�ufӂ���Z�
�����%d1�-j����TBR$��Ӕ�6T�����
���ؖq �
Oi-������[��l�%��D�f�!"c�x��SZ�0֍��k�,ySЏ%#��F�M;��cd��e�
fiM�� ��f-#E�qpW�TG�	F
�$.����'-z��B��X���Y;z�$�T�M�� V͛�Mr�>g�tD+^%����XF�v���H/ׯkײ1����H�Z�O�<]�_=�$���8����lA�QG���!�Dk�O��e�'-B�n�ס
�
��� ~�Z�w-��{�[A���7�b��=ӂ��
;t�?FYYj穑�:�Y�Y�q'����X��Ћ�x��K�� h�@U��֥�(�8��
"���zK"<���4j��n�����p�
��M��89=�9(kk��TU�l2a>�����k�D�p>�������)��ZlY��� g���Tx^i��G�qD�$	I�`	�|�$�RT� U�Jjx3�3s%�l�����;l<s���]�7�"�����]6|C�w�����W��ٯ�&GMAUhdܐ��������_YKq<f�4���%��1�ܲZ�gs�O;ى�����f��E<��42bQ,�\;Ǖk����r��HШDQZh�í c���.�]�;BG��_��< 
[��x:a��d�T�eB��f�UU1����^�x<孷~��[I���'c��>��?����[o/�,� �B�ьR�&��Ŭb<Y����g�oqq�'��N��e7o)
�r�T�F���P]��1�������)���Jy<]�g	��c_3���1��.ax�Y6n�μ��k��bDU��V�ߕҁa�����#p���i��IAT͉7%6p��2�\�u��k���uT�$��՛���W�19����Yv#�P�LPU�I���;�sE'�z=T� �ֆnQ2A$h����|���հ(*W��?��^�A��V6PIO���-�>�d��t��}��D� �H�Q�*/��R�3b�/+@H���q���?��M���>�g���K/��։=b�H-C7ǘ �޹3&x���2��*�A0[�Lfs���"���(E8IE�\�R޻�>^��g���a(#���c�,�-���]xx���L�G`,����fcK��&9:�x婪���1ˋ�!С�&�����Y������p�������r/������K����P*�P;��0Jmp�B��Y����g?V��S�V����e�} ��SR�|P��Ե�SU��;C�}wB����,��+V�l{W�w��g���#��0C���!��2��Ɍޅ��:���[�	U�0EE�JzW_B���G�������!{�C�dc�?���^P��GXI���,�S"�Pm{�8A��ŕϽNk�ƕ\Qpr<�(
�Ŝ�(���M�˂�x�E���:;;�y�||��ݏy���LO�Y[t���Z���I7�'��g�s���&�Z����i@Eq����E��qR���͵k�1���{�'ǘ�x�ͷQ. ��Zcc�&���O?bMI���7�ϿF�>W��ٟK���S����)qJ�)�e�\Vm��vd�Z{���W�cms�%j�]I��2K�stw�N���3��N*��GEk�'$BaǢ�IB��wg3����ڙB���\�qHw��n'��i��y�V^�%�]�ݡ�m����J��X��ziU��:��b� IB��:_y�/��ކ�����}��x��[|��m��{���y����FDe��j�?��k	�	l�����"P$��\����]�`��?a~�I�p�r�����?�&��ptr��������Ṹ��7s�6���AIY��(PT�m���ʗ<�}����@ˌX�1Fe�BS
Ci+�Y�6դ�M�����(<=�b���w�_�38���Lõ:{`��0����`4$��u$q��$ؖ&:A�b ���(A��5�}�7��.�����}���/���ŠZ�&Q4��)
���e�/�$	Ëp���M�pH���8�	I�����4��jj�$b�j��C����7o�}�̖q���o����9��mj4��H��S#����S� �T���g1/8><d����i����ᕦJ���|��|�����N(�֙F����Ӝ��鋈#[��4Ja*C�!��zC��L����K!���'�"$ΰ��H�k4��z�20�:�B���2�+�-�X��S�R �o9��xڷcdw�?*S!�o�	][���P��U��Q�0��t�q�WZ�]��;��z�p�L�����ٜ]�<Uqw��n6.��4~�yn�/Z2^���f��ھ�����=�7����{2Z��Ni(|�Mm�������}7_D���L�xYD�lJo�֯_��5�|���)B�]��I2�Dihu7u�v!aqu�� @�t�֮���u4�!B�&k(5����:C�>��GB���8o99:���ch��h����1��3�t��s��eq��"�%�p'���dQUTB��o��a��`L�Ϲs�C���� '7!����v.�D�3lU�Ӕ��))� �}�dȸ,�8�]Z���/�dc��~�D��+LQ���a�Mݩ���R�J��Y�i���>��8����pto�_��qF��\0o,�)�ޓ�Ȥ�E�x�T�"VU���S��O�:-y�������M�t+#���Bh�UUE��O}�.Y������2��-��t�v]�aZ��Έ���� M��,K����?��g~��;�1���bN�ؕ�"t��C	��3�2"�3�2���$��k�q�[����y�����Ӄ17��y�O���k��U��g��R���j��{�k��и���������T�RKI%<^i$ANus}�iY@ hU^ �-*|S�Ċ�6�M�oj�2�49��H��w�M�(k��z������12�8[��C�%�A�P�c,�"/��!�~����"M�%�a��l� EG c�.�Έ"�H���>��d�>��� {=\]1��br�j�#b�P,ʊ�l�����}f�����MN��,�C{ERU�霩��p���Φ�����<|�W(a[д�.4{�8}��{	FB?�a[���,⠛b�����<�^$�>��y��D���b�HQ�Ф����o<˽8�l��~�9����������d�d��-�}�9J߰��!��Ƀ]�{�l�Q�܊���(�8T�@�^	H4h�Њt}�`�������-Zv�mϤ�.�J��,d<���Њ�y� ��[l�lAhEP���(]�u߯�v�u��Ë;��j��� �?#�.L+�f'5�|����Dj�hgh$�uM:�n�;���\��L�ѻ��x�����g���Yv ܙmi�v񎦱\�7{[����G:�aS�|B$��5d�EU���CT��*"�l�
�Z��{��x����'$&N��%1�Jpb�#dL���?f��9Ν�F:���&�S67�E�8�i��>��1����XL��N&��9e�`�K���B&i*��!Q�\�پ�iYr�(���5yY��lG\��"s���#�N8||��b�M��1�|�4`q�&҆��F�$��`kff�,��[Y�G=��~�7	_;�A�ޣ:=�� �j��<�)��T�Чj�7���g�P���V�@�-,��܋78���98�,�o��
��}�σ''�����7e��l߷۔ݵ;љ.�m�f�;�C��4��$��/˲�>��!DplEp�������nĲ+н�1�^��x<&˲e�j�c�A�����=�!�d���o����]����Ǥ6�0�Q�nZb[�ujk�OI�6)�)$u�p:ͩU�/����ǌ��_|��W�MflQ��	�������p�k�:b"��h�����GC��.\�ĹKW�'�y�#��ޡܺ���"��>{{�8�{���]����c��57T^8�E�F�Q�����e[Gl�ŉ�.rR��e���: <U0�{}�j}�$�����i�-��&OȒ���o|��ܿ�}*��MCTCR;z:&���$Ɯ��w���_������D9���4��W5��ќ�H�h��,L͢��g%�t��K��O�8�,%�Q��ل���5٠���R��&�g�����H��?K@����BI|��X��,c^F�z2@����t�nJ	^z�uv^�<��YK$>�3�opp*Y�/s���P��c���ο��~�_r��>޽C�4;WoP��<:=���d"#	(��Rzd$1ґۚ��(S�xlm(gf�2�kE��@�=��]�o�93z�ƛ���=��H-�-\C��J(�3o[lC��r�-�8���2Л�A���҇@ȶ��g��*�P{PI��A���!lVD�0X��ܙv�o+��sx�|޻�w8'Zk����~i.H�_\xY�C뫼ҡ�TŖ��n��^��1��A�@i>��O�{��\�z��ׯ����`�z:%Q�����;X��L�1���Q��[z�2"�:MKCa
t\q����א����V�ސ�\����-��\�֘,����o�ҭ��v����Y��oA� �R��&�/szzʼ�Bb�!%��LJ�����d�}�D�:\Ԇ�U����M��0�/�&)�7��}����S�R�����oo���	e>CkA�m�3$��Ո���Y`�D�E�*4�7<HL#ͽ�K��o����>9���l'��RP��-)��9[:�C�FK��#�4AS�C�"�W�z������N��(Pqry�x��_�$�č[���҄/�k�<���;��dQ�]�taT
I#Q[�!�����UW��_���x֒ �n�&	�s���ϖ���pA��]B���t��e�{��.��A�jj��x*��ʱ�a��E���_��?�C�1����;w9��Q���dI�o�[ Y�#�ȡl�IT,4�$6R��{��}��֗9�Q_�Ʌ�@�'8�@|��?���U�}�s\~�s<��G���Fe��.[���op��͵���[TD��G8�37���M�EE�-��!�͈�������|̓�w�ܿ���}FR����%J8�pD�$I¢ȩMC�Ҁ�{tz�|^�H��^���/r���x�x�����,`l��}�z��Ҧ����Z�,f�>�My�.z�(�)E�g��#F2/j�lDE�h�����fB��P)f�6�/m������9�T��D3�`}}��\O�����{@�(�݌/��8瘎O1E�ɣ=�3dI�8kO�����۔�'`mA:0q
�3d�J���9Gv�2/��4�#f'��}��lG���JXo������5��ןe��ќ�풙�}�?���нsp�
O��[/]����I5?���6˸z�*�4���K�yMl��Ƈn���U�`�&���1đ �
W��((<�:��kq>A �;g:��\���C�����}���H��xf=^u�X�@o�1R%xQ"P����eɿZ�V���ګU�J����|_t�|8���}B������EK��gc��+�Ϫ��W-�)�x�=�@��m�(���/%R���?�2������a�i��"*�x2+h�&J2��8���X�XkEYW�)O�@{�M����imp�CX�"&�\|�&��=�mm0�5����Q�{��hf5��Q�5�h�~�n����y{��W�_�y��K�0"�c�	nM��4%�� :T��hĠ���� ;/����,7oG	G�'����{�T�B�J�U�C#��FԵa���ߤg�����%���_��)�ia�m����z��������,rUT�|�J����#�J������ݔۗo���=>dNʕ�_��������G�?~¸.���4DB���b���)x�ַ򻬎!V�ere}v���b���J��s��zZ���k����n����9��\㨋�Ǐ��p�c�v�!c�_��q��Z�T��U8��yCH�=^5�z)"�T�SI���o�~�H~�u^��94=���)+����n>�:�[�㋜��?|�}�&�П�wl�p���(��K0eAv���L9>�1�҆[�!u�3x0���]����}B�ܳ\��"$?�d��@1��=�s�ݞ������8�<��<�?�Fr��s�x�e�/]`:>ac�Qn�y^���8�]�a�}�7G�=f���'�XIH��#�AI�
�֊���"I�}~���)�u������x�[����������,0�0�ϩ˂�阫�;�����d�_����$I���.��~�x�K�,�$ƚ}����"l0��˜���o<���h����a��J�C�H�dI��c�VC+�ҁ��f���L��)�� U�/���7�D?*h&xp�k^�ڗ����o�&��CO����d�8�\���Am��DhF�J�]q�O�A�������B�):~ƣ*>�I�]'���(��M;V��Q�Bi��g�g�g]W�%��Ӂ���OH��r`��z��~��>��|+γz�u~p�Rз�E����`��0��bI�;{/Ձ]V�\)y*q7�r��/1g}��W��
bVh��$��^D��j�
���H�d��W6���E�8��4��M�*��$I2RS�z�n,�X����ѣ>���ڐ&�H���l����>Y�Q���)^�J@�(��4� �+Kʲ����$'$M�P��hO�wk��4����к===%ъg�^ekg��sȲlI�R2�M�T�v6�6�X�U~���K���l��y��_�l�z�f�^;ǯ���y���>aF����|�_������'�[l^��ܵ�B�%�2Q�p)O�%����0^�(�(Ix��r����y�P45�_qt|��'O�I���t���)	-v`y]��<������r]~�����2	�~9����p66����;-h�+
|w@�Cl��?��������pt�|��>�:_���xQ��kb�����/���Jy�ƤY?�]�����G���{<�l�W_"{������=���9�R%RK�W�����B5�,��i���=v����[/��=���b�`����	IU\�v���+��˷�?�s��96�]�>���{��"�qH���c,�֚��"M��3����s���x���x�)Z�\�|���y���4�6�B�`rJ��(�
��A(� 	*��3�(��ϙO�$2b��>��J�_Hd#x�{������{�P	����b��)�%M�i�g.4�����8==���akzҵJF�����Y��"j��=����sE�8s�g�>��4xoy����!w�}�\��Ō�,�\[gm��_��c�Px�C>���    IDATP1�f��HQ�|���ٹq�k�|�j�2�u��e<�կ�}p�˿�-�����G�~/+�`C��
T�[�*hx!��B��R��r���'�OG;yX��ҁ�W��?u�a���w�ݝ�����N0��ﱜ���ç��jumY���+U��˙eWi���:��3j�o��ُ.�y��S����34�<���Eh�ϵ�}�k?kn�B�,�=����̫	���~��S�e���'�5�74�2oj�8��Y��Q���%MbT���N���*��� +{��u�kk��Om�8|jӠup��OBPo� m�4�E�X�\�i۸V{�W�ֿ]x^b��M�ꪢh�<g�a/�x�q ���?5��lpdr���-��4��mm�H)K�#n����{�f��-�p);���^c���{�=n�)�k�{�s윿�}�fUi;lf[�K�g-����*YO�n#z�Q4G,�akm���1��Yߺ�W��:�?���%���f3t��F����D-�s�K���W+��d���
��� >@������/�m>��˽��X�V�����mr�mh[%PR�[��鷹�����>Z*z�b�w�)�FH��m�J�6�PU���"{C��q���������y}J��+̕།��������2ɨ�[������ۨ����L ��.��~���8�ҋ�x���׆��c-·�����\�y�����ѿGF������)��,��	n���,��k�{Ȳ, �F8H���j�6�I��(��P�9;Ww�r�"�ل�tJ����9��b�h�IG��ۚ�Ԧa:����DJ`�WX�H�}jӰ-+b������?���?��� k
�d*�+�H�kO�T�$���ܹT��z�����46Ŗ)�N�"�8���\�*멬c^8>��w�=�q�s[�/ao�l�u�y�f��ݝ���e5�l������,*�$���K���c�VTdDf=QAP����XFXVcɖ|%]�����W7�z�k��Օk)n\�sw��^s�1����$I2�kW�N�ǣ0o�g�E���#�Cn�����9�;���L}�G���r���]��ۈ�&�W���_�>}u�%Ʌ�\{�H�r�z_����x��H�%?ŵq)�Z�#/���8b�ϭ���8�"��cA	��ò��r����we����->�A��
<���<=[`�CX�V[�������c1>p���ъ���X�=��䳺9�np��)�ǟU6ѝp^v���F ��;#p�s�~ޣ�l��h,C�J�8F��Ɣ��A�`�ሬ'����qLK�+
1b3�p��)%q�"�@�45��G4�!��RX�^�e\�y�cGGGHe]QW��=٪1�jb>��k+V+8E�I�2���֜���ЪZ�`��Vt$�~׵E����.�a��4S6A�ɒ`�aJI'_Ct�x�w~�[������y�����p����W>ƍ��!�׼�W���ɯ�)����Qᮕg����只�W�I�\x�v�u�b6>��K��H�$q�Z&�1���q�+S���$崘Vy#[2�B�1�M��W-��Ž�tv[l�359h��Akq�R���{���,�je���L�T�-6�v�Qr	g.�]�ch�Q�ư-�2��X�ٻ�6����8#ڸ�����Z-Ћ:��|@c�XS�(�dK��(�s�w�u�6iz�Ym��x��<�q��)�o����{�ݾ����݌�BN|���_z����y�h�o��7#>�O�'1����6�4� Cc�4 ����1��#�1W�\'R�x
�o�W��D+���{�y�a�E��q��n߹�|2e:�䱠������L�UU2B��;�ʡ�����a�3��qi����0�9q��s����^c��mTQ����~�����=ύ�W�E/L�XO1�RNf̧AQJ�����$�8"%���.�L-HK|������ӢjUP��S�&83����~�*��-�7��������ݷ��__�!��IW �W�'���|")���k�~�:4���~�c����ظ�,�'�����߼̅�ߡ:z�����p]up҄8���DYڀ�SU����4������zz~V��������=��}L�U�����I�����}(ϟ
��� ����g�Y:��^�T���p����[���nI�;�}xS�s����W �E��l^_�j)ֻ'Їż~���@Z<oi��n�e=A*�j$���#4L��� g-6��H��#r��R#�[1�Lp�����XS�IE*=��[ϑ~SяD�����=�'Ǥ�g�V��F�$�ڀ�8g0�&�F���{��M��ČX|5"\+��L���$qK�JӠ}�|�Vx"fݥ���՗��� ��pg��	�o�BS�q�Cz�&��e�����&�~��?v��?�:�ќ�ل�|Dck�i2CK�m������Յw�shӜ�{�,�����bo��k�NA�L�f��fF��26�>�PUزZ��'*��A��_Mb�_@«��T
θ���E��k\$�lPcl�)1�i+�3��"�^�.��g���N9�<����������9�[Aˡ8a#�Ȳ!�:�VRI�����hD�E��6���^�z+��4k6/n��7^�������Y�t��^�1����[�����Ɍ��S�cd��XNw3��˔I��;ֲ�{?}���~@��ܾ��n� K;�M�l6a��#�|�M�ׯqtp�������{c��5�b6"^��Z�wz��c�dYΨ-��	J��K]�r6e2Q�%���&K&̋����R`kA?�$B`�
W74Uh��y����(Xg2F�`M����e�qݸ�x\�FB��{������Yo@�$�I�d2a6+���FK��!Qx�`��K��0���|D?K��4"�y�^
l�PWk�xZ0�k�u���dFYΘ�s� �=W�\��������M�����n���YV$UMBD�R�)�`����iH͌ٿ~��B�*��v�ؗ��J��|>��?�w2�x���`�=_G	Q,i���*�J'�XG��P5M���$?�������+�E�^����<d�3�} �+��{��o��hQ��O��
��U�������xRa��8�B�,�Y���LPdqb�!E � �'�~�Moyۖ�b: X����X��*�?��p@)d�Z�g_{d)����i��A��H��ł�ݔX
�$��(��0��!�$:K�\��	�	��x:�9���/�� �"�>�R�%�ٌ�j�t:D*�J�3���g��u]�Ҩ��P�g���uSA�TkI�D4�n]�i2��KW&�2�W
>TE���ˤ#H�:��$�b::"S�^��"��/�2�����A�5�U6�]����wx@)���D�FIO탳�D�����|�;|�&�U�U�9�(NjE�t�׎y$Ȯ^At�D�ьZ9�j�>�W�"��.��\A
D�E���WoV��'��k7�+����童��ς���r�����@#y�s�4����錍��+&4�#�(��di��P�mhR`0�� �"�(���jt����3<a:+�G�s>x4�4%��!��#�O<��;�p�������'�� }�����2-UɃ��r�n��k���XY��qA�*f���̽�鵎��鈦�H���1�iA��D68C^�x���[H�[~F5�q��6���l���X__'"�����ho���c<x@�X�(Fk8>:m���p6p+��Q��뚐�;O�$�1�VN6 v���}N���&$Qޣ������XRzC	VB9�9i�wH�~�O�4����t�bG1�NB{'�i��:F� v���c�ݰ�!	5��%����+B ��4u�p:��(�<�V1Ͱ�<@צ���+�<~<��׆��}�����sz8�����1�0d�9�����+_�m�z�X=�#^����7�>x���.�)�"H�Xoi��M��5Qۧ�&�)D�o�u�g��*w����]�!L�%�Ok^�()Ck���vΡ��b3Y��<cpK���������Kx=\�v�#��yZr�����^�p�z�ߗ�y�:Vu�/b��Gۦ
��Hdx#��7-��w��`���PA�S)4�������8dG��֧��IK=���E�8F�/"�8#�L�
�l\�$��j�r�X
d�!K;zkˊ��*�4���0�����8g����
!Œ<*߅a��
�w��,���A`���Z�eEQ�4y��d�1�<T�n�A��xWUx�ё��&��Svw���3�3�����2��3�����O�S>��_���ӽ����GDN��!�s+B@+D�_�|����W��y��h	Vh��"�v�O�������q�{�}����=��)���Ԝ	�<M�y�/��'`�E@^���Id�B;�L�E����~�Z<�i�gq�3Z�<��.����3*7"N���@�a֠��Ne&�����΂:�d���"���v"|]0+J�|�<N~N��N�q��'�~�^��wH6���a{����p[����C��$��!��b��M6_�$n���d�\8���9Y3�xx�h2���P9�m(��C�՘��7(j����6���ϐ�1�dƟ�ٟ�����~��x��w���~�/��o����QU	�+��#��U�x6G��H�^��dƤ�H"E���u"��G�$��L)�C��4��G�$x�U�u-Cu9o�:T�x��):���{8�#�{����yO�3 V1�+��4���	�q����Dy Ӗ�5i���L#�& ]�ې90ΡZ�1�8\e����
���,av2��p̝;w��1ãcb�k}�(�����xF��8g'����f���(镂8N�6w0ij��x���&g�<t���fVp���+Flݹ���YB��4&$�M���qΜ�N����J�?�<MY��},{�+�ku�Q���r�+�w�%��%��_YV�pO��چɦ�P��.��;».�Rjh!х�N���O�Ow-4,�i��hZ��`-�{ჷ���}�Bx�=�P�/�o�儍y�I�ZN"Bڶ
X���â�L������n�!:�~/}�
G] �����PGJ<7�e i
qTR�"��f���O�ωT����TA:�8�Ɇs���?�3u�X��$1���>Qa]�|2iq�2�4��{��l�d:A�NF"��j��38[��z�S�`����Ea�C�����ե�)a<�T�X�9Hc�t����k��`\�4���~�/�}���y�������&������l�X:�����$a��L\� ���V㼠�6D�s�I���"(*��� �9<���FR¤BuR�tUʤ�Y�q��7����w��Y��]���@��9�L�5u3��B�ɺ�1k<cY%
U;0�ZA�D�UEACb%���ƌf�Dc�%�cb��`=�0��fadIj�H���k�nƤ��eT�̥8i���j�)6�N@|I�=Ro�V5�VC��5f�2�z�sc1&�.J<%R��Gb�g���5�@�$��K(f��ԑ����uCS[d!�Aق5�����h�ᠮH�.׳��	�bF�3�;����sqv��(��a\�l����[ě�<���M������&�������v���TUEY��֐T�(�2lP�K�8��~��>�⧨��p��g��O|�y���^���%F����߂Y�BДe��4F����He�7	�K�G�����*�i�2��4'S��LEC�A�j\�q�
��hQR�v1Z���dJ������O�����̊�r� �%�ِ4YH���51 M2F~�kD ޵{�u�"{ 8kq
�	mY/Hb�@T�?9�(+.\�`�B�$�A@I+�7$��(�)�!I�뒵<g��m"7g]A�OP�a���D،f���9��	�74v�H�Lb�-a]tq��8������E+E=�����Ѹ�L�$&��V������<���A�@*��J�6H�T�V��F�[�<N�b7&�aqm��/��PjbJ����"�AF)�*@�K(s�-+���Y�p��������t�ھ�#\� Z�!�f�o!�%�B������c�7�Jx8�--��'��G����;ψB �BX��vW���i�F�"�+Ic�.C�.*�hS��	�q��u鶴�8���G&	'�[iʥ�Ϣ�{hQzOB�zg�,�g� �zrrĽ{�8�Q%��%4y��jHK7��Z�@��&�S[�u5�L�u��P�51r9C����6�=�<qd���{�1T�W9ts\Ull_a��}��;����?��\�elЧ���p<��ʷ������?�PL�fc6�M0G��r�@o���ԧ�����>�^�\�H�us\��M���I|JZZ��'�y��?s�=��c"�b�K�.]d4RNf���t6EGq��jPļ1v��.qR��:��0)J\���#cEa*BP��8��qB!�Ή�.�M�#-��ݐ�&I��,�2.k���N�a6�s��e&�o+"Q��cr,r:G�"K��L�'��$�����	��k�r�*],��� ��0�$IЍģ�Ts�'3杘��dY
Y�� UF�G��3����ݜw~�]����S��C��p��}r�o_���̚��h:i�(�z����T5���O��I������kW��/�R�f�ol #�w��9<>��>�ljPAut:�1X_�����h�h<�i<�>�"�[̊���y���	Y���3M�d5�i1��5L���1qq-��gi�����`|TǔX$�e9����QM�v
Ӫ1.���V�iJ]m���1���Hb�M��%�ښi�4 ߮QOCYW�ʂy�<B
�sԍiG�$q�`]�6��!5ND���C�y�n4����C��E�)�1����L�����x��y�MT=��� o���*P&Q�,>X�j�Uv%�'\�qgqpu�Ї?�L~2>�����d�m�����X���kG!��)B�{�%�~�9ƷB#,���p���X8�<�'xr.7�Ǔl�6̷�Y���Pއk��)�&�����u�]�}&������{2(,��L�=S��������Tٌ�w�7��>�pDQΰUEGH�1��*�h2eR4�G
��X�W�n���ú�)�y���X%l��I�>����z=�,C�*�vy�t��ѷI��0��i�Q�lt;\������	D�#�����HR[A]�E�t^��*�-z#l
BIDݠ�0O��}	����Eتfv:�Ae��R&U��x�����潝ׂ����.P�\�f��Ox�����c6���;?a3�p�0�J*R�����xHx��Z�W�1joi��+��Ԧ	�5Vh��w8b'Cg)W/��w#N�?$q��.����o���}��w�Ҍ�������g��98ݣ8>ft�\�*�����&'e���+|���j����샇H�f���8i���h�Go���T�D�z9�I9ј
kn�z�KWo�{����]F�{�Y�t{�/|�78������0:��Mt}�Ƣk���L�4�+�i�)j�����>�/np�p�Y�@h�ܜ���iIi+�<E����2̄��c��>qe�;]�/^d�a:i�����\}�<��_�׉�5�KۨT3+�4�&�?��:j��U��w�[���J�E1^{�ց,�""!���������:Y�RU%�{���/q��M~��Ox�����{4�0Mpx������_����?���9o��3^z�_B�e����rIZ�Z��9
����i�x2��%=���19>f63hl�w���.���@ck��N8�
���GH��K�w�d��!��@�5!�Ǳ�Yɼ�Q�t��HF͛�"��=v��/�YQ�x/"��[,ec��#�1Y�rR����D&��;'p�bm(��7i�G֋��4�s<EE]��#��j�͔�ŌA���#��υ_�*7_�����K_������b�V�$�QBP����g�`�ɐY    IDATy��)BPv���K'��ں(e?Z������fO+I��o�t�0����WY�E��� ��jo;��W?�\�"V_����� �'�����'9���b�p	��6�A���g_���W5�=gH��9.Lo�}��քˌK�8A8|&)WE��N+�A�����&�防,>�8M�ZGa(E��DI�:��B�\C��AJMfDY�k7ﰶ���������fvcC?�ʍ-����b��E���qzt�����#J���ÂC����y:��J�ӒyY"�^7�)C�X���:=�e4�Q��`0 ,����f�ڔ�$� ���5"�X�0�<ż&�
gj�ܐǚzR2�xm�GG���=��]��o`�ǫ�Q2EXl֟Ϩ?��2s��~�k�d��y2!1�!�)H#*%����|�+>��pwDå����{Lw�q\�ڗy��B0����o2�?������?�����ɐW^�g��2��'d�����lݺ�����k��ʫt|᳟���N�d���!��.l���_��H-x��AO�=x�K��y�4?/�	N��:�k��;|���������>{��`8�7�7����̬�����������˷o3��:��Gd������We+.Lt"��Z������}J�=	���l��k�����|�k��+c}�Fg�O��A�`>�yO5���}���M��}FUæ�3ҤK�R�"Im�l�K\dKe$Y��`kk�n��p8����p�Ԋ^'��Rt���s�Xs��%^}�u���#�QS�e]�PH����A'�S��4�=�?��rz2���(�	{��A>ϐ:$@J�IYU�u
ΗAz�B�0���l`�/R�f1�JS0�M�F��v�b,8y�'������,I��ӥ�A@��7�:'R�i��@�J�
�@�WZx���xEP@��
���lhM��BOB�lp�K�,��Q:B�	*IёFi�L5&Jȯ���W�+��)�TD1�ӄ��,�()�]�"Y��r��w)?���M9�-���@*�.$�m��˶�ݪ:.{�"����-�S��'��2>�r��G�R��u������Xk�mt|���be��-���Ӳ%��<d�$�H� ؉V�WĊ
�_fyjy#,��a�Rg������V'HI:g�7�9�Q/R��[eҷ���Z<�������_�{�����t~�w��ȷ郀Ѩd<}���y�N����8(�!b�H�,x�ԁ�([�K�9!J4�ٔDK^��g���MP�ئ��U�q��^ଧ�*|���)�NJ��\��b������A'@�Jd��d��V]�d�s�u�^�ù�������hX�� �b��xa��&02��I2X��X�d��˒����3�cvd̍/|��������������p%�Ƽ�?�_������������_�w&�Sd�I��L]#d�
%�2~��[Emg����D;v'�hG#����i��	#Ar�&W��o]'�-÷�޷��t��Z�ǣ��Ï��%��NY�sRc���������x6g罷�{��`�b>�ݟ�ɻ����蛆���r�?�9?��OP��PL����S߾F1�Q{�l:a~z�h�!ۛ=FGCNO������;�X��F�	�k�u�sF;�Y�t�B�u{\��d��ؼt���|��ь���q}k������v�AD`!�d��c�Ǉ��E�?S^����J��Y��2�U5�;��.���O|:G�P�55i,�e���h��Y:Y��`���X�K�i��t����:�m,W�ֹ�}�+�����I�$������!���E�t����@,��������;�i��z�ݽ�@��:H9Bˈ��C|�Hy�8���-I�ι�{<��z��n�}�'DZR��7�ASZ)A���q@�i�[���H�$���'
�e}P����:Ut��M��8Ak��} �1TՄ8�p��Ҹ��O֒�-�ϳ1셔�s���8�E�-��$d����L����BA�wTKdUaM*�l1H)q�;��m���9��^$� 1�'�czL�����c����S���d���HӔ��1ƅi'�[�|��]����":?!F%]���q�oO�?��0�$��]z�Jo�c�A[���.g�R�b�Ћ�� ��:�ً��������旿�-�p�XlqX�C��-�]D�@;�Y���	�o-e3�!�^�
[R�<O��^������O[�;@��Cz�������I�i,˚�6�ź�f�׭iۗ3�F(�!��O�!�47o]g��6�8���HQ�F�+$�zʺa8������c��!n4�99����y��y�p<r�R��\BPVQXP##qR�v�"~c��448&�`�p��]���#jk�4�`o:<=����g��I�%�"�X����Q�F�s�ӟ���l]{���<���N�Q{���^���˷��y�HF���c���G; �^S���V=�m���w{�^p/����R���(�o��;"��!���M�o�Kvy�T%tֺ��a�oP�'Y2/��?�����?O)6ӈ��c����
S��V]��(�o��Uv�S�pm�#ʂ�4a��}�����h"͝�=����Ç��/��!�6�sz�f�ۥ��H�b^�o^ANO��1��姯�ʑ3ܽ���لr6B65��:G�a|z�����g��D��C!�Wq9�`8$jR�(�p���cSЌ�Dq�*�l��	UQ8oH�jkqRQ�Ox����s��:S��ҟ�F��N��D�o�/�_��?&_�c�E�P�q�b*���l]���z�z^�u�
�����92pgYU�����<õ[7���孷ޢ��D���DR1��/����2N����ܹu�+�.��^x�,�y�x��a�F�x��@Ɉ,��usz�^�6o���a\ʹc�M��x��a4��0~k]4H�(����b�,#�c�8&V^)��ԭ@X�� ;�o�gIKR�ަ��N�.���7A/CG�ZG�͇Ϗ?{��"\�
�uMS/}:��кQJ�Ě,3�X���X�XSl[��H��B�PޑV_z�#�����f�gos�wo�IKÈK��e:�ܤR��@9���B��`N�D`֟����^����Xa�Z��)��j�X��͊v�Y��d�i{�Xr��H�ǹ@�xC/Crz�����lW��rg�܇����� �s}}Z�\;B C���`�[>,t8��ϯ�ɶS �b>�`��z�O��T���ZѾ�j�·Ν�x��w#3�Bā�В7�C!�وDX`UP)��r6����|�v%[���h�6�أL���ɔyQ0�L�'c�����S����<<b��!�x�7�x"�jy]�P�$Bjڱ{J$*��z=�N��	dg�ƭ�lnlb��(]�������`:s����t�L
E1�0��!�	�J�>��F�Wh�|�9�=s������7����c�}����)w�O��<��D�������껯a��Z�xA���8/���GT�އ1�����wX+� �<%iK�{d3��������D%+��`n*R�I+C���.%]�f�T��<l�u��+�s��'��^�q8��G�r��-�?�d� ��(8-<���<��K'�g����%���-
�1��F{ŕ+W�r�r�1|�.�[����{�GLf�?�܋$�bc���o��ostz�7��;q��?�����N(�C�|��ko���	Jg�6A1RI⤃B0�eX�ί��Z�8�B"Lh�Ԯ!�$҄�ix����c��e���8�TUMGF��ϼ�%�[�w��v�!��;��/x�]D��r��-6��)�MiIR	H�
	ݼ�p8��a���l�B��w�ec�2Y֡��t����)o��U>��}�R\�t���S�vvQJ��v��89bMIw��e��7�7ll��kʹ	
��C$0��D�
X��H���^Ij���-#��A�/��jH#E�g��ֈӈ+�/���I��xo)����NN�"L�"�!ip�XG�ч[d��T(�8�W��Z�KE��l]��t������hL]�qR�e)�,02��[Cvl�P���Z35�x�ݿ'.�w��oy�ګЙ��;�e7�˕_�5>v�*����"���eY�TfI�S^�{�"F���������_��}.����d�޾[�Wci������o�R�/Z��^���?>=�-z�*\O�罷qV1?��_8z� d|x�M�d��>:!����g�^,�����8�!�	��+?��%�	��/�z1P,��U�_�Th�F޷*Fm�7\�t��t�AE�$���	��Z���E���u�j^RMG�R0�����;��%�9�8e<:����x���q�A� ZӸ����'�MYKb�d�('�A-$�����B@Z�_��@���q�x�]��F=�U�I���>��8NpR�]z]�3�U���6es���q]R��4e���c�O)DE?�3zݜf���[/��/�e5���gs6���ɔw���_��?��/�n�3?��K�R���K���K�G 5��ɶ���_�9��FX,��N�&9ESc��n�G�Ԥ�F�F����n֓jOmas��d4����̌!J�a�h|J�e0*+jW�uB):q��e�$��`i�[�<���ŝ�êF[C'�L�Zg��p����m�M�/_�2�X4�+�[��Ir�RuIk�������6�)����7��1u&I�WWx�Џ4q'BH^��$a�ux-�w�j~���G:'�<��KT��EЍR��~ i�n��ڵ-���xg�3��5��:~s�Bϲ�*WЈ�5�a�&'c6ok�<��/�$�,ToJ�U������	uYᜣ��2X�39>�������� �v����p�!����_���}��p����?xĴ�18�V����1�5E���3���DF� �P���$y��e8��"��8�X�-!��uMYT��s��_;�r�b]�:���}�67x�S����=r���d8���{\�z��4�q�����C��.ei����R���Qu�S$$q�TxϠ���ŋ\�~��~�zgʚz>c>nh�@�(��ABYkM����kE���o��^����X��w�D�aT��.�sìz����9�ے�ӍJ'�eCY׸Ɔ��)$���ʦ�g$9%�-(�S�����DP�[�G�R�ZX�/��I���;�q!�S_s��ڧ��w)ĘhQ�Me!N�ib7��y8jZᕂ��o��[V��f	_�Yx�{`
B�,�B��A��혝]n�
%"j���	�k^��@�S�# |�W.�ʅ;�w�J>���ZO$C��hP�M�Ռ
I���ɉ�`M�H�Q��w+�e�"<s�01e�K�
bs�i�7���w��A9�h���Y|A�ykZ�-����U�#�p�F�Z�amh�ԍ�J��#���Fa�7�(Q������1[f��W>OOy���lL���n�10%������G{�J�sME�2Qk�8�'̊#��|)倆*3D��Q�t*��>�E�є�����R(��$��0�'$F���l|�'�A�!�"�ʒ��6w�}�aQ0{秘��j�n�9��"�.>�L�[�2��5t$�����d)�����tdM��N�Q�TJ\7P:����է��ȣn^�����#6bn�\�WΘr���S̏�f�V$��t���R���(�y����%K];��w���$�Q��4G��hNy�IlMY��)Ӄ�̇c̅u�$���w�1L�1:� \��k��WX��6���bP+$%/[R#+���Xop��xEn$����߽�s_�
ϼ�YW�pZ��mv�!?�ýW�䗿�En����o���>ɘ�zC�ݍh�l#�ڍ�k�f�C(�1-�|����1�P�&$J����������v3��X��%[6��t:�VB��rD=�yú��L�Z��k@Ť�.�>s��{0�N�.�hN+zk��4��M5����f\X���0J����V%2r�DU�x�H��N���KRƲ��,�h�ڥ��N���ŭ[7H:9�9�q����T'�Mح�S�ǀ;ƛ	J���d;�Q�0ƙjE"5�k�KG�H��cTW􁍵ֲ.�l��W/q����HΧ����h�w�c�Jht��6$T$1Ra�+k�͌:�tO*�f�ދ�"]�fm�ar��<x�.����2��e>�����r�WN�xD���UBmTK�8a���h��P^ Z¢}lE@��jj�l9X� �Hv�8��İ"'�-�Z�� �2Z-�-��@���
�[�P$����|(a0*	\ν�����4W��O#�����p���V��PG����gF�#%���'����g-$�J�!x�y�U�?'K��؏�y�!��)&�R�	�xgt�b���U\�2,Z�i���8{�ɲ���s��Œke���lvSM6M��DQ��F�@�_l��"
0�7���� c�`[$����	Q#����a7����=c����pndfU7i�HDVTDdč{�o�.2�UC[�8���C(���<�*�m�RIs��M �!��px�;�F	A�|��-18T�tmHf��!JB��g��h�p�y��s���{�g�8�[�R�{�LZ�JQ�E�ֶ׷ϓُk�h���f������r� -�p,��]�˯~���ʽ��6�S�⡵t"b���䙧 ӔM�Y��B`��Nn �p��x�:}|�d�Qo-(�f�(�6�`{c�����Ss�Z>%x�y'ƈ��@*��4�c��锕�y�G<z�M����ۣ�a)���.:�&6��>Ǉ�ƯPJbT��dJ�k��M����6���טh��h�ɽ}���ݹ�W>�y�w�����3�Q"ZO��X�[|0,G���dd2�_�X[]K�J��q��X�Z ��a�iM���$ѻ��זP�!�B*��X��Ny����O|���)��ښ��K�W��W��}��<�ɗ��(�:�b�ߡ�O0t�UM]�x��ʠ��lT��,\�4)$�dP�de���	��}��ns�8e4S/W������t���4Y,KE={��0HG��HFnal�z��&���[tmM5�(v7i�<|$��j6�6��SFf���,w��0��p!���h
iP��o;�stV G���&eQ�R!����(�y��g�{慄;0
;�2麓/":�r��y~��Ⱦ�=����?>!,JS����E�*�$�e
2m0yN,3(3ΜA`���a�z�ܞЊ��dN��#N=L� e�Ѵ5R�2��la�F�8y��Z�a����W-��"UE}s�O����_���s����9����v�l�p����ԧYNr�\�8�st�κ;��.�'����z��p������?gu�*_�W�����ֿG?�N���˓�~��m��/���@�[��q	�u�!��:���J�Q��3^�K��@wn��EZD"
|��5]A$ ��R�O�����mr����Hx��O�1}��\ 6�HHu��T�4�L .}~qNi�YAn{F���Qs}�&������t�vUS�]��7�dYA㓤���O���,��mm~�Sp-����(�e��cE���cc�
���5�|�ζ䃜n�4�G�鄍��%��L�y��k{;EE��t͊�Zn��v\���k{F:C��b��Ǟ���{��>�ك��]O�ߍ���_��/}ڎ�7ߦ>>%� �I׺���^�\L�&�B.�$v���w���1���R��u*3(�Q1`۔�ERź�H@�ȏ��x��4�ӷ��+�Qh�s-�I�	�Lj�����B���>|��kr�(�9;r��;���Z*����fT"�݃���W�?x���ş"e`����������QB���uqr@�7�#oV�*Sk�\W���{h"D�6n;�'�(�D���原D�Ͽ�R������#�G���/r�Oq��������7�/�³_�/��W	F�(	�c~�7����;��|=��i4&���5z6'����ENbt��`]�rvt���!g�Gd}ϧn\�l��Ç�x��6�＃YP_��    IDAT�*�_5�~�Ggf�X�L%��#JA/s5�d;7�޺�ͫ{D�x���Y��P�v��R�z�!��)�������_��^��f��g�z������eL�5�He��D@^��`�����= fuG�i��VH"�Ct-G�����wɭ%,��}�~�:��Ry��Fr]��Ǩ<#� �@�D��Z"uN09Ս=@�]�eAČC1;ǁ�U�@2�(��h� G���ʐ�<Ԏ����>���*�x��׾������E�<�'�x�o��K_�֗�*����o�C=��/��."�h���S�1��1���t���s��sz�Gş���C""O�/b�G{crl����וO|�\��/��'����x��5��|�MD�dh#�� �8��Z���O� ��cn�"|�	��lH}��Ǔ��(p���E�0\�+?�
�v�z�s�������=��t�ଠ��\ �=�>�+<����bD��k��C�x�R"�]C��p��m{����ı�]אI����S��Ɵqz�>�(��m^���d��/Qw��L�ѓ�("M��:���cr'� )@ֿL����h��)��*/�����'k;���Tx�Q��I���o�M��o��ۿ�˿�+<���| �[=N�`R ���������a���P�!F�� .l�'��?4'
���P>��p1�H�J��չ�0Il��1��
��Qנ;~��5���C)ä�X)��ǟ�pCWHk�F������G����5��@gɍ'_���s6ێ��Ѯ�("��s��гٷ���~�o�O�>��vE�ϖ#�2��9Fb6Gd�lwFW�@����p�q�X&Бs �V���L%	ϵ��ڛ"x?8�u�?<����Mlے��%��)��$�ܢ�����gW*��?%/|�K�q�����=~�����9���d*�2�j���4t�w����&����r͢^��?������3�A8��L�4ǧ�ݿ���Lۚж�۔@XO�u�c�M���H4yH�e1��ߵ����?�{�mT^н�6�K��$���G�8{�]N��i���ﾈ���ߡ;�'���:0�+L0v*S#Dp}���)��}�==�oP���yJ����R|D:�[���������.��G�ݒ�{򲠩�Xv�m\Lj�A�*X	�
��9�傅�~I??F���Snl�O&�c��j��)��\A�6�񴀾%����('9!���U��,��4rmr����'����L�=��f��,����>���m&Ͽʕ�=�8~���=�>���p�������CR )����!�]gJ�K�����}�z��F�]��A>u�ŇD�\_����Ÿno_�� ^��?�T��,~0�C�C�4h_<R���rkQa��־IٕLٿdm���B��)�KAZ�T�?ǟ<�������]NxR?�D%�c�/$~׏�B$żH�h_:���
��d�B���y!P�z۠��T3.�]�::>���v��2�d������9DL���h�P9B8%hE`e;�q��h��Q�<9v���dt��@���u�@��l�����:g�FA�Y�t���4������̌	��|�d��lu�O���M<���'^��+�GĂI1%3��w<��w����}�ED�!�f*��@��ć�a���A=,Rb�A��0RPH���
!�u�z4� �Ԯ$yb>1e��I��k:��hcP�C�5&t��&1`��"�ئ!��9�����d'L�@���mZr���k�;�<Cf96B��s=A@�5�mX��0�eN�:�f	]��:�3��d�"�o��Dk���'��"z�h4v�'$bHd/U!���ǐ�q=�K�W�p.nD�1՘�dd&�N2M��|�Z6��S���?���������XAd��j8b�d$�G�;�r�����Yu-Z)��$]�µZ
��n��,3rm�j����A�@G��[�T(���~��:]+��b\tg�<�����>%�Om>�26<|�5L.����C�r�	���NJ*!	��x:\���+�B�������� ��(��������w���_��O}�1eq2'oz�b���z����]��;,o����JXt�&�Z�a	h�q�Z%e?!1F��,=�]�����C|�2�v������LʓHAg=�x¡J�A��"ט�q���CKP(F��"Nx�qI�8��ߧ{�>�L4y�d�
�*��@��� ��E��uu
�C9�:Lc�����Cփ'!���D�XS�׉����#�v��5RL���N��]
�5:8��,u.=�r{�2�u@�DE
1�c���n"�N�c�$E$YZ�s�K�>���`����\:9i�'�*�� "ka�8(%CX��������u񹆳��s��ɧ]��	qYg�Ck��>&B�;A4
��h~�]��S��[ϲu�:~�K#>X�zE�X!�b<!�%�Z���$J��v=�b�v�b��n{�f�r�+�I��$����'��]��Wn=K[$�������G�2hS �'v#��X0�$Eቢù+�U��JzH|i)���{������-�1�Sch�#�������d�bWG�V"�E���TdԷ\��h������,h��@���]QZ�R"�h�8��{�A)�L�c��ɾU�D�@�Q����?��Kɲ�Q�4��Q��B�^�2`��ipD"W8�*�|GO I�IפΗ�()�C�X�4�ـj� ��� G���<}�h)PHb�ڣt����B�D�B0-�D�:42͛�P�D�>�/�IP��+dJ�<�2=��.�/���ؐ��Ħ%W�����'���KE�`vx��j�?x�U�@iX�m��0��l}�%&g�j��KoF�E�:�"d%M�$e�Pdt��pNq�:�c:�:4B� �z��d��(G�I��,]MD^Z�"�I�+i	�=.��=-8����e�BQ��4��lEC��Py՘f���aNf���Ŷf٘�)�	j�Cv�G��J(���q�ݷ�����C�~E5�y�?��c���^ac����z�����5���I&��ؼ �� "+�b�-�1��*FMO��+���8���2��d�P�g�[�2���P�o���Ţ���E��is�G��3�<��Oqg�M��c²�W�PIp����]F����
�/Ų��'ʶHĐ�K]�p>c�)�\w�/`�ѭ_�����p��-<�G���'.�1x�����=�����3Z��/��b�n.��/������D���b�M1�	&/(�JA�y��W/�]�o��M�.�!8b�1�=$ܻD"��^]zO�ӝ~֢k��ŉX�|ئ���/|��C�!��X�������c
��@�1ȮֶG�r��d;�����K��1/�FWp�%D����IT�2G��)\�� s�%zK'$������ۖ\�MKa�#_E��n��=��2z"�޹�
�Ԇ<+1EN��QdFQd���Q�fւz���'���P��c(L���`l#Z�5�lo��������W1�M����32���Z�	������sZ>���$�u���>t �]��kC
���S�*I@]�I�X%?� Y����G��HЃ]l���%�D�#L�'��x/@e��"et.,e5����:��������;���w	<�iE��H��6��U�%�L�w��F�ƈ�h�qJ��q.Q1 P�A�ࢢ��El�\��>�K���Fbr
!������!��r�㯲s�y�ʜ��S�;W���s��|��~��/�;��^�}��Rh���*_��xx�6�޻�����c6�v1��x��p<?÷=J$�!��k�����@�+�U�s=&F�j����)Rkl�.x��&7�#66���%�k�"�9.�EF��lE���&�Y�M����8�P�neY������Bj�� 6�"66麖f6����L��(QK�)�������m�FYu��{�NГ1��m�?�ؚ���q�!�h�VW�eյ��f��
#]� g�]���G�с�)�\fٕ]��m<�&l�\���!\����,K���A���}R������2�����Ӛ�%(5����#(&��xg�����<��Q���vd��ݺ�̑M2�$)�T-�3B��tRA����(À�\����;Lp��1k��k^�A��x9�Tg������� �Ɔ[��}�&(�GgOާ��0�^��E=�6�&�\����3�Wn"���|D�	�a�B��������>��#���]���#Ȉ
�F8)�J_�Ϟ����I�e`��5�S�s�].�\��=J�h�c�a��%,�Zx��d
1�&��{�ƪD^�F�s�|�é�:#�D-�H�@v=�FFFH��D��1��E�#���4MoɄD�M�w��SV]��F�e��2�%�(���C;�P���
b�8zt��m"Iٯ�GdF���W�L��D����S\�L�ڀ�{b�������}���:�
Ĵ�|�e�EOӁ���[\�̋�~��dA��3������{��=�֠��I�R�J�,�z<1V�O�.�ԉ��[���Ja�����D_g�dI���L��I���'4qu]�L(t�pxbJJ*S��%���֢����%��N�R� �G����)���2��R��	���Z�)�!U�@�-Ӫ`%#*Z\�@�D`yvJe"&�IV$6A�JP
�Q�l�Ud�h�H�tށ�ĵt�ci}]>�SZ��o�9@�I����۷�>��/�*~T�|�5�`�y��*n|�kl�W�m���?����\�ԧ�u���p������'G�F%��F��Y6<#|�U�|���USspz���n��Η�9Z[s�8&�~qƩ���tdJS�'�7���g?C��$t-�pL�};��aS��"gu�@
��n]Ag
*����6� Qj�b�
�vlW#\5b���G�:�a��e �̰J�o��/�]��"ֶeF״�:�`������͛���5�Q�Hh�5�Gf~�bF3[�sM�k�_bf'���k���'.Z�0�׹��ϱ���p�T#�֑وo�n�x'�Dd�96�ф��)F#�e�F��C*
�]�mP�C���J��r��[<x�v����o�w4���K��&�6���C�n<���6w��{���ߒW�>~}&��0B�<��n�:h�+�������*[���햏�����@�E1}��g���.��ABtĐ�4���c�{`�L.�-�w�r2��$Aj�w��^�4W�z���#f�����|Mh��O�h�(KDQww�|��[D�P~�Bp��?�=|}x�̵8)�At�UX'p}��"�|D*�fFq-r�>1j��F�n��5(0F�� � O�M�d�X��L	�r�A���4���f5��ӧf�D���d^1ζ8n3�~᫼�o�[��0���c)`k�l��@�HV7�lG78�eEZ��`��{�2H���˚�np�MA���?�1��~�`�*q}�jl���<�k���L:��5O&ϙTc�4	��$�a��f6 �י�W\/�9�~R���Ɍ`kZ�=����9��ߤ���Ͽʗ��K9_��ſ�������+���ɷ7Ț������O~���w�3ݻ���c�lOir��j���p�����y	���#�1B'ڧ�=�af'.Z�1F��=ZhD\�\���(���Y���3�LS�,.sH���� F)D�J�Z��wD��OGR�\���FK�	D��W��y��R*B��8�r� F���%*HbP��-k��G�|�BK�,��Q}K5�2����1�S��nW�H��85�U��LT
�K�j�O��G�P�2�w(a�Ra���p���w�������L7hC$�3�_���oxtg�=�����g�g�Wh�V3�B#7�,W+��S�AVT.���E�����[�8�8U
��m{�M 6���������8?�佟��{��P�X��s|�d�|rb���n��H��Z�mK)V�f��3)��fm�`F
U/������a��~��ܜ��]d�{��%�ј؏(��u+�ﰲcak�[{d��"���m11�j��NF�Ō��{8-بv�t/�
r����?�<��'��G����B��l899c~|�.JF�{�DleE�1I	�(��آ���8��;��!�e�&-jF�当'{;�ÿ���!�w��W>æ�N�'zA�-�fxD�޻|�/������J�g���akr�P��}Q*0����C�߲"���"��� �мL�E���=6�\$���0Q18�(���1X�\'���B��0: �(ː�Cr)���a��<�'�z�[�y�� 2O�������H�{v�V�a
�愽O��/�ȉ�X���[os8�QPd%=Ѷ��$���bkw�W���1aT�LL��S�2)*^��K��5�o����ȦL��&ϰ�Ya�>UmB�{���ϡ�'>����;O�vL�v��rr�Ok[r����C�AP/��G�<9:7��|�+��(
BZr����}�)�]�`�l�-��h3 K�eJE�6e�>�M��G[�s��� =ݨ�L�p�:�|�dk�c���o�5Z)v�\�����2��-!�Ҍ���kP�#:G'=�����ą�'�
c����FT9;��.X6�{�/}�w��7(�b���_|�lY㿳�g?�/��o�h͝7~����ܽ��+�0��g���{�G��'�
$AE���ϳ��O��ĵp9+�yY���P��Li�Z�C�u�p�ne�"Z+r���@#�d�@c1��@�q��(�u҉	��L�Yr��DBL�����^�t��׸'v��� Mߑˤv�q�jJ)79�/��u��FI��ۭ	&���u���5& I��n�P��qm�?�/�#?�q"�`4��&�F���h�q��[�w�*����]���d�ʷ̏g��mrg䣂��n�Dd1o	Α�{�}r.��'e�6�4m��_.��O��!��>�XI
��h����{{r�yk���,�m�4
!#�Pt�eٶl��`�B��b2��ƈ�Ye�l�U�U�"SHͪ[Q�%yא�<�R�6$a��5'����������a$��DY��mKY�3ژr�[|�,�}�&��e�RD���t-E5�mhړb��⤓��t�,/��cm�����[����h��S�ؐ6)c�m��*�	hC1��EU%m
mp�[��1k٘v2��s�w��f~t@���0Z���w��_��믑�;�S��t�G���d9,�1h�*�f���wP�b��3ٚ@��Dh��2�Ds�L@Ui�* ZkTn�lH��(<�g!	YR��Q)�D������>�':�睆p� H	���K�
�)�'�VZ7.��}�z�W�h�)'4M�c�[������Y�����=�j���_��K����o�;��������8<<���{���{Į��愫;�d�np��iʂ헿���s�q�����l�A!��Fp��Y�P�3��u�<zp��w�����ՖQ5fgg���c|tI��h��cO��;C�&�M���F
���q�<���r� �zt��I��E�Tt�݊��4��_�9G[7�}O�%�+V��zѢL��D""=��SV�S�L�s������,�kX�S�]�T�2x��h!�cjv]���bT1�)Fy��h���紽eZ%9��{�"���y�6�,u���kרON�̧�-)�^�������޻���?��po��hk����o���~�?�~��ho?��I9�A'�q��]r��,w|�P磟͒cD	^�'�<�H]���O�N�q/�;b]�g2���H	-|H�RBL��rx_������s�1�zL�J
r%�$ka����(�$۹���$I;�aR�� �G$蜅��˖���%��~A��MG	��8�h7�����{n � � r��4����T�!�N!��=H0wA�)#��qc��Q���O��O~�Df�¢�BGIk]��1w��fU#�q�ko�    IDATM߅Hヮ��}�e��%NG���u��]d4�e;�B�a��|�u��G�� 86i<��}�"׆��Y-W��1I��p���Sh��섾��4D�|�Q-^vT�g��U�999"��j9;a��3�cw2��)hۖ�k�F#�Ɉ��ш�d�~��-gH�#�e�Z��e4���-���G�����r���U0�
/C����w��k�ELƪ��<S���)�GR7Ghtf�Z��!�Jr]��2P�'�le�E�V߰qt�t�'<�����3�w�9����gT�l�ӂq�1*�x1g:��>��ǧh&�+7�����`׫���v`!�ď�X�ѡ�G②'��R+b#�8zAkd&�A�$x��v�������f���2I5[w���Zh������}XK�^2)x���⏆m0�e�r&�|���/�c���+����_y�?��;�|���������O���[o�Mx�m~�iKAq��[Wyn��Zp��?2�_'�v���n0)Ɇvڅ]���s�/�����Ʒ.��+�pα�-!v�����a9�QێL�BAg)2���ad0(��$����c:���+"
��9p�/���?������6u�	:��AKr)�c�J$19]��z�¶]-�H�$]ki�D	��aZ��q�T��EIVUD��������	ڐiq	{�T���%QK��F��5i4B���֚L'��-ҵt�%��O�����/}�Ljhz��Y��	��yݡt�t�C$*
��W\����������_b{c��N�<B�L&�H�5��5;�96#�5j<^Ŭ�+x��F��p�:hI��)����3]o����6=�F��4�s"8p6���b� <��L-|�N`=r)��XˀVIxFĀ�~P���󙢐�X$��2���m�s�F�R(��EϚ"*�F����1��
�w�cA�[ƹH��P���%����w������:Q$@��~2D�!t	$꩔	|�u�r"�Ƃ(�MESMx��_���������/Z����miږ"7
ں��x�h���wt�R`脣��՜���y�ۆ��;�µȘ�,��پu�2��nl�)$�Պ���xB�-��S&���=�09!2�Q��9����ΰ����X�՘�(�2bF�xzʝ�>��}���i�s�����x��<}s&�~fɲ�|t5�L0�0_.��f4��[��Q�a���Z|��='�N�ҫ"c����=�ôΰT�QI�ŋ���1�VH����(Rgpm��H�F	."uҧ��WJI�3	��阢�0E���Zl������8d%�����Wg�Ң��X�QW�ޑ��9*��U�bRe�E�Rg<���JJ��)��}!Y���"߽F��K>��g#��
���Lگ��9���f����h�T�*�m�<}�D(��Vq�.�[�G	�'�R��t��M�k�v�/
΃������ɫ\^���*U�M��W����������1��W��/�.ʍ���1���yp�����|�[_5[킝j§���A+��?�nV(�)��ń"B�:��/^��3^Δ���x�q(l���C��d��w��Dٱ���h2��`���W#J	]ۢ��]�(]:�)���jT��"��4*�����$Q�rJ���|����P��(5v����>µ5����`X�Vt��
����i��%�Yt1�9���Z�E��ְ�YL^�	ɼwآ`z�*�Wv�x���m0&Od�|H�{�n���{�AWsU\+X�? �"���[̛�B)��H/�nn��=�O�y�S����M��}��1�SD��^!�b�
��(�a�`kA�Q�.��?��sq����kG�Z�!$�����@@�@&�LB3	r� ���l�T �����c�����5NK��綧RD�(�ԆB����!5��a!�@�QB"e��P"${�(�2QV�^Lpْo(J��%���mL ��K|lM]^g	�:P_Eb��Q"}Έ�G�ŹA��8!�R���Vh1a�i�[/�����Q7� cO,��u���\\�t�E�HU�]��mR�$�m��)K�w���w���9[�ȴ�pt�>G�G�N��1���z�U^��_�4B2���@j�]�F׶�OJ��� ��^6x'P��xDI�,KDt�)1��'}�\ �sB��Q���Zy��6���o�_�u6�&�х��׃�%4����s��׶4�2X���MǢ�Q&c�W��	]O9"�l���=~��o�޸Mt�%�EA�y��_�"�O?�l6C���Q*}�L+:��s(����|�DWJQ]Y ��5�d2&���^���}�u�M2�E��=�gR�D��Ρd�P�q�<ǅ�����H�e�����u���W�����s/�v� �	ڌ�YN�-�1iNt�3��p|L������6��1���^RD��O纵�� �[��K{�$�o�?�{]y��=2���?~؂t V�	��~����x�v칐�� R�ܨ�����/����,�-~����w��x�?���~�O��?�Ώ~���n�b5��Wx�s���;?�'�Ɋ����Harz�by<���Y�ϺO�w�h��N�����&8�lL�޹�j9��}��f&9FY��"q��9����k;Z'�M&C�_ΰ�f4��S�[���W��ֳO�C'��gۖ�bF=[pvz���	���r���=��n~Jx���н�(�@���68Q¢�Co�Y�V{��l�
Wn�d��g����ƈ�yY���԰�(D��z�&ǟ|����}�O���8�4m��� �ݡ�?H<��ib��v��ՂO5yQ�ԫ������>�_uc������r[F)@&yg���װD���=>�._+k:ˇ�Kirf�ph��r��f�D��x6
:��	���:�%#���L5���H����]I��+I2^�8��.'������\�vRr�NL.�U#�L �F�#��+eƶ)@X���q�#� �$x}/�?2yzlL"#k����Q� )*�T�K�&K:��'�X��b������%�̓5�����Y����ҷ�鞽I��ABB�X(���C��cl�JR��rb��3���];T9v�r�Rv ��Hb�2H���H0�h4KOO/�}�w}�����ޞ�� 8]��������>�9��;��w�P�VΓ*H�KFR��55�� )δ���@L�Y���jPƀs�vEj<�H0!!S28�bw�`�2�,m0��o��l�X��lv�rc+R��y���iʍ!G�����%kgQB�B|
]��J����x@m<y���}'�W��������O��w|�sW�����9r�6�R�I�������>y����Z.���<�9BېHG�b[l(�kQ�R�%�ŋ�����A���e.ln3$�\�I=�i���Ȑq��@���u�$ӑ�+<2��JW��#�l�h��V����'�����ԝa���e���1�̐*�u�Olr�	��2��7�b�d8N��Ү*.�l�ki�{����?����e�E���_��K��+����ⲟ��n�+��O���������3w_�޽���W�޸E}��hk$�2�4�'��\=� �x��>%����:������<�	��	ޅx�?Yx�͋�������2�_g��ϳ�縻p��Kw�������H�?;>�}�S��_�����?{�ज़s�_���{�a��,^l1����E>�<r���࠳4��x��V��=������r�>v�o�&����#�<r'�� NYc�҃�R�hE���{�E�L�������7(�=J������@�O��'�6Z��6����]��~χ(68��q��ٻy�VB���C�SԚ�&M�tQ��9l�'[�<�0�褢��d�l�h�i��k;�siF�et�Y�>�s<]QqL��IЊ�Y1�ڡ�������V��jΓ�z�H��a0r���k/~�G�{�g���p��[��)Y�x=��.Dz�q�=���X����Y�˷�n֟�J}0���amnq��$�@�I,����K����P:!#�]��!���rq*k�@p��Ѕ O��#���<��P��s�t(!��;��E�)ВP$��b�U�RD_JC�xL"�2�tg��z=�8�]q�9��y �-D�'w�M�<
�߿^<.J��m(�9Y*I����Χ?C��Y�W��1��f]ͪi�F��`��6ض�5��S��=�l��9�1L���]�͒���xa(G9�@kjv�|�[n����ѐ�k�C����cO2n3�Ni����ٲ�jV�m�Q�#t�Dc�����-����p�Td��^a��%�Ҍ�#=S��bUa:Kj=�ݻ���*�f����.W��!ÍM�����f3��Υ; L�S�'SV��8��p��Q�iV�����v-��.b��I-��@���s��n���pgD�D�P^�7O��h%}�W �G��D1(Jƣ�(G�G��t�D�*��.˸�m���/}1�"M 1D�l)�)c:H�I�ԭݲ�H�"�$�b�I���۰������O����O�GA����?΅x�G(�����hB�{��P������[�K/Ӽ�2��-���mP��{ʚ�����#�^/'(��Vs�����g[�:��{�n�O6������U�"`I�� Q�����l^�'�3���K�o?��{���}�S�|����?�?��oy/r��^�p�]�fwz���1E�c�d�Z�)��Mq��9����7��C�V	�[�h�M|�ca!�J�����>[�66���SVՒ<�M_��SK��vΣ���iQB����%-�*jaI�ٮm��c��w�K����gZϙ蒨��P2�t��)�}��2�t����{��@H����,�S�U7a�^��4>Q�_`�s�$�|���>G{�L��a��,K��`1[�{�>��=���+���������2H��Rh���F�,�!�^��co�s��X��f�
��3��;���/�"n� +R��x�I�B8�T:f𮧐��B�d*��LX/�^�/寥,�?�-��%21!�	!�B��MuB�C�7:y�s�VR5���y��Z�T�J^�B�Q�I�L�\�XW��v�8E�#��T���N�'�
�Jk\��$R��A�Gۣe1d~0't)5J���3�
G�8�����������/�:�A���������.�Ӕ"���#Z��)43�i���)���%^��?c�l)�	z�E}#e��5.?�B'����Ӄ��ߙ�+a-����l��f�s��+6�C�|�����sWY�B@�2��˩Nzs��L�#�>�5�0I��ߥ13T�E���[/0��f���MV��h�����%��r������ӨA��j�B`����LIT*hWG��[��?�3d{���\��3� �jͥ�W�x�!�՜�_=�i:�N)�4�c�:Ҽ����;h��̧���rt�7���sWɛ�k�,�1�-,��Ӟ����i ��=���t�ι�/��ۣ�?�k�yI�j*��\�J>����K�}V�Os̨`����aNP�U��LR�!��S��G�@Z�4��C�jq²�Z����|��������ڿ���;B�տM��E��_�������]���7��M�0u��[iG����H�^�鸾����c>X���3�3����`��8��A@�7fY��ЋP�jCR�iHq�Nq$ٓ�9��s��g?Oy�a���'�iA~=�������?�>�K����|�9�&�~�2�����-�5�l3�[ж߂�S��}�d}qDT��_�DG9���<�ݡ��k����,sjΟ?�p��:���a�a��U]������^�U�1�.iɋ@���eF�f/�lڄ���Ҕ��&/��پ�v>�Y��yQ"�g�����̎���+/��hz�r��Z-�ꊍQ�v2Av�,������u�,6x:��?d�Ҕ��}\��W�򞧟%�2��N��pT�(ͭ7��>������댇��S^�J��a�HjA'[*9���Ŕ�W���'�'�����[�!��f�^�2�?���9&W��;�_��Ĺ|�M���0�|+�֒g��eT��J�%XBk��1�5��;�$>�ŏ�GF���+*Mlp"Z���6�Y�(2I�����ѡ鄦m:����Nuԟ���[��h�Qx2�Ht���2}HMc=�W8����Z0H�7��h}�_KE4Jr'-�%��8"��t@�[XMW�&����.0?<�:�"|A�5�8��ŷ�7 j	}���:뵶�zv�t*����s���w�@�*��HH|Ԥ������(��$L&�AB��B�]z�_��ԏ?��{��>�]�G��=g��]�x�U�jE=�s��]V��jŷ~�'����)(��9�~�7x��/���S�S�5�N�!
G5�b�!�%�f�%��!�Z�)3�b��-e�s��y�T�u�m8��ݿ���v���1�}�<�}�$Ys�F�p7�#�����Q��L&Q����	�������˘ʲ�������Pd9��c"�w�l�r�*�}�w����b��٧Я� ��[�@G�H=�p����O��c���+�>�s�{?�{�P�$�S:'��ޭ�T�#|۰�ګ�n�d��1[9�?�[�^��+�bgW��J�s����`F2�������:R��X�"2�L�54 Ü�wh��J��z��~ �������A����g�$����D�Ǜ��I�u����o?��9�+����)�=(��5�l��[����s��{&� &�:������%�ka������v�o����X�u�m�0��+�~o�=�K_y���������?�q]~��?�}���;�_{�������+7xx���,�~�[*�i;\��A�V3
n���`�v�[iVg��dh�o���ի���c�AʠAh���LʒE���mDV�����!E�PI����l]z����-�v%)1�p���ml��3��)˜@���[���/���-�w��o}��b�'P�5��c�m���XD��>�^&Dt�6�F��%��߿����o���_�ȳ�<���磓^��TBp��C�w��>����?�`���r��A#?y{��%�m�hrv�x���N�IN������k\�SV�)�_~���=C>~���~w��D���"|���N{����5���8A�.���{������� M��X�`"H�����e@`1A�X��4�Et~oUwUU1�lnI�(gPx��F�� �b���c¢��f��2J������)_�Ƞ�Ҥ=�y�<�ͤ�
�U�"�d1[���^#ORu�}gq�Ğ��eQ�@ʈ�_�N���[=�@���lcH��]�z�\�|<�� ��Б RMP!,*M�s0= �)�ѐ�.1�Lp��%M�l_��N$B �c��]n��*7o�A�6��կp���߿�l���;L���H�h�꜃�K�癧�VՊ�ʰ�����M]S�%i"���e�5��F9�ul^��p� �)j��]�R�y�,����ͻ(��L+�#�T�9A�[���uv����,f3��l_|��E��`����gwx��m���O��w?�+�	�R�f�bgs��v$JE�$��r��A�b[��}�!������Xۂ��	ʓ�9�Ʉa6�GGێ����SOp��C���$E����H�χ�Խ�{-��� ��8�R�Y_�3H(Z�ͺ#<�$����Q*����������6�<�B�Αz�ߛ%��F��E�Ք�5�i��*t�F<�������9�?0|LcHH�S���/y��3����$yBgR�	2�P���k\x�[��/~���?ã���7�4v��?����������7���c6ꑇQ��C{�r�#�Vk}���	���4�&�����шF&��N�8_0�|�nj2��BiA�DE2���t�z�%k���v�=��x�Y�q�]�ծx�d°j��~_H�N0�u�b>����LI6�c��GT���C0�    IDATx�#�d��ͪE�T�"�)�;���b��;.��_�*_{�E�u�).\����fr�Ѵޓ9ן|���1u�$�#E�T_w�Z��Eg�z�����l?�m�\#N�f��o����i�헸�SRn]����	�z��_���jE��$m���C�J
R_�������F�\��\@ɞ���e�J�q��j��v��xmdڟV�i�(�_7�u�s�����k:��R�giZ677�r~�Q�hǘ��)��r��"8MD/��e��b?#���~-�SE:�W�T|�A���O�u���$C���:�S�h>#t]u�����O�b5�Pz���'Z ��'��m��=@*5�����d�P�(���@��K���h�(I�ޠ�!�m�	����ژ� 1A��!i�-g$!��1��K\4���7ys:�`Y�4[��x����������J�봲���,����w�p���,��W�9�X,8>�RY�1u�iZ�
�ڒv��K��iIV��DB�f�4ï,ͪbvp�l��C�r�_�A�C�wv�f�|����dX9?>G�T��۬fKk0(���i�,s�<c��#}lٮ� :@ſ�D)�>��R����"稪���22�w��Dg4m�J3R��%L��G3��KI��h���.�`yᕛ���|����:l�����m�On�����F��FLKB���V�\����o`/^��P?��b�������{m/i��)*C��*��}&̛��ȣ	���-l��x�'�g�q��[;�HN��g{ԑҲ�O��H���[������ן��&�>^�g����_����7��|�������?���t~���l^�����f��mR�U+��tz�h <�3<;������S���G��}o�����dE�x�����&L%��#��h%N�k�r�F��֕�l�6�W���?F�ķ��+L��h3ДN2��t E�3�ɔ��L��*��UU�uJ�S��1�� 
��p��5��]	!�� �V+�$�,K���͛�mK�Z��1-B����<��O�[�3�*�WUE���J��6C&������=�m����[��)߳��kn�|Ǎ�dp�w_�L{�2��+���U�n�s�e�
i<}��O���11�KE����}�q�H���}�:3�ꆗ�k��5MF�Z;#鐬ږ��0> TJ���:�$��KLrA3�'������h�s&��ϿSj왾��}2��k��(�'ON�JB���?��8a*����(�숀Ht��ɘ�l�g�5�q���iE�?T����I�Ɇ���sgmnp��-���t,[C�(��h�k�XemGYB-,m�^�0������ʕ�d2�6�h,�[w�s��G��S/�Qs"�QQ�Y�X.vHF��-�H�t���֐����Ӵ�����8��,�wܹs��|�	R� ��"$!���f���'�%��$�뉓*�;�hW]ס��h����y��{�_ۛbL`<s�<+W{��ܸy��r�7�"�YE����s�����f�%:-p�Fc�u��u���t�(����g~嗩����~�<Oq.p6�ޭ���;�JR��	�x��K��Z#� K���s'�����NL:��Ht�@c�$8Kb*�t�S�|Ͽ�����D�M�gGv�����|v���U�XN�C'D|o:hZ֧�u���Y�9���;-S+��	Q��,p�q�$�H�P���K�\�K/���.���?���z<��|�����s�ů=9{�G��#.��4SJw*@sv< f8}�t�9�u8�O|����e��ҭ�8gY�j����E>�\iO)2$A��� tJ��hg��
���Γ�����^�G���dw�>h�\�x�Ӌ�"&Z`L�[뱶�mEElLg�#������ $��w�i��є��mn����#I�1 U`<����Tx��W�^ess{J8�i��j:��M4���O}���1�0}�k����]����v���s��9�/�Vc�Y�'r0&��Σ�@�5d.�1���u<�mL�d��$�D�vol�`���z4��)�O~c�X���?���i�w����Ⴚ�"�>ͰZ�!]@Iؘ���Ls�jư���!��p�li��9�������2�3}��=;�W��`T� >���%J�� ���U�H'�'%|�#�ޙHK2=)!I���ⵌ[�����v��;���>�'�A�t�b�1����lmOP8��+=�	�|�NI�Q[�(4��:�LRF�	�ł_�����O��C����ڳ�{��o����7h���e�̆QV8x���n�1A%h��F�g��I�e�	�9+,���'���s�&Q)��!�r���s�I�'���,G�%�zEY��7��SL�����$t6��J�U��P���&bP�px�2*3�D���X�c�xݳZ��{vwwi���`�u�����{l�7O����h���th��9��Q�߉X]��N�j������D3��/?�s�����:��t>c�l��fg��9�jH0T͌z~�sa�<�F�.��'y�Щ�dJ@�Syez��(G�2Z-�!M���]�x��|����A����7y\����oy����gvD{��2�m[$)g�4=o��V�y0ߏ��d#8���h�@h�C	h��h6.]Dd���>�]��<��߬k�O���S�������o�2<�0��p�c����d瘶���x���A5�}�-�����ι���������0L��� o0[�X6+�J#�FhI�T$i��RѸ��^Qd
�x>������-��\e����"���B4m��$�O}��4�~��!�,�K�B㥍���Gq{�5Zk��1�t�1��(c�k�b0�4�)"�lp�9�q�c䎠,�ႃ��+I6�`0�qG>�:jiQ)��1�o�&�/�ɽ=��N�ē\���ټ����_å��,�
�J�� ��i�$CwI�"U�� *� �$I�Fuo$c{-��ҠR
�o�ޝ�KI){��F%}��:p���tuK�to�ll�)U����2(2�e�d�P� Xy�Ga�����e����肃�(#��*X*)�"`� b�am��q�Jys9��3�D}z��~Ih�������}h;��4��I%#�x�D�{]�b���N�2
X�����.lnеG�{��&�QD�����Ķ%źRa=�x�h;_��~���#�t�7n����/���G7Ⱥ���$K�vxR��� K*�� 4�(�j�#�ə�e�I��:��$�����%�W��h8����%X��dJ����R�x��Xע�����h�Ӛ�8�"����tU�r6EiA>�����{L� MKQn�m��W3v����c��f�G#�4M�t:EG[7����Ɋ�s��욮n���	ΝԙD�1Q�Rͪk�VBp�U�k�|�ݽ1i��j
C��I���J� �i�"��mY��g����a\�����s����A%F���ld�x���4����%�>�]S����o��CB��{�������m�G(g�U��a�z�����z?��ݟ��'z����N{�'e� ��к�TD���&7P���O����ώ�>���_��O?�s����K��V��w1;s";�|Ҁw�g��?� �������M��e�"�5��M�Ʉn%��Å��
Z(z%����D����h�%�$���-�UC�=�L���Rg}Y��) TU��8gI2M���'P� ��c�����{+<B��xg1�=	�k T��H�ٌ��,��'��eU%5I��l�����Z���h:g�\⍣��f-��
������x�Cd8Q4U���=�7g��K�O���i���T�v���q�ݻ�����<�Ĥ�"(��ړr���DY�������2�)E-r���g���)�TQ�C��A`��� !��S�S�,Rx�2ckT0�R���t�y��r���� ӓ9)k����^N�ºL��u�[J�<-�N��k0\�i�JD.��!��� �´]Lx� IL(�R���(|d*�)�՗�טyR	!*�<���v�	�k���d�F;�xo9��WK�4��@X6����5˻{*a��e�����Cn�|c[RJ�3�yk-i��dB6�(��z5c�\�&��`m�.���'=` �	�f�*������� 8عx���dE��?�1�ʘ[k)$Z�D���dV�X��l��	��)�㺆��@�D��9Ǉ�8��yJ2(��4�����67���ES��j��i����f1_1��Z�����!��H���mɓ�,ф^�&IR�L	ї��r��ZDlnnrX-X�IT���	�x���4 7�t��b0*)�\ehW-��u-"Mq֜�O�5�\s +:D���kH��7�p�������G�����a�?z��/|�G�+��8�Gw�6�P �á΄�X�_�-�[��6�,�ln��4`���mm�,*׈L�)7v�r��Ǟ�&����x�'��SzP�<��X,��9�x<���q�=�['g�[����g?[RQJ��`�����?@H:��;:f�u\x�Q�=l?r��C�у!��sl]�D9��\�TU�����A��|��ۑi��&IB)tR�2�ԫ
�ml�Ȩ'���,�HӨ�B��^,���h�+�yG����'I�j��=����!m��US���EI���b@�=��n[�.r���FW�<g��ɾ�}Í7_�/�P\x�ݴ�6����3?ŧ��O����'�j-|��"ae:m<eg)�#35���,I:�m@�.3WQYd퐵��9Oj��$Ρ�E�-���V5�j�M���ب�^�4�]��jC�����jq���З�C�=T��S��<�xSa��d"�ܖˊ�u�6�-�$��[E�z~�>�8�`z�"s���{�I©��)F�4�y��E?�=D9}�iq�Cz�&�`N�F�̃|`���'&I�l����k��<XD������:#02G��yt��#���5�{�$#w�T(�޽��n�_����h)1�Ś/���"����#�&-G����P�)��E�;spPZ $��(2�DE��re���M���x�|>�_�/|己�c�\ $y���D�I��(�`e:/H���t��`Jh�i꺦m�jqdYF�e$e�C�eB�u;��3��BHA�J1Ǵ�a�XFIf�'�s�mn!�[Y����	6���>��l��\�A�XV/���8L�Ȋ��hv��-ZKD��	ɢ1,���*6�/HhZ��q=um��8ƞ5^;�Wѫ$�	Y������C��<��3������= 㱕��b4z��ܡ3�"I���g������y ��R��Ξd���nUB"�gK����&m6!\�#���?���z<���x�������w�FN!4�7��)� ߟ�Ύ������-`�u� ��~������F0���?z�]��wh�KFD��e˂�����x�5�$�!{Ë���oݥv���9V�(%pb�VK|p���$8S$�T"M����tBx�rx�DJ^�֔��h�d
���Ig�z�WD�q�Zᄥ�P�)�ΰ>���}�l� �,�9�b�C�nH;���NelT�]���M�[��w�ń��}���}��g�xt�����
�����9���vX2,6�v�2��\��p�j���Tm�v��+���i[J�XoJa�d�k��kw7V%�b�^K�.�%��`�2-s���y��,-<�(h���u$���Ƅ�R#�%�^btJ����j�2�;�J�y���AP���e���K�ӷނx-���EL(����A��Z��%�:�)I&�x�B� �BJ�V8���2�W ��}�>���]����ٚ�mp�~�kc�F�_���=�u�n�o-*YbE���S�[[���H~0�iвa<�hT���36�����l�QR�yU�1�m��
�5E���D�DY�n�߬d�2ԇ{\��M���H1�GHODŊ�����K�G��(��/}�U�r��h���`Y���	���z�R=G��.����r��Wؾr![d�$1��"`�9*#�̌�L
��bKx:��v���C�����+�.�"�k�jE]E5WI`4�(��9 ��PU�"��OVdg#�(�S4�����%� ���VL&���	i�S�:ʲe\gI��%t��l�sfob�;��m���4�@.4��F8r��uY'89c�W��@����ğ�����u��}���O���������W�G5��,�B���"�n]�Z�v5��H%$&�Tk胚�gu���@����cc��kEY�ll��\�o0.\{�����g��WAI԰�����[������7O{���O3ȷ��ק�D����kY�X�1%`چP������\.�f)%��1��}^����w=��o����$f���T��@��d���0ޱs���ߧkb֜x��f�m��e�$��0G R���|eo�`��t�	:�)���R�h���6����8i 8G��Fn�o1U��>�zv�%&d:�4-�i�����on�Ե����f��9׮l����O�c>P9������}̫��
m#��ݴ��4E�N6���`��,���y�V�;�D�����Q��u5��i�=Y[�:!{bCP�A��52L$f���RS�6�;�soQ�#���Y���!4�E�؇M��G�zf@ �C���7Xﱘ��E~^��ɾ��@��׷J!5�Iȃ=���f|=����{��5p�*�G�ǖ@X7�Ϯ���:�>=��_+�0�8:<doѡ�1uk�w��7K�L>Ax���k@'��[����}�Q����v�kȵ���HS1)���2�թ���"ୣi:�%�Y��8c4�Ŋ�����(��Hr���(vo�f�x�D��9�n:.^�̹�;��%"�����4-Y�P$�z���)N	^~�k��x�#c|ב)�c�ø��X�	��tm�o��m+ eY��:Q�1��L��4m��3-�{�aA�
%#�:)(u�v1Y��V$2|���̠4m�������P��E��Kq�f��Q2;O3��%XK�%�{�lm�II��x+��㮊��'{���h�[���RH:����K�H��襟z[p�#�p�Sa��wí��ٻI�K��7[����3C�@N����pV~d�,$i^0�l���������_{�UB+� G�-κ�yk�_�w:����F���0]I�B�}����j�LS|^D�����,KIE�pX�������<c�x�NI���ֈ��T�Omۖ���X,LFLjɷ��[մ�JK�AN�j�eRJT�o<�A:,#���Y�psª��V+�,�����ܤ�3D�W��X˂y�R/Ե�Ɇ���#��<-p�$���|���!�7^����!�O>��7q~�3�)������+��ٟ�¦b~�M���&�LF�Tp.d�[^���ي��q��K�'���|�vh��Z��ȅI�`2�y��Y��?�[Vci��AGH:FY�ְ`3aj�z]�qw�T�֊������0��@�*�"aT�d:�L�����:�^�%{%#O�h�v[U���$��tB��48�琱�.�Q�����@/�=E��t� ؘ\���6�X��F�h��$0�9j28�������@P9:OɆe�v�KB�Ո4Q�f�r����v�1�W�ie�E��B�A8�d8`Y�[G�����ZB᣼���i�����>�6

��[�uE���,:�C�>ŕ�cw��j.\��PD}�Q���߀i�Ya���A��8��8�s��xU"�hum��j�0�
�<�Z-q2tU�ЮI��1�P�%�Ʉ��!���:���3|���I�"�LiR%Y\���G�&�!	�! ���V��#ӄ�k1��x~@g��˒2O)�RI;;��*�ihWK�8�o���ƶu�F�w����`5z)���Yk�JS�l�q�����pr�!�g��?{���������W_��Я�    IDATT"���Z��wd��k�L_AY��#����u7q6��u�/ �?��[��$M�����b��|e�D��@��tݢ�@Dc�տ��,N��V��$Nˌ��n�ֿ��&(�ړޕ��n�x��tԘ' �b,�YT�3_.�[c�$�H�]}��l����\{�J�;GSU̧Ǵ�a��Ҙ�ί����1�������y�T������`qB0%�O{c�g�D}�kW���3O3���a�����.�g-NH��{h2�\�����&�f�]�$��g�z-K�;�ߛV���ՙ�M5Ð��,J#�l��#��X���l�������b|!��̈� ɒ)��(�l6[���RW:i���w�sN�&G�(j
U��޻��k��y���E�LmW�o~�ce�'X�V#�R�;c���ֻ\��M����$ڀ�
#4hI
�C�����5O�T��߂O�QBcTbR����\z�
;{{߹��:f�E�qi����'J��xĖ��,�>s�6�R�-�Wu�*%�\<ϥ�2�*Y���{�vf;���v�4IV*��q�(�IqrPM��C����(2�|ȍ7$r9�.E�0�R�{�Y���j!OIP�u��"8�ڠ&p��!3iq3��h�S�4�Q]�l�)jf�a��&W��!bK�ωG����Be'4,����#x��1j<b���)41f9\�PU~�0�;���S�%B$�q���.�
��d`�d_�xBl�"�B�DU��i�#S��5ͳ�z�t�ó/<K���WK�mI��H��a������򉫗y���i�?�m"fuG�u�mK)�A����PR�w=�(�^})� TU�;�hi�s�v͹�� ,�K����R��2'	"�@��J����"!���A��s��ք��r�eY2*!���VF0���(��]d°k��h٭jjS��C�0��yd�6E>dGJ)s���3׬޾��+����Rq�[8��6���t^�N������AJi�rҷk)eN�J�#3�CEkɩ��)�V�!�pԩ<���q�gH�S��=2����O@8N��+�8����qR(�.|:�S�H�;��a�S)e�{rCzQ8�p,W-��B��[���a��E>��O��H2P�&cB��K�߹�O�')�����?��6�������,N�ٳ��s'1�[������J)yꩧ��+�e:3�NI)��p.�j{۲Z�X��,�5.8����`qĢ]Q'�vl��x�8�d�/��>���������t숝da�������!8�W��$��6�P����C��(R�������0�c'�gIi �Lp���Z�T�����q��>�j�ؔ�"�e��(�%^��`$[Z`��s���
ڤ�w=�²��晗��ʳW1"G������v�T�����3�6��E�9c>A"����d�z#Z*J	c!��B�L�TRS)��b�o<�S����j�2��O)�b�p3<��o�����f��A�$�s��u�*M�A����]���SV!)z!�a�����Wx�%JU��3�e��e�x��{��s��e�����Y�<��i@��?_�4+VM��S��� 3/�R�� R����C��]�6��d4��Z��7HB���W�\aݬXV��e�-u=)D�ш�o��#̨b���M*�آ2�����y����w(�Y7}�x-���q��L���x���>EU����._���=����7n���=�mC׮�1P���hLQה�	øj��" y��)˂�e���m>��K\�x�g�{�w\��Cp�q1������f����
��۵$�Y����-�I�\���G�����Nn�h2�D�P���1?<b����\����G{���N��tB8t9jE��%��-p����s�:���E!����SE-gn�a��G<����!��Q���ܹ�
�=�M�-�C�����:����YW�G_�t!����+�Ć4�HF���'���]c]�v��z�	��������S���SO�QO���儽�/_a���;~��HU���,��ܹ}��k9��~}f6*�I*�x���̞���+P�!���{��킸�S�F�>X���m[�ݚ�r����4��dU֮�쩆��]t�E��������̯�*���7��Ã%����N��_�����?S����g�߸�(�kTI�Q���7�M�ș�C�%�R	'���Rt�l��l91��(�p�e��Gi&E�jE�R�DA�("h�e@%IIVA0�z�EV5I�L�b:�[r<?F�@%5[�&��}D����i{�ڙ\JI��X�F�SꈌL��.�@Ҋ����Dk}� J�|����t�	�H�I~ñ�h���=��zz�����_2RS�n�R���e��	�lK�5�S��Ԩ��XU�z�P5)�<�@Uɹ��ĝs�@m*��_b<��{��{)%�[V��o�����{w�RhC��O<Ͻ�#����`ow�T��G�IR!�B(�d$Pҹ�������QՌպŔ5��3������=�#xO���;,Yk��2Y�J�I�1��h���J��XL�B��((tE�S�\�z5ͅu<*���S��x!�(��U�'_�,/��27߻΍7�ٹG׬��2W�f��3� ����HRk}�1-W\�;ǳ/��'?�J���EӰxH�j)Q��*������}|pD�tB�w?��ʭX����y�&I�tK�!�Qx��8%�*!R���S�w����o��l����l��� rvH��<^��D�*�H5�HMs�k���:��fg�qS�m��-��0��_�������O#F�1�<��ܣ�����w�gf���G<8��!H!�_n^73�}J�F	x���}��;h��&�L+C�+v�\d���ڮ
EB�	Ѣ|kQ]K��~����;�v=�7G}������E>#pC��ͰcLCX�Ô��@L�J���^�;t�e������>Ef�N��٘I9���̵�*�x4�,v��E�6k��gy���H�����q���
��aM�)����������{�S��_���PG��[� /Je����C��s�?Dbv�8�lK��Dp�Ѷ!������~��6�ʀ��^B@�DE6��B����h,M�!*Vѳ�4�1�st!)�	.�v��%��I��tm�-S�6/��P�+-)��*I���J��$Jm�ƪ�r�R&H�6�ƅ��^����>����5��l��T����B���;b�x�<ۣ+,���7��8�	��H�%Vk05Z	�]�@._�����SO�޿úk�x�"?��W�����Em���\ƶ��#���o�����G����w�x��ݛ�� �IF�d@ˁ�հ>�x�qYv��bIGĭ�W�a��y�qN{�!�syk1\�h�]Ǩ�h��#CYU��˳n�18B���a6��������Q�1�~�KvϝG̶�����X�O|���6�0�!:ۨ�^@���^���_�o����~���1��Fk���!F�d�ߜ�m�lMx�Os��S��98'E��+O��5����< �:Ѵ����(Ƴ	tkV�CM�y�/���߸Υ�P)4�|�fpi�qQ�$�"��U��ݦ�:|���;��.��'
Bd��	We�N=����=���^<Q�KD���o�x
���9���mXϏu���[���(�1��G���6�K=��G!��G�;[�6_o��f���u��6�5"C���IK��)6�!%�(�I���S)%�Z\��H��z�߼�Xo��aqD1��w���Z���Պ�耛ￏp���ۼ�X�>8�?���<F&�xaμ�S?Ƽ���e�xg�&F������moq��E�j�12��bgo�3�)5;�	!$�r6��Q�"oڮ�=�i�J��&����~己��K��4�Ǟ�{�nr�O���/��ӻ��m����	2jt�Y������8F�-.Y�����y�3&5�'n�-QE�(z�7=�:�5�ҢG��P���(��خS���g��֓�b�KvzM�J6���#h\"z��з	5*
�T�A&�N���W���]��e�(BD��A������kA��K�i�6Q�O!�Q:᝜��L��:m �3�I�,�c��@z�3�N옫�&
��tz�s綰�!HK�z�N�lb�,y`<��ra�y�>`�ko����K?�)w���`TWL�5�{�����Y�.�0��}�%�z�-�޻K�#��C�n�%�f�t�5):��֑��c��L��l�bB�w����g<�e��HJb�ʆ=U���i����lG�,B)�sL�S��{�.{]�Ӹ�'	�Rdӭ~}H�,��E%���������{|������8�dV/���޲8ڧ9>fq�w?�Flzl=�R]�)R�j�ل(%m�捓�� ��K���(�U��(����L�S���|�����r�CtE&�^I���S�ݽ��~���y���]c����kJ$�*�aE��,#�;W�>��?�|��:���(��(�{1�@��8��e��ZR�B��4��G� �@�$�����P�5���`��O����_�H�cy�/�k�,�"�jRג�.B)OBh2��I����'�μT"�� �'���ov$��S�{�R��hL���!}-<���%.�[��ɘ��<u�&�x����]����4�9��1v���L�$n}���:yj�A�	�
A��͜���z�o;�	�[#u���I�Mi�H��n����yܢ�[�;��#v�1w��w�GKo@��G�W���}�Z���N��׊}+دz�H����z�X�{4c�m�(]P3Fs��0�F�8C%s�Bni��S�Vd��)rZ� �,Y��L�ٜ�͜~���9�<%��TD��8�B�EV4�#JJ�q��_׸(h{h{��!E�?�X�ƱS��[���j�״�Y)��d�KK���R.�jcw":@���X'�� �Ȣ��X��B�f�e;:��Q8����u�	b:�0�r~H)��@�8h�!)��&���!�1�lF�2.�%�Y��,��Q�e6w	�4wԅ�����h��.����������i��Ã�s/��x���+f�mb��Gk1��E:�t|�us�����/�5݇2�-j��ܰKJUH�,�4����25e	���d���O�8���hW���1ٮ�}g������[�����*��RaXU�I5��U�Ry"ms�Ȃʲ")���[�����z�M��ѹ���)~��Ȗ�?�i^��Kh�A�e���� �"S��r����������׈ﾅ<��tVrW�M 
�����q驫e���#T]�h-��Fnm�G�f/����%v��2�
�v�%m��z���K)E��n�jG�Y����5eQ�n%&Oo3��*�H�^��RN7��;��U�b�F����!��k��X�����������GhDC[�luAɨ�{&����)K�G�)U&�
��bD:��#D��4x[?2?�B�L�w�"�ii�~Ľ7��勯���#�\;�7�����0�$�ǽN�W�L��Y������O�+���G�]fq=�Z��F�.F&!b�	�ːOZ�(����V���(��Dt�<2E���C���Ȩ����Έ�l�3zcJ.��ۆ��H�)]��&{��Q.���&�6|Je���Ώ�jXG� Mv�rC��R��Q���[�v�V������#1�q�ж��H�`�ŗ8�S_�;���H9�Ex�J�UAun?�HL۱=!��&	|9�5�T�����\�g��Id�p����L�M�(�0F����Ѓ�MR�$�6$z��}��AnȔ�S���7�ˎ6���(5^ff����J�Ͽ���(9Q"��mFz*E���Z�TVڴ}�h�q{a�����#ųS�n�0EF�-�^�ф��h`�
��gU�v#D>R|<b�����f�(�M����!�%E��0$�%hC�Кp-���dٙ%F�#v��QB�z7�,g)�����ki�9}��N�h��4�5�slᐽ����!��9���P�\�JϹsS��E{����1�R�X̉2�J޿�~f�Fx�h�kL�p�1�F/<γv=N�TB%�G�6�^���Մ��uM��NPVn�ޖ�S?�9.>��}C�%��L�Lt}�[�9�����9���-�v�u��|ݢRI%%�?�].�s�Z)��1��0N�P�h�1�j�����S��>��.]b2�h���M�������oQBP�&��R$D�F���)I��F�D͉�u�^"��xI)Q)�c �����,��鎗��+���v���*ʓ�(�jyƱ6"E�`��;a�A3��]h����D���B�@����ٹ���{י^|��D�O��"�sl�(]#�v7�a������F�Ǟ���Ʌ���f��3�dc�#m��CR�:P���J��TW��s��將Zw�(�i��u���7k�vM�)@���=޶���J���&:�^wL:˴�(#9J��*���z�:��
���E��6Kn���ж�q'r��낲�b��/Z!i�����EᛎJ�H���r�3���/���+���L˚>��z.|�%���}��(g"@H]dmvL�I�L���n`V�l�ъ���S�غ�ו9���њq�)��i)ddRVh�IS�2BJ�ݚ�%:�C""QB����+�$d�R�$�FU�BPhC
�-rRH�@�y#��5��1�M"EO�Z�
�LV��DRh��!C�d���!��k*ΐ�b�GG�j�%v�����J���_����!�����@>�Db��D�  ���L���q]���T�7-���q�E��T�g�F�t6 �DK3H�����|�b9'������tK�*Ҕ׶H�0���0m$"
��$�{�*y�����В��^��/~��zε�|�\�hZ�T��'���KL9a4Ҝ�p����.9~m�A�A�Ct4�9�:�0� �FW���K�[���u������s�+�8��5;�Iv�#�m�@��+l�7���M�姮B��:�F)�l<Fc�5#Q0���c\*�&[�7���wL6aY�VXk	Gy5?<by<'��&S�x��+Fӂ�H�=�DDԈ�s��čOʣ�s�#:d;�AĞI!i<��Ï^����o�)���=�� �l��c��^�Ǽ�Ɍ^q�l��Q�?�D2�(��0�"Ks��׸Yl����Po]���;��ꗏ�8��r<���2����!�<�1|?�����l>��OlX�b��|��2���j1x��l_����B�-�s1J�dYX$֒�[\��|O��������;bJDr�\�o��o��}�qY���â���Kl��">b�-O��D�e4Z	�utM���!B�TƠu�v����QL�3B(�KT�=F[�N���|�B���6o���PNvx�g����/�*C���,"E��r��׾����<x�5��PF���6�CuI��O��8_s�y��t�3+�d����qag�3�u>/}�O�YX�!aà��XM�������[&���t���4t���a���@���h����b���l�Z�䬃B��\��i��S��z\�Dm ���$��b�yͼ��E����E�,U+�x���r��#��|H��9�0ϥ#>A�Erm�m�������d��a-4o��;\�ݺ������v�r21ѯ[�G��5m��뗜߾�Jo����5D\L¦��$Re���#�LY!�f��.Q͒Ż�eK���>|�5�b�*h�&cjS#ܼN���΅�H�����！xp�2���FCr,D�4���u�-�[��i����׮��̳l?��h�#fWs��v��]�Ժh-&	���?u�������]D9\�7%֭��I����C�GFjD��uL�d�HR��}�b��[�2��"
O�lom����[���/o|��װ�c��Ϡ�!�D�̇@)���)QQd���=Jk����w��<�{��xH��w�#�    IDAT��c���!��� �g�C��*ns���	t� T�>�y1!bN��"�F���!�aqL{��ϼ̭�_{���r�GR�n���o�������j�먢��t���~8RJ��'C�O��/�?)�<7���g�C��)w\""��yt��a���R�T��$>)\���"�G1�����l�����{�����]l����^��$&C�[���O��Or�ӟ�u���Q@�
?huuRx����UubX��B�Pj��i��Nq)Q��JY�k��1*C��ڰ]*>z�u��`����x��a}n��AE�����w�����f�'_g�<ŸB���Qf�ܤ��O��|n�ə�#���w�AF\�x���E���H))J�w�;>;�� ���ږ�לT�G�'� -41%�%�(P-�.Q�g��8��ad����z����^S�]���� 7e5B�>�u--�F��h��6ЯIm$���	���cA�$�=�Hg�1!�D��KST�2����	E�Q�ݣ��C_��b��%�Nb"�DYWhJ
� �xG�9��R"BOX���>���'"�Ii�2�T��<���%��w�F�r��TZ��)��L��V��F�5kT��]˞�)�,����� (@׿+^�������a2�H	Z!�>��,üS��"�T�v]�D��&x @=�[d���]ү��$��B�e}p��7^㎂ŻX�V4�%��=B��AnH�Z��c�Z��&�޿���me�Ibm�ͣ����QDZrr�B0O��떬o^�^�1���m��Ǯ�l�mEQ�&��s��XOg޹���w�Ƿ)�=	Y.u���9�a3����9�D2�i�g�*9����e�x���o~�Ŝ�t	���x�
��E�(j���So�!�t6�� [q�+������(K<à?:�;�9��O=)�����~�ս�/}�����qt��/����^��ަ�s�1H�,	y�~7���I��0�_��G.8��M�Jn�R��}����=����$����"&�2٢�� d��R;?�l�C�&��f�yQ��1@�"�D�}�͘����^`��A��Ĭ�hb��j�6� ��0.+|���0��!JJ�$#�FgǬ�B�i}���P輩)#223����L�@�e�#��mn��Wx��AH�ňX�ip��0��J�P#M#�%�J���G��7B��w��t������4Rh���$._bww��G7�mK�?l&z/Xv=���DJ�!�eB`m��ђ���]�H��Y��L�����CH��g/�(��1w���Ɖ���/>�D��� �\��a�P��5��l�Z�0X6��>Qr��I�	<�:˨��������"&F���7��h��qʨΚ}��>	";����"����Ѕar�2/������
���m!�V�f3�>��k;�v0\2]d;j-]�a�CEA!MC���)QI�⊱.�M�?O%8���7 v�2)��&*��pNYh
i�%�ɨ[:ee��v�BjCR#D���-J<��=��ضa�{J�'8K�p��{�;����T����b�\�>��]��E@:G�-B&b��-��E���e��W�M�(����9R�H
-�)���#��X�"���5�C�@)"���I�W�,ǽ�n$�Ai&�FW0��j�Hx�("��e�>���Z��o)52ETTt&Q���{��������g�����M)�<����R�:�	ZA�x�Ǔ&�t���cr��h�!761�F��a!I!��cL$��4��(����[_�*/���q�����w�~�/_}�s+�����_����U�}n��iW���Ȋ�z=����Z���I���!+�����c�<���$IJ!�$GL�Ƭ�����`���1��L��Nn)!�Bh�wB���CG��1e�����dA%RDnܡT�^怔��Ϸ����ڟ~�TMKY�(FctU1�ؚL�@�n��{���TEI�s��2Y�(]����8�q�Ĕ*�,K�.y����u��I:_W���Ï�3 �HL1\0�%�"�z�����A$�P��"^��N��yL�|t1ȹNeb'P����A����M�sKb1ƙ	�����Vs�n��=MX�=��Zg������o8O�DP^@�n�����|���ۄ.}KH��vV}���L�I�{\%��(Ifi�����R�6`���#Lh��˶A��Ai0�M,۞�)3QX�����8
R�X������^��>^`���N�I菓�B&Ɲ^���ײ��		��NU�l?�	���g���@�YvvvH)�3��x���t�9v��Y�	6s�����&�	�6�����	1��6���>1�%+	�Q=u$�X��s�l0T.W��
�G�Xg�b)�����3FQ#��b�]�$����W���'�6��)#jta�,�����`w��:�b�d�#��.��ۄ���)�X��������z�;^!G#�hD5M��dK%��2�Bj���B�H��A���icr���	�G�|��HH$)�.Q��Y��:9N����N�c�#,�p����Ql��K�ʮ�J��:`��^�����_�׏����������W��{@$�11z���Ա3�{�>��^zx����c$Iy�m��24�S�B���ֺ`=_�ܼ�������~���ʿ}u=�x����_{�/���ۯ~���%�sp�.#`�9����_I�}��o����*}�������B���O��ic>���HG�#{J�"n�'���:���S$�P�P�@O FE��6��(�&��B�Q���!��J���b��(*������{t�c�LiC`>d;��)QAe4��4�$v0"idQ`L�G�)G�U�ָ�	t� 56zj����l2�ЮH

�M���rV��hJ��!+��J������P��:����N�6��3�II�q�Y�WJ�<�03-��m�)��{t�r�����sj�����N�.)tQ�Er��O�2�	�GHM�����M�޹]��RcYܠO�#]�XuEv���jVQ�@):���Ao��#^��Ȣu�U�������Z���D� �M�E�b�\#(�˒�2Z$�Yۆ����.B��^|����/R�%���s�7(�{"R�q�̣����H����Փs�4��k;�VG�;>�l�c��%�SX�a��GO��D��Ӗ��D'pn4��-](1�����&�1ED���y���?��[�d�+*�����3��Wiz�YZV��)(M�ozJY�|��vk	2B��$zg�uE�K�	;)�Mp���l/�һH:��
a*:�U@(�)k�P�w.����n��6Z@߷��s�YM]���vuL�h��_g��T�eϑ]$̦{�$q��4�,�~��7� C�!��0��s��\��UV$�@a;G�AW��P :	zo�B�9`J�Y
��4�c�{u�q=��9��ЮW�.��H�6��Ld�3r�C�i��v��V���7^��)�.~�Q�)%����{oQ=��	A'�aԗ!��#�3(��?t�+��"'���3��
 hQ$�#�v����!X��%��_���k{����߯����y�s?�C)�_��_��������/}�4�����{�d��ւ�;�*r�W���$b� ��!@`󁦔B)E8q��	u�aC�ܩ�$�I}b��;�S"J1��-BH�n4�$[ll򉖂� %�gP1�#�^�&������[` �HTT�Xd�U�
������5�����b�#R'�XJD�I"�ݚ�Ĵ�̒�!
tU�UI�Ȉx�s)�(�5Cg\	|ʤ�@���j��Dq��(\�0l֬(�O �@���O\T%�o誀��Bj���cL������D���b ���sQ�I t$DO|&� &%tH@���I��(�) X�a�Ɔ8� 
E��_�DlZ�y�;���Y"��I>GҦ�)���4r�3/?��g.�n�$�]�T�B�\�y��w�HD-����>���mM]U�՘n��s�gb�.jR��?���L8�0�B�l_ܡ��al;^���ؕ����78��C�[#d5������ɼ��]�Y����"ZiR��AJ���z�}��-�����G��+�p]��v��]՘j��Pe�4E�l����0,�1{��R#L�-�J+M�I��VqM��αՂ3#l4,Zϋr��)dt;��O_����9�D��(LI�Y�HuY��H��0eAY��tx[�𪪧6�#��\1V��Vjɹ�ĩ��s��)}�a�t�p|�lg���6���j��Q�fg4cO��c�%�H�튭^P�%�E�`~D���������2�Zz�h����~�Wy�^!h���Q����]ߒfT�h��:$oE�V��R!�@��(J����ح����17R�_r!��j��9O�Hj��hH&P,3jp0�l���������O�����h��I��?x~���`�M��yX��JlL���Y��y	$�ޓl���RD&|���I�Y�	� �ʄ��}B��Ќs,�>����6����/~�������o���7���~���Ɗ��w���o�O���������2��o�o��.���(	)K�|�]�V��=e+n
��u�o��:�?;�}��;=��0)�3��S���G�]�5�ٸ�[<S@R�䇟.�q�amP�Mo)�9�?�����Y.�d���"B!�<2w�z���~y�s�G#�QH�����)e����g��?��&jx�C_?Г�%�=��:yl|���>W���Y���Ӣ͏��ʹ"o<9�XCȡ:y�(3�r�E�}��(H>P��o��x�����m:נ:O%$�Z��/�1ۓv��]9� �
���O�$$�L��B���!�G���k��&]���o��{�~�[\c�$�ш�9yu����2>�|o���CE1�xB(��g#\oQ)�"^��;��U�!�re��b��
50⅒�����^�9:s\0��a�[D���xL��(��y�^3���x�u��_�3���w�mM�ܞ2.R�x�Q�ʊJ+��հ�.)��dݕ��5j����=EY⃅�4^#�k����v��w��{���{f�Ҥ��7�6r2�ٔu�2�H՘5��������y�-�y������,wy۬�g��8�%S�Bm�6˖���$��?AA� �#:!0p;N"ñX��I�c���/#g���{���r�鮪/TUwu�s��p������]]��W߾8���b�0���G�52_�ܹ�uC�Z_�Jw}�ю�̈�x{���8��ay���g��a�� ��ީγ87�.���ln�ke6�3[,q!�k��@gQ+X������zCC�����,<�B��2�{,��ZRZ͵��o=��_�}�G�<���?\GGz�2���֯Э�#���.���%OSt�$^��Y�zez��<z#�k������L��p	1���_N��k����_d�:������/��G��?����S��{���������_����_��=�?󧾛���I�/�F�̦��xCln`LM�M�\c����[���=��4L�=�qz��(�0��g.�����`$Ĝ�!��o!8��˥Q�͂Y@Gk�a����B�<��!66KXT�\c`��㖫��n������ֵ�̙U��s�ڙW������LR۲�����\4Cd�+��ξ�iPe�5N������;v�U���(Nc+>%a"�"ɽ�8j��XW\u0v��7hO��u�;.Q�w's���7��5�f��%��������Nc�=U�˟��o�b����T��p~����֛���+��U��6��}dJ�6�ާ�/���I�x������jźuxױhj��5;�õGHw��5Ǵ1�}�tG��� $����x��+� �*������K�G����yM5ߣn���k7���α~��Yp�->�0嚝�r�C�-��ei�m8���W����@D���l1��愝���+*�qZ��G��O�ʗ���ڀ�Hŗu�g�u�-�4��%�#�]�5�H�!`�C}���5�7�f3;3\�@��=<&\~���En���pr���7���O���N�l��N0��m�qG]74�K�����y�ut�5^�f9�T1�2�n�0AY�9��p�_��DF���J��P�YH��l����o<��_R՟������f��������gYqmձ[-8:>�Y�!���,��T@*��i6)�"�>G,�j�� �4����c���/qk��=x��/����Wx�G~���У<�ů}����폞���^z�߬��W���_����~�S���'>�_��?�];���_��^��u�-mbԥ:�)B�253�F���-��d#n;�1���9�|�0f'Ɩ���4�	��@�"ģ  }�b!��#���>W�S�D?���P�a(���8kSÛ,����T('��������!�7<w��y��3˺[Q�E칮���Ab��	.a�?�`^�p���(T��6�TN_�S���wʦ�³i��D�[ i�hj5��D�Mo�'W��>Fޠ�$�L���6l8��&�28��z�17[��.X��N�5�������GQ����gb��R�2v��q�yc�z�	���!�W��HU�i�Q�)�S�|�g�N��� �]��C������g��G��U�0�@� !��'H�Ӵ�e�Ν�x�����}�=� �9a8x�2�~��\:ڰ0�\S�l;�ٚ�7ܨf�\��~f]�����M�p�v��rC3(R�EMfhk��X����J��ڰ�Σ�.��#�|���:u�c�D���2c�X�«�^Z�:�ɚ�d΍uMwp3�onn���}f\�j���\k��J���^����x�e�IK+�1��RU�ƂG:�7��`حgԪ���f�ˈc�㼏�9�68�gO�~�tw��8*�V5�W{�(�l�\���:�=�����~��g��1�b���������[6�F	f��;r�6%s+Q8֬�����Ķ�ek�*ֱϵscN����ƒ"�������oK�6;�ivgx�|���_�շ����?Ȫ}��߸��o��'>�w�],.]����1��_��������;��/|�^�~��;���ٟ�I��n��-����.����q�#vL(�hC��0!�i��B�1ҧw��G�Ɯ&D�+��-�ަI�Wi���)&���&�J�'�\>٢%�A�$��U�j�ͺ������sƻ5�nt4����qW�]���Q�$�XJ��ޱ�@Y� �'O ��bҜ'��j���~�S@����Qj���!��B^b�!�XK���˟Q�ռ4���P�|<��PG5���i�t�[��h�x��U�_��]��]�*hvf8\PDb]��c���="�\�9fK_��'D�'k�=�O��
����\��;�%ө���6�=hXASp�sQ�&�Tc7�Lw�o���,�&(N,�mp"8�ؕ��*�X.���푃�~aB�̮��@u�#c���Џ��3?��[�vkv��x�
a����.��lf�vp��3n��r��{�a����?�ct�<����_�lZΝ��4ur�t�.Vt�k��%}l|�Ժ��i�A�85�͌�߰r���ªC���j6]|V�d4
)�$��ڠ�fwQs�>��l1#����9�Y����w��������O3{��	t��gT��O������X��T������A���c\��-UP��!���7���j�T�\�Y6걳�"��9�L"��e�Jp��x�sZ�"�Oڬ�"�g!5�y�!�2�������_�ko������?����m���G�v���?�kO�����o��]�Wp����W�;s6W��=|~8���-Ir���u����5�l�I�P��������޼��1,��C7-��U�����\��G��{y�v^���[����폾��U��1�z�o������o���>���r߽��?��̌r�my�[č�<C�    IDAT+7�n0?�����zx���ַ�Ӑ�z# jc�P�Al��,M܅�z ��̌�Z�6��߯��gg��?S�|���=��@uV��N�"<i�2�o���uX����hd��<�G/�a�(���teV[.�-yX�M���{aŲ���X��m����M��=9��݄>b��:|d>�0�m{�͕2��{�V�KM�9k�9�'��$�1R�8��N�|!�����
kj\P|�XUf�$��J����GG��[�1�5�U���W�����H4��QC�s��x�,[r��$AC�G'3D��B]UQ�433\ ��Aƴ&k�Ӯ��=����ht��sYjye��]�1S��]�oŌ#�$�R�"M�$J�r�B!�-A�5�T{\;�G~�G����p�u��	��~n\����'���C��=�)�Z����a�oن����d������Ƚw�ҋ��@N�h;�nS!p>�[O�!
C&Rv	qO*oq.��R�8�QpA	��Z�hlWl��a�;�+u�"z��y��_A{���3�O��������w|��y�{>����/j���*o��$W�����k/������ɟ�><��g_fvpL[՜��?�]|���"'{sNB�l'W���\�nW����>�%�o�9W7x�Ҟ�^3�u��G��ؚJ<���L�R�B�Bߒ�S�L�]2���9�To>ϋ��������z�_���K�w����k�����>����s_b��rmp�Ҟ�+%T���Yil�W��,t'�(5�*�?��J�[���%�~��$�&�+\F��,�b�x�<oo�Y�\�7�S���^9��+or�3������A��v�K�}w�ރ��_]`��13��~���_�ڕ+<��3�j�~�P-fX�,ｋ�Zn�z�X�[0jSQ[��1'�g���yd����˷�to�q��\����,�R���I��U;��˙HHBYa��ɦ}�S�DIm(�4�lC4�q��QLҌ"̼*ZW�Mǥ�S��1�̪�������8�e4J�Q�L=���2�[�`���cs�Դ�͂R��T�ضO0�<���Ef��汉ztO�*�H�0;�*С��`U�R��)����q�48	8���2׀�]t��@!��
h�胲����Z_0�A�c�֝���$
�#r.�*�mn���6�l꧟~wʢR�x��c#��I\� 2؜.�7Ifz��6���=T04�,I����.�|��Ǹ���'�䩓[p~�>�<�����G��S�@^ycg��;�﻾�����B5cs눯�Ư���~� ��Œ�۰�,��t0�b��$+�@l&�����y�N#�M����<>cFl,;+5<�2E|tZ6�Qvvfl��,t��M`v��<�3?���pp�%���"��%��� ����������_a������x������
Ǖ�����ٜ���K�3�fE=�,4
Tn�Os����?�/��GϿ�Nepj�lx�݂v��"TZ��
��1KL̈́~���{)�
'�����֋O�n7uy|���?�ο��^8�����o>|㛟�'���o���.��X�^��#E����es�����e�Ō���AS��39Ɗ�ʂ~��>kV%�U4�����l�Ys��?�ԭ뜰Dd�|�CX�G�s���B�	Xw����Y��u*S3�wYԻ�}Wò�����+��	��M��Y��`��XíЁ1��NzSGE�q���ؘ7�⃦�;���4�$�����1�i�ۙ��̿�Y�ҋ��~���*�4l�1=�+d�(��������^� ��S�f�*5�	O��ر�l��M�ٔ��Y�[{��EM"i�Vb��rZ۶�^��H�T.�_
O����v;��6&T�/��O3$b4}n�������U��ʫ�57c�u����-�V4f��@c*@�����;ܷ�������M�J'�]b��Zb��b�þ<t����2�<����ƺ�-c+����X��)]�@W<����h�^l����])!���J����F<J��Ēh:hmX�Q36VpP<&vy��&0�y����������+Fx�o��(7^{��ц���7n�p�{���L�8�O��/}�ç����,w�d���[S�P��j �Xk��-~EB�sŅ�l���u�Pi���&^j�r��G�
���`mEmRbkb��5T��t�������#�p�e���/�����Ks��>�?�=�����'��!��!��\z�a�}�}�u�eړ[�U3t�q����.?���`�G�:dy��؏s�w}��8D6Q*�AfP��U��:
���:Î�@�,����+E�e�Ն�A�������n����������~�+��K��=|��绎O!����o�ܸ�G���_��;����k�2�8ٟ��ќ��a��u�YE���(`e>�������0�>���m������9ʾ"��L���8IS�� Uo�F�ZΥ�t��+��Ҷ-��8�jkh��\�u���8��u�J�xU��.� ����]��1�X,�K�7#bD��f*!�UT[���x�����Yi��?;�di_M�th�Pj$1��x��opY��h��x��O�RRSh���-�A%k�a���i8gKs��������F�gJ���&���l��6�����sQN�F}��],����3n
G���1�F�ɹ�:T�lf��f�0�������G�n25��Z`�y��L!ܕ������۴�SV�,��2�TN$��6g��W�&�6��(U�N�� RWt��E�P����]2�N���a�9:���?�����M���]'ت�s�u�:iڱڈI�Wt�>���E%�)r�2b`��;,�/V��[����n�X�<�S���8;��������n��YI�,�EcI�bO{Qct����1�s`�&xG��ص��'0���q�8\��wQ_?b��K|�ſO]yv�5��s��#�w}�ø�*_��K���o���1��K48ZjnՖs)�^��>�S�ulk	���5f�QS���Y݀�
�Dw�HLÊM�t�~�T�f���"(5G͌��$4��+��g>�	�]n~�Y�|�+���c�q`��囼�~�ko��c?��8?_p����݊�n��гYV쮏y囿�l��V�=��?��{.V�����gv���tu��tq�jwL��0�
5���Ұ]�E$�c%|�qT������\��ھX��9��n�d���/�g��[�?������?�������?�=?��)�p����ˏ�����W����_�+�\��z��ۗ9\�X�̙�C]�R[wb�1�����eo Bt�ZS�s�-5s�[DԦsiS����gN4+��g�{6QN?ￏ��$�O�ڼ�ſs5��t��~�
v�xR�ۅĔ�M���<dҢ4ϩd��d�/�;k�g�����dj��ZaW�GT_СZ�y�^I�c������Шa�����»�x~���;X�b�:!����p��kgi;G���x�!�y��}�K'�F�ŕ|�h���9���]��4��ɹc��=�g�ܗ_���,��W����^�\�j�[6�Q��ž��ǭ�uYA���Fs7ոÜ�.?7����S!)=t곑K&��=z'�K?/w;�?k�2��F���_���!��e�;d����wq�\pН�g1�kg��&��T��>�?����c\�r�Ǿ�x�	������g?��?�4���u�RuZ�k�o�t�\Bp�]�cS[W4�ڝ�J�Ҫm8��nS�Y�`7�cj�/wؿuH}n�����U��u�m����j���>b�س<��G9��\?>�2v��t/�=����n�]��i���]�O}�g?�;t��\�/	��;�[/le	.��y��o��< [����c�6'kB稟��E=>��������?�;_\S}2T�?���v޼~�G �rk�ߺ�;9~�l�~������O~�.t7�㯾oS�;*_�A�Q,���V�(����Zlw���M��v�+k�@ʗ=�~"g ��=Z�u�U���r��}��&��,�5i����8Z���g�?�ۺDS
�	��m�L��ސ�@�B�X���D�TAc�D�~�}U.��G���(��3� &��^b@� �h����kϾ��z{����7������t��W1�)��1��c�S<�����Z}���?��c��L�|�yq;�L�1�����Rt�
I�Ph!��gaI�j���w��/:ش��O-������Gm+5m�q��tNA�^�3�v�!��&R��_w
/����6�J����ǲ���gb� ���Ӗg���:iSP^������,h�U3N�]��Ϲx�.��9�n�ij�[aW�RR��A���?���{8Ys�{��]�Np�w!�1�+��\���r'�	�Sk�>��235�V=jbS)<m���fͷ���І51��;;@�:�v�y׻�͍�6�t�f���"��j<��[��Y.]���|��+�egv�N�ci-]�Q���;����y�s��:��_�%���������l��i8٬b�U�mZ\�Q�Cu�o��7��4,B�A�jEc�Z����/r���q�=��λ?���Z��Ȧ��#�9Uex�2�/��Md}L�Z6+Vo^#�N�'�>�b�J��0uCf��Y[YY�@����=�t��UeM<��N����&�������kl�v3���]	�12
��*��0�q�V��T���ʜ��1��q���N4���O`;1���s��ޏ���5��z�}�*���ޟ�^Mj��؉H�z��MǋϽ��6�l�g�
���%�}��VR�)�k���<FIoOȷZ+�7Cszg<x���=q��������h����a�qZ���qk�9�\��_@l�[Ѷ����<�肀Ԑ|����9�����:R����~�;�=�,V��-�M�o�pu�;<�*R�^���`;kجZZq4��f���i6-3�\_\�qd+�Պ��}v/,y��ț_��wp����C����>>�S�Ͽ}��z�]���ê�=��:��A������֛��O�i���竩,����c��9�{�ON��;a��s!,�x�[1�k�[#'G���!T�*��.M8���.�Vp�Y�������!v܆�>�;��O���XB`u|B2��B-��/�,E[�w4��2ݤ��|<
6Ů����A���6�>K3�1?��bo�P���c�9�p����O�hW��x,�����K4�i�x�������%"ɥ��7!��n�������1��~+�?҃Оx����~�mf��f�61�@�/R�_6�T&�G{�.����	C��.nwm�b�]K٦-������Sߏ��~����M~����#���7��<�B+ۄ���a;I�l��ZW���;�x�M�I9�;�]'����T&�"�����L� �l�ʰI�jz���ꅳ~���'�܆cF8�m����߉]
���:Ì� �5��x�Ȉ�{T<�������2�,�(���N	�جM������$��*Ov	�Q��6�2^�>���ΐ�Bs�B��Ti��������3�,<�(���������fya�p���/p�R������a�ܓ_b�ݝo����s<�����`�y��?�ݏ>�+�>����9�`��3��,��,7�k��sB�8<>a��1���շ_�m�`�R�l5��
�9�*��{�=� �T���T��	���:��+�[�\I����!�7N+e��J=W����G������	��	�����_���u��n�NN�>Ԇ��i�#lZ�U��Z�h�k
Sz/�����n��G+Z�>�TR�L�uR��^����o'+և��)�%f[�Ϫ�Jb��
hE���߀�Bc+¦P0�&?v�����4c���C�g����F���D�)�G�Z�ۀ�䠝�Q��MʹASy��S�1���}B ��MV�r#s����uM5q�)!�#���Ҝ��,p�9�&�|����k!��_�� 
�'l�C�^ɀ�cg��[0y����K����J��6uC5��c�������3���s�X����C��ޤ��jf�������]Fb��Ts?�ɗ{Q�m���řȵ��A����ɵ%Y8�XN_�����9���c�|��6�ؓuX���|��MQ45\�$2X䌎m}ڮ�G|W�Ǚ�m��iky�߮PQϩ5b�LI��g<�c<oy=Q��h�G53\������g��[�p�����������������o���]<��?��������xϣ�g>���^��+�nR�[��.�W���0��去�į[���:�E���{A�v��`�7�Y��A[vfU3Cv�S��/�x��.0��.��ជ��3���q��Wq���.��朻x����!;�oۖ;���|���,�ޒ>�����g8�l�%�c�5B%U�|0�(�BSմ�bV}�.Ֆk�`~[�����&YՔxN\JH�`��t���kX�����VAL��hq�l�X�'hL�^b!7,�9�s�Ԑ,*�%2�^�˚|��K&��F�d<��{!��+ж����24����cm�}�r��i�,�����r`�9s�߮�wXSj2��( ����%�ٖ2�MЉ?��}��&u��d3k��Z|����u������O�@!�'E��1�3J�4XkY�6m������_J+���7�B��~��r�6�ߓ���tn��8K;��{�瓹:	�r@��X�9�)~a:�@�f�<�	���g����۬��]�TU��y蔡1O,b�{]�d���W����L7[ 㪶���5��6{� ��P��o�z'\�v�?�|��~��[�1�C����\��S��������h��:��#GW��7�������C��]<�������>b�9s�p|�/��'���/aև�ΝG�!�dPaٵ�F�+�X��9��
�v8}z� ���%�+K]��u͆�����56o���?µ�9���#"\z�A����޸A+;�������︈�k����2������>��G���'�����ϸ��	�obv�f��X�!��QI�$MZl��X݆q�z�y�{&8���]mV,R)���EUqA݆��kQ�upxϩE�"����ǢNjll�k*p���a$e� � ��l��ޘ�W�`�����"&Z��}U�)ˈ�{]��6:�S�q�å�}A�����jRJTD�U�oF >��ՀļޘGI�@��~�(�R�)�k�~gA�4beM?���b�Z����ٌ"���W.^�7�ȂX�ܨ�{9�-Z���=m͠X}�.�&Zk����Gd��e��s�@u	������o)����H�)�ֿ?�MO3�&��z߉1�W��'�6����ͤb�P�%��`sj�/��fM~xf��x&c�����&|�	�
����#h�p�]G%��]Ƃ���h�1��1�~2v"�Us�q���!J�&W~_^F��l��p����q�7��?3�W��5�Ն�>�\k�|��~��>���Si�;|�g?���Žz��kG���Ǚ�s�=rΟcg�����|�����o�:{W^��ތ���9�g*""�v]���u�����U6�U�v`6�)"����^[����3��}�<����G~��~?����9>���}
��*�����A��nÅG䑟�A��y��ޢڽ�ރqt�U���_�����s����s י�e�������fV��|��[�rۚ��6�W�߾��hϛ0��7����
*�5M��pX��Um����q8צj��n����xUASC׍�ۧ�Nב�BHe��
 a���"��V\�:���U6��F�F~�/h4M��g
^#cp�Mҗ���5��c$��ƭ\%��Q����}u����sx�����4�&�AH��Z���F��ܘ�(~�\�  � �(~}�&��j�
Ԅ�Xa0y��'��|��,��y𪊥";�R�����KG�ؚPZ+��ҷ���YM=�� e湪im�    IDAT�T��7i�B��נx�}��lƚU�)A(��K*��������lR]c��m]�ԲP��U������0&���0��D�OOL��[C�f2����*���V�&uRցFc;f��M�R���C*�M ����*�:��Ezq�Qi��Z�=�o�1Ǘ����w���}ã!X3Y �=7B��eq�����Q�S~-�/�HAi����@���V����w%�Na�0�=-��8�X�A������gY�s/M��Q���_��o�z�*���c^���98x��`ynɝ�]�~����WX����}N\`o��3G�] ��)E!!��Z�v��.����&�gvR�T��O条�w�ݚ��cg3�|�˼��+T�~��G���`�K/��淾��?����#��S	�s�v�6��^i�չ4�x��M��Cf�+=�����-���KTf��*�ex�ͬ��Qb�
����<M��}�scA���h���r���4$�Z��X� �����M]<A1�4�T�9��E�Q%6����Y�;���H�&+K��R�j$���<jt3m*�=��n�bqi���Ȑ�zBU�=�W�0b���i�L2aOJ�V��"}�:52|��S�`��@#1H�Q4�2 @�b�����RN�d���1c�5�䃍"`zF#�5� g�!tUH؈���H*���|D�w��(=��t��M���^���cF�^ (��ɻ��2�PX�B��ҝ?5���9�{�oqH����"���
!b����%��[��x{�e`@�=�(?=$s� Q@��`J���R�H�gt(�-Ƃj�ed����&�	�P�� ���gl�šBYY�4���h�.�̏��qʊX��N�=�����w�l俳��@gT���Ѩ�����M�<����¯U�y�f��̰��٭�NY=��|���c���w���D������'4	��\�]Z�N��1�J��l	�.��h
H�î����ڷ��k���q,ko��@�����<d���'<�/�)�wpb�u���"���kC�����x��	3S�O�ys�	kzM��x=&1��E�:�H����CbZi�m��v���1+F�|��3��%�ޟ��!)�f�#y�[!��넀	C��L�!/m����Vz�\��'++�7e֓�4lа�ާ����	GVV����O���_!5��%_)Z�N�ʔ n3y[,� ��O�El�4D�O6������P�M�G��������^���Ӱ.�[��H֞3���g$w=N�&}���E���;���$�ng��U����	�9�4�0��52��"_Gf�3ĶK
�l;�����NA�Ɣ�X�q/)5�K灢�6Z��e�.�����N0=mXlQ!~j�^�.e@#&�Y���;Ef���t���t����3��N�T���p�4�d����1;j#�F�	��1S��do�ύ�!"T�eU�᾽s����"�5޵���V��-��c����Κ�'7�2�OI5>΂�"S�~rՕ��#Vg4��=k�9��}�7^���%�k1T�c�f5��p���W>�.�F����kkt�8~����nc1jX�V�1t�b�ABSLW��`vw�1/�02N/��Y��=�3Rƛ�+B�s�yD���3㌡ms�r�r�ɥZ(_
Cφt�F�FWrt�+�O�p s���`���c��QD8�ç�I���6Byzqф���#�f�9��D�Y3���ء�����w҈�kĄ2�J�L�R��L�0��T:�����-=��ACLI��n�LK�0F��V��,�N>g�Xv�������ݡd<2��I=��N�ߪɌ�z,��/�L-p�L`>��R�LU����sg5���</�w����=i5Q�ġaM���K�GN��d��%�9�i?�,�x��2� �CWŬ)�r�~k�p���6�U�ƘΫ�|DS'4fP\�k]zZ��E[+.x�󄠈�(ڶ� �T@�!�dRo7Ufs����:�Z:�p�1����h��:h�NJW��=)jx?dMd<<K �p{�3��0u�ߴ���yݰ�X�;6��1�?8��9�+��p.���jF���*�@�zj�p1t�ۖY���.�Y��U[>�=yOR
\ĵ0:?�ّ����S��r�����O�)1���a�2����~^K�9(a���w�d!f2F
Ƌy$idYk�/Mz��3�(�yQ������h<?�6�ƹZ�D�1���0e��"`��I����ArĢ�Bl�� {��|�Wa�T���%�`B�dp��>���D�C��ˠ�DA"�2�3�5�g&sJ�D����KEv��o��֚��C��vbn�G\
�Qd+����O�f �s�b^CTm�2��DoG��{��.q�����pl�HOi�e��s���ِ��G�ǿGU[&�����z�H�s=`"�p�O��R��X�ςS	��{�d�x�>�8ߛfA�Zd˾�{r���e?���F��� �� �!8%t�؋cP�����Fb���)��m�x��1���1��[cM�x0.v����k+�R�b��`��w[5�w�n��Rճx�9Z�Ҿ8*Yҭ��i�[���b��{�<�x�l\`#�z��S)TM��u�i{�$@F�%��ٌ�_�V@�R�Aŏ�Fz#��\�R�֭��o)?��%�.�H�˔���XQ�0��K�[U�7�9Ee�A�FO?DݗZ\p�5��Q�/Si��Jm<��l���8^X�U�y��$儐�Rz�*Z�)��K�K��n��!z�Ǉ��jBxP��V�`��I3<ҿ��$-��]��S
 z�RP^b�3�^H:�A����e��Ж��"ogE0�4=b庡\m޳����$�H*x�`Y�4ǲ�_�_?�X����0��IjM9�GH���h�3��Or���/a<��m�?��gae����Y�Ϧ��t�OQ�}�^:Cy�4�G�Lw����#����șk�odd�,��b�H�-�����{7� !��K��2->�h�~~�Cq� �|�}��y��IP%u4hXQ����X�k]s|�f��1X��Q+X���4g�j�BKO�{ׇ�-��m�~�����v� f�<�8+�X|J��.�Jf��'��c
m�=ud�jT��5f�Xa�Y@[�8Ϭipm�.(k�6��Ta�SPX�"k�y��Hnn=��dV�g]Kr����m0�O����mV�OΈa���l�FW����
NB��K��MD���X��0%��[A�%�a��v80��\���6�e۵����	�mFH��g$PU��/+���@|ۗ�b�B1Q�C��~��k.e �iN95CDFf�Ba��� ����N�����|
F��;�7�,M�3��p����0E��~�BH���
"B�b�V�ߗ�8����� 2Lb8�cS2�%���4n�O��ʈ9L���8|fF�gig�]j��[�If�!�(h!Ȍ�ʼf��;���Rw+a�s.�sa���/a�)�;Y����`q��� {s��&H�-�$�#�Y����q��Y����0�*�~|�Da�F�:#�S$���X��(�;���14H��]��ǊPױZZG��.	e�bd.�����H1*?�<�,�����"W^uUc���t]
�6�Z��������n�Sefp����t��*j*o�@�:lUG˦�x�w�JnQҴg��/[i�>�5��y5���T�J>oy>_f���L=��\��4�fz�9���|��%�(���>�0TJ�o9�ؼY��sZ T�@�}֥Ij�p�A��>̩�Mk��Y{F��U�4����:�sTs�|�z����m?Ŧ~�is�S��� �E4�����i�HL(1��\��U�!@L� z}*Ѐ�9��,b����gF�#/��'��'��Be�s2��ZO�UO��0sGm��3қ��n�~�������� ����t΢%����4������宋}[��&��s[��Ո�B`H��a>��x���Ê��D��f^SD`Y�=nL4u�6&��NϹ_�����WP��K�C���VN7%�J!�l���m����~���������A`6����fk]�)^R[�ڮ%��������6T	��-xPk�eZ�^'>Vz���8������г��xou�a4�
� �V��77Y�`B�ewg�r|t���kq�JY���Z ްZ�]UQ��f���kDR�ƺ����]ÆM���:��Vf�Y���Fi!d(ʔ�z%�Z)]��aVfٜ��Fgۯ�
B!��P�ҋ^P��l4Dc/,����ɋ�.�� Fcd��04�|�pT"��/�����Ny�@�n�63�����h��� �{�m0���a6��*k�Y�����hN�y�u�!�9UUE��E$�d�U�O$�<_IE�M��4rd�q�!־D;:�!H*���-5�L��*Y=��̀:DY柝��p��\��ѻ�H�
!�گ���EQ�Ǜ�H 56z�;�(@��bоpR�2�9���7�$��Pi��M�п`N!d�H"#�AL���-����_]b%V+�mb � P�A��,tq1Gׄ����[��/<���/�W���Ѿ�V���}�t���)d�F���B%Ub\!�c��EWָ��FgN��2�ȁ����UrF���'!���Yr{谦��3���hza8h�t�^���ArC+�F��$!:�h)�yo�Ƹo$%�i�^��
�&e�	���Z�,�7�4M�+R�h��sD�������D�Q�����V=�q11��w�fFc���	�E�}��EN
�Z޳��g͢��h �
�`����,�;lB��#.�r��
3q��/��v�u�5ӵ��u���>�:�=��¦�S!le(�X�o{��ު�
L��J�Fx$���~/�w���)z��9m~����̛z�ؒ6��0�%58Ӵ�$,w�%��.�d~T��I4k���M'_JP�Mg=sZkʗ$�,���RD����G�N&�����]Ef��i�4��nǐ�3D4g�%o[ԦB�|"!j��w���/?��,�T��*h%���!ˡ���� E0X�W�^G��G'�aq�SM�$���A(`��P��5�^�<w=��M�͇4�,��;龕5�<^pmJ3`���j+��{!�qPG���fl��:�/gp�.����{�����݈���,h�7��S��3l%�i�K�������CcƱ�C^M��M�%�Tf&$7:������Y�>�����(@��n�1�!�>'٨�AP!`��@�'�#Dn����Bgd0��ۑ&:��1!�7��ˠ�T,

)'����cA5.l�Y��BJ=�#�`�C��-R���\���!���ͮ�����A]H�؀�"���2ۊ.gސ�F�3�ĺ	�z�Q��rAzd(F�n�pk'�y�d�DV*���:��8CF�U�m�'��FlLq��P�3M��fd�^y��1�1i�9�j����2�0"1�Lu6���o����n��U�����E�C61���3b%�> �$F��T>k-M�P'��b�/���)b�sf葐��l6.���_�
ǟ:���9/��E�����62q/��1C�aS̫��|S��Ϗք����ZY?�YϜzm�B8�Vy4��ؿC1RE��hT�%ٰ̏�#�%��3/�y�gf�X&U&�{�s�=4U��[��'����g��J,e��Ks�a�~�ʐr��a�UD�杪�eKSI�EHn�`C��V�`���O�������Ĉ�r���q6���T�K�;6Yx�Thj�@B�j�0�5f�ы�"=����T����O��;UM�ȸo��<=1����oo��"�!�c��s�?�O�s�f��ZX�b5�E�_������Ć�N�@�1�`L5��4Df�^0�k
���(�7���#@K�+8�t�h�a:4��/�ջ1�L��S��3TcS��,M�@9u�ƌ|�1K�:"��¸(�=NB{!0�3(� ^A�'øw]����,��׿���g�"X6�W�X���J@����x[%��N"�����w�̉�R���AN����i�
Ӌ���Pr6�DI�Gٳ���`�!�L-����Ĺ@�����5��ȁE��B�hp�&Ǐ�c7�`�+�T ��wnI7��J�"���ǃ͠� �*�i��͒s�ҳ(pCKI���g=(���N��5��T��Ϝ�P���>��L���"@F��%d�B��b��>�T����q�����	�DCtW`��0Ehs�>1��R�H�u$�7U�����1D�M���e����X�\&��KsL��ʢ�\-*�,��
�(��S���|F`�O���A�s���lnV������ُ�����f����0P�qK�����G�!ƚ��b��Г����ݦg��2��>�C5
�Cy��
�`e(Ϡ�8�k'[�����I:��3�}_�9��~��t,�|*�L�	tܕ2�n��[���)22��6�qJ�ma��&��TXp�PC$�����C�~��OT�:ҟ,@ga���q��l�0I?Mɦ؂�w������H��Xb�4������ݣ���
� �E�~�^� `� - �b�g����23��^3#�@�̮G�H>S���~�yxxH��9�>r��Z9�l����F� <�{?�q =F
=���Ǜ�WkIn�	I�ɉNptJɴ�G~�J:N��A��ч��D\�g[M	C��Ci��' Ɍ�>��)ұF�L�mx��~�(�����G,�F�����PV����m|��;�/�Tn�ÈtOR�ٟ'��/�ww�w��f�g�ObD9�ݣ�����"Q6�\�&��cg�>�-�����\t�[��|TA�a@��Ȋ{��+!����(Z_�W�4(�E:5�O��2�a`ꒃ{�a;�3:�+�h�Jk��!(�d�u�^��P �NC���F�C�P��TN�[�u�4�<lR���A؁��v:8�b�����?:T�����:uB���/��҇�x��e)g+�Ɯ1%?�	���q�12+���[�e�p�}� ��n<s��ιI	�f<h�' ���].���}�lY��N�Hɐ�S�n�������݆^�_<�?�s��� b�KN|v��(�]�4KY�Cp?�	�8)ƾ'/ǃ���qp����~�#���ID ��o��^V^'���2�:�vD|t@�?��?������w�}Jɔ��6Fz�����{�g�����(������@����F�|�Y;胛Ï9��qY�X(1A�M?��Kc��؜1V4KE➤��!�nl����Fqsn?�۩(?QPE����u���8�z��[W ?��Ǎ�-���	6�����Ά��C? ��6��P#�<�cd�4�YP��@��J82#��CWS9yCы�H�Rt�">����B���"	��!�$vO����$��vT�r6ҽ��{`�v�^)�����Z��ܧ����PPN�@뼆���u��AQ��b�
,�c�:@�����rms�'rM�D�v�9~~-��#:]̨G���Vܙ�~}��f����o�*P�av@���r4�#����2�7+Rv���x�l�����6�1?�	�`|�pK� [��y �AY��.��^���B��l��g	Tr>k�JW
��@�L��5&Ip����Gg�8����)'{>��N�$�>����60��71��A�ފ ���ݭ7�z?�_��Cp���.(� �<xS$�`��DuD�D4�)Mo�|M'䉱�C�����Ä	���`M���N��A�?�>�}�R>�@�"�piG���=�Mon�Λa��u�'}1}4��oc^�� �Au:1�����c\�ł^��;j+�L	�Sk>�2�����'���]�^��\�v�\`l���I��ʾd�7p�`qc��Z�C�?������?�����A�ܙ�)�P�s�"BN1v���9�q���g��{w�)*�y���`��%�����"#    IDAT�b�7�cYc����\���Z��:TfosmF�G��;��	�)�hZ���X$�{'Fg]S���XO�΋�X��m�BUL�Z���C�6�ۣ��;4�_��Mr�;C���Z)���z���}D6\�	�[u�� ��O9p�UZ���e��X[c��t��Ck�U����gaMS��p��} E�j�V1瓃�������!0�Lc9Y�aahü��D`c|���t��pL�{3�������{�?Z�
gc.���=^9gl��ǩ���٩d����dm���i���6�	���·��F�p(�RR3��%Zv��B���3^�c�V���g��	i�sla+�f�4�����B�Cyx��gG"r����+p��
��g-5Q��d:W��h���P=4���*W�Ίa����A[��I�#��|�E�4���d!'n��)l�(ሰ�H��}�
px�.�A�"L�$����Պ�*l��R"Y��o� S��6á�@5�\����gҫ�=z�6�/����U���X �T���2dV�2�z�42�Kmw��(��ƿے&"rV�s
H\�a���-׏���va8��_t2�T��hvD�e�1��6u�Fn{Ygs�O�y�;|NE���A	�p}Oj�2��8�j$R_0'k�j������{#��We�>:.KM�;�f�Z�n��,���k]>�he!�>:1�q?E�L�|l��"����}��s�~6�M&��:���_mNʇ����s����QN�=V��f��]����g��FQ�+���t�ugԶ�Ef�	�BG�ָ ���l9���,_3/V��u33(g�.$�Nu�:uBa�����z�"As�^py~������X^כ�o)�(!U���UpSE��;���?���_q��P�H����ޚ5q���=�C� g{�.���p�Ƈh�n��r�6�v��@����w���i�"w+c��*���ؼ��`�*	_�]�MF�y���B��4���(z��)1�r��0 wj��ٯ&�.��3��Q���hI�`�i3�jl>!c�����յ�����4 K���_�J�G�j�~;�	�l(�U��q8�����Y�8ٳz�U�>�ʡ����p��p� H��*���tj�KA��@i$O�$F<��lƲ����Xf)�(���M0���h��)��!�g0"����4�ӈ6�)3��ض���Zt7X�ε��X�L��/��0�)_ 0&�vw�|�[kPG���`�Rpt���r(hK�֡��PkG�^@ʨ�Y�^�Q����W2�2;U,[���j�ɮ]�E���N^ƌ��T�ԫ�������!�I�nN��j��Q~��{��ooo�r�t��$ ��+)e���lA���`x��O���c����Z̰}�b��e LYwCU��I)y���>˶���l$��ɷqm��ө�t�L�3;�����"~�vAfF�t`�# 1���Am ���*�w"�*A3c+�#)�$8�qX̩'����:G�3���lz��H
\K�1�J��>D�l$6}%`�^q ��Ղ�C � ��ݣ�V�`�d��G��ߐP�
y��A<����c{2h9�hḲ&�v!�����;�\�u�S6������n��V�� g�@ZOx�����Ě�$?zj�<��!e/wA�~�Q��.1>N�����\Ԁ2�v��q�D>ϗ&t- �+F??(�8�8p͑�%�].˦ѱ ����(r�h�9JN#�!-�B�+xx��LeJnP�3TGe�òIeB�s浢<� p�M9�C"�B�H'A��  �w��Tf�'�P�w�ȕ�@a�մq��g.ڌZM�(��yc7���9X���g�5��`.h�Z���y�cs�\�NPZ����m��"��ldґ]PI�/!>�����`{t�8�����6	�ŮM���FG۱�l��"�I@�� b<��V=�4�pGC�&F���$�Y�!0�TȤ����
�^���&���$��"@r	Z%�9,�w�趔�.v�
8É�@�
�����D�h�&0�[;�.��k�è[�CL��jx�X�o6y�6�V�^�!V� #sf2��{�`��@*	�a��99=/��ש臭�ަ�Q8�#Y"�Q =Z}���*�z�5g^�uE⧓=P%�6�D�T�G:ɜ��5� p6���	��v2��ُ�%!���dG�zJ����044��[F/%�����@��߃�D���f�lrNh!>A�˚�0t��{�����|=~xr9'��W3�M�F('�1O{k�D8�������VG�ތs�A�zN�֙à\=����/_Qoo�r�P�М3���e��#3:�gv뺘��̐G.~�Hs��ilV��"�ɠ�1����b/	{���duƦB����N�PG���o�Y޸Fk1��T�/ش�{������� �;�G ?z�xߡ9!-KŖ�Y0U97���6�׵��$2)T@,�(��J�"e�#I�Y��lh�LU���d�>��V�
�^��{�j������{��ٝ��@�&"��n�}Y��O ��:��b���8Zw¥d����q���M	G���[�5�NC�� �n�V��[��b��^�� m��^�|}��<-#w�X���GN���9�X�5��G��ԇ���f�b�`�p�H:
1n��%h��l䒑��`�ޱm ���������㨠��!ӅA�lG����Rg�&�u܉G�s�&Pe�DeΚBXQR#�*�RL_�h�u?EFw�՜�!���wCcΨc������B6P�����>]+���߷;>�'�7@ƳF
��>WiiC[fJf���y3�Y�q%�c�u�y���6?;v�ws�������m۠��j7��BT�j�2�<�(�[-@6�ު9�p�.�� ����6Ќ3�{�S�_��Bnr���+�
T�w��GC����A�O/S Y�Ŝ�sB.N@�2�-v8���)����+^��YT����u�!�W�{G�&��H���j�ʶL���/l^JD`�ٴ��d)��5͉�m�^6#��9Oeu���Σ��z�U�* Sg��|�޽��u�Bn#"�H1�� ˵�I\�Z�wp����Q�;�10��Ύ��3�_=��~<w��p�9��� ��n���Q���C�⠜6��D@�D0b�w'&�1��w8�S
�r���m������R,��c<��N��Z+SJ`'���=�Y�L��o�����'\�i��v�U��S��̜��t�&���rI(ŌZ��R����;�6�l���;R!���I���P�/��V �޲�$#�u�@O�		�u\K���97碃����tttb2C�͉�"h ��!?mH^����� �]J~o�����2(w(
%�PTgAuhjv�DC�k) ��(?�5L�]�v�5�ۻ�:"����L@ڐ2� � �#�֠�S��HJDF�+�{�^v�wyC��?_���w�ү��5$O� ���*c���ɾ)%��X���� �@ɢ{��gL_�U��q@�5��~&�1��&�m]W��h�91��:���D82���J�8c��9c��i���Yp�c}ϒ�����5��Qn����8�������l.���� ��{Ux�+�5���y���K��<,\�z�����z_9g(�P�Skr����Z;�����p����uG���V�s��_�b9����ʞ/��}x�� I�?��0�Q��/8����L��d9Ե�	�Q�+Z�=���mТ��a6Q�L�P�K�ɍ\�y��is �����ȼf#���\U������k�L�e���0DF��vsqc.�`{�(���B1�T��J��aV��2J�b�VX-q"Oi�N��E���(G9"2�Bch��a��K�`z��[+���w"�*.x�$s*�o߀���!طY>5	Bs.A>L5'�vk���5QR�y�d9��8�D�mk�9�JwuI�咱��g�qTGE�Q;n���H_Q6[W��g���7ʟ��;�"ؙ�f�'d9�a7��L��}���v�X��U�%���B�q���w�
�:��զ�(�v'�zΓ��������}����;n������ �6��/��ۗ/x~~�P�///��n(\Pr6TQ+������1��r[�W;��0�5���?��qX9|ƥ0����E�`K/�d���-�i4{�eS�/�Xh6���Q�*Q�T5��UG$�[3\1�P�H����Y����Υ2�0�<��z3'	0Ni"HsG��^Z����0H��������bj�W��W��H�v�#���h{yƏ����ϸ��,t��vC�x���o����m�a�U��'N����-|}ư��b�(-?7�n�����ٍ�Y˗��4kMil�x�ox��7%��>dF�jz�2h��A2��O�n���6G�t�l�s�h�����R2Ja䒐[���1��@)������E�hn�uR⠎EDoa3����F�$�b�*<��G��ƺ�W1������	����f]������8�0c:a1�����g7�v���Q�DD����q��ĐK���E��˩X͵�~����h7���[�cYg16aD�݁.��:h����@�'�u�B��-�7�lų9���n�:�R%���^1�p��/GɎ�@�WD�_�������M��M��j�wH�͊Z#�d��ao�%���ĸ�\������d0�/�����]QE�(8:�W�@m�A��`f( �[~;����[��w2%#��\��g1�Ug�'��Rv�ځ����h6Ykuf��W�gTvZ����nJ��� ��F��:�O�Ƿ��@����������o)���ߍ@!�����$i�t�HA���MMc:��>Ά17���ׁ(�噶3j���x��}τ�cYe��`:S�v�k�����i�
fsJb�[`1���w̃v�˲n���J� � �Y���?����X�·���3ǻ����@����6���Z)%Nx�W����Ox��dN���ϟ^��� R��j�qqB���BŏX�"!�������,,j��S��o����߳�r���㘌���夰���K�{+���^EJ<{|Ƥ���F��c<BW�~�������w�����O��N��<�7c���;�NH��h1*�TŚ�IN��U�ci3
�ذ�ߠ�"
F�-w��̖�����&�D��fx�F0c�5F�f�n J9	.��@�f����^"4���L(P���C%-hM^����[�a��d�����5(wO�P��% �4Fr�  g����i��ס8�|"2�5����a/���H�`Pݚ�(��P6�N���SA~@1AdN�H�.�l� r�������"$��J����5rZ��w�nw�	 &\�N�ׄk�z���p=!����u�!kC)����j�{�3ZKP}��zE*-�^}CD�`�ɿ�V�;23JI�vX������P��t ��+f�S�Q����r��׆�8F��֚�&��e��9�6$�u~�E�W��8䔰�+jo�v{�O��������3������xzyƧOW��rb|���H/��A�w''t@��8�8#s��w?ܷ���X��G����ZW���*\/� ���(�� �^��)��6�hDg'$ C���6��0�jG���>�K���qHH��#ؘy�H���������P��v�.U�6��w�m"9��l�"�1*8���!�������ҹ 2�S�������xz����;�\
��`ˤcߪZ�E�3&�(�����c ա���'�_e�I��V���8NY���&�/�����8�o�}@���������o�921�x���	e��j�ߵ�*p��E��K����׋�6���p=e4# J�w�1���'t��l�]/&�::l�r=��܉z�v�=�4�E�q�^�o�VI ? ��v&�LF����lHM��|a�#J}8�<���~U%h�Z��U#A�LD������A��P��Mi���*�k6]u�Б��ӎ^j��1�cԲ�Ch	�c��q�g=w��ɟc# ή�.�y6d��<Kyqv�Q{��W'����wU�5��mL=m�lH�-׆���������W��V���|��d{��8�dK���;�`?,��@�-F���x��'\.WH���Ў�[���7����>�e�������Yyuh6r���r��pI�Vz�q���|��u0[�u�M�Hd���hM��ml����L�D����;c]p;���m�� �t�z���v�ض�?����~����>%�O�=��@;^���=v����Pu���=�R���R�;�����r��6�7���[���>�3$
��E��- �l���X��zX�s�p�Ww�u��9��+T�M(���8E��L��_P�c焾T_l��V_ޚ�t��h���ڸ������)�z�I ��<�c�^�F9�M� ^���itĀ�lU"�[����(�)~�G�����������~���G������gO=��X�c��d�'!KFG u��\*,��ߊ��m����x���U	Xxe���Wθ}�Cs�ԙ�"5a����o��KY=*$4$$�2qc����<%�kX�D��x�l�b�C �j9�.��mG��W1����`(r!��H��\��sY��D�ީ�{�&~�p�C7T���t�@�hL�#�W��:0��}�%u(}�8�E˃����`�$��b��"D=�X���w�1�{F)�����p�ߖ���vMCR����7�y�V�T�,fx��	@dK��t_�F,�V�a.Q�;a�5%+�S_�#GO��� :R�H��n\�{X�W��ބ�֊���^�}計PK$�S`��ԑ!!A���m����W(��%����V��N����^m�
81���/3#��U��6\Л��2Ϲ�1��3}B����'�����O�	?��)�ʆڌ�B��wq���&�+z�u7#J�+�p${�ш����(C�pH�ܓ������-��*O6U�~�A��g�Tj,�!Tk\��"�"j-X~�����Y�a�;�5<��r�����\���(�H"��W?�o��_q��� i8^�Bަ}���]	#�����47�U=��ǚR{L^C۠Z���@��Ti0����!�~P0h1)mȻ�L���
�d��p� Fg�Д��v���<�N�! �ͯ�)�DC5P����d��e%k��#�ł�>�����ɸ�����y����I�l8�����}�H���M���_  ?��w������_�2dM �� (@ʄ~���-�����`t��<MiSU��'�PXX�]Vt2A�ڻ��F�� �����w)gפa�/��"���g"rr�C* vt?6H�l0b�l���)�����vǠ+��h����  ���4 �t�`�w���&(+���,�s@ᑷzȵe�@J���d�Nv�Ӭ#�9��U�w/2��>�X@D�A܊�&�?��h��X�o�BPX9�v��QeK3h��tO�� ��!`<��$�G�CK�I�q�3�2o�Hs�di�7��K�ziC��D<R2q+OOvPb�2=X���@Nb6���?~)/���PwxI�0R�W����S�dr_�s�����!	����K�Ag:��s�"��$���v?���������3������������Z+���S@S�S������`J�|1�wI9�6�қ�Ԗ�>k͏���@}�k�s�S^X�ȫ���b�ďvۍЕj�����lͱj���_�͝��g$$����O�B��n�kQ;�u�n_��݆�LQԶO��(g�}l(D>�r�6_�S�	k��o�C4�9��������ў�=�����Y��1j��ľ���$�>�����ZO����Vpd�{���F �2o��b�е{m��+Z;�믯 �?=��aŵf    IDAT?��ׯ�P\/h�*	|���ۓ�&G%)��iST	9gC?#�7Ҭ*#�����/��'Y������3�b?�;�m޽�sɏ�� �7��ƟCn�fÕ�
���a�@eA BH���z���G��g
���K��SJ!l���v��e�,-uB'�H=ڴ����7b@�`{tzX�����s��������ߌ(�!�1�?����o,Z27 ��9���Cǿ4�����~Y����Z�> !o�6)�I.R� �(�SS9��FS3L2�^aez��&h��0x^^�s�I��G�&ꅓ�j�ψ7Bb���<��>��@=s4|��(*�98ϭ��/k!�+����Xӓ>�#^�w��<��չU�j�8��j�s������xI�����O?�� ��[|�����7�# ��ik��߉�� �ߣi����@�;�x��s%~t�H����c��+ P"l��w���@�^�� ^�W�Uu�^������@ �8�t��}���7c�ݰ��@+��r�^F��ԅ���Z]X� T-��r�)�%�c���'�v$�vbHNe�$Q�.X��a��YY���<�8��ͬ��UnS�U���p�	Ȋ��c\�h�������`�@����1�f�����v��� e|��{���O�����+>]/�D @����r�`x���Q�n�x<=/%W=����O<�#s�',[;��-k-����5�? ��3ֶ�7�ҷ	.�����_ф&��:C��YLFCf2r	�fu�D������ßH�C�E���a���3��d2%E�0k4�P9�:��7�Q��iU�;��x�ǧ������"�	����Qbwި+�?�K�:vM�\N�R1�T�IHEܿy��9z����8ǳG`qe�G�9	˂�;��7���|cS8u.c�s?�'֯�=&�L�o U���ad���������u����Q��])[Y�Ґ�D��w�P������C ����ˆ��'�Λ9�s��?�g��|���JF{�#��nС9랎&*�rd�X�&�ʊ���5��5�mH�e�A>�[���`X�˟v�Ł𔇰;���Z6$f�0���	�d�^���='%t�9Y" �!ok$ޙ�	���i"Vv���H�0<s�LW��4�[�v�:�S�﯎�d}c���	 l鷵�mL� �ѓ��8?�p��w!�f(�FN̟ߜ�8Ё�a�F�f�wo��A����#mf�j��
��	a?:�02]�U����B�?��;\?7�����M��}�n�6��T	�@�cs\�A�GH�N�+�E��]�6^�u�GD�.�ә��I������sB)�3�F:�����"H�:P���ѵ�~��������1^2���?�f����T2��vbӯ""V+�'�Y�e��Qt�u�G)�O��Y&bc�� .��2�/����\eֹ�-_CD�2L�Hh��m�1o��;m��ВXO�^�u�$�GZQ�	W�����>M' 0��/c}6Q��j^za��]��]]��GB��}�O�o3�?5G�$gC<�����\�4�}�.��u�#1OY*�Q^h�!E]x����c���T��#����wT�K��*1��������� D��Ͽ�	���//�H`���+^>�jf��0�x���q�l��h��s� �̣S�ͳE)�Sg'���B'vg#D\��ǡ�n���G7��m�`θ�"#�s�y�^��J�C�!��~`�Bw1���B �c������9wz�A(8V�."�2�ѵ���u�S(��A5�r>;��Z�C~���y4��t��֪i�h��p���^O2侁c(��c��x'+�lp�&_�n���_�k9m d�o���߿��w��>���������8��y{��펴'Q�(f2!.����Ï�<EE�c0�!�܋��jj��:��+C���I��A��;�>�n
�..y�>��n)6�2�d��8jGu�"[��nQ|b�-���b���8��{��PM�|����'�皚 �k���%B6G!A{��pIU]����ڈRslVǡ��պ���}I�s�_�)�ń��=��p��t2����Ѱ� ��S�j��}ξ�D L����8���}<��q(4�{RkR�q/�5S�8��D�9�ҍ�g����OT�(}ql0���יd*���/7�){��~� nS�L�ddԒ�����bL��6(�mzY�z �=��m����U������� �csu��[��km`��@GQF)���\���� (�#'�c>�3�/c�8 �}��ŧϨ�kF}�������Ok-�>��V=?'Ԯ��M��d�˛��L��G!�)��0~?����e��3�FD
���N�(�X�(0�p~ҴaK�\�;���f"���#`*&+��~VTG<��a`4[�C����A�$���]�l4�Y�.Ӧ�� �/D�5x��3��M_�Mb7�|�a+�\2�M�Z3aۮ�ow|���?���O������؏#BҰ7�&��Db��j)��Г��:V���Ε��2��o�7����T� sz|�ѯ
r�z3�	������d�O)����T�0�g ���p�W��M�A�����Ʉ!rNȧ�4��1��V Uq;*:)�:h����kD^�;�q[�m�w�v\���-�{e�&)��{1��[��rG+Ӛ�Z���7A�uH�o � ��#!���<�&�,0���4��{/a��Ѭ'p�s�&g�Cာ�:V�8����,_� �FN"c� G�q��6J�z�f$5�F![���@r�ndC��)�3��r��'�C�^ �q��������C�s.����2��p�j!������m~���UeJ	ʕ�v(�a�	��
p}��d'EҎ��@�ݐ��F�M���^_o(e�W�A T�+	kp� �2E��e�N/�~p}̏9釶QU2����5��y��uqxӣ9��6���l$�f� ǫ3�u:h�S�CDS����C��5��FEŪ��<�Wk�ð�X�xU�R�c�h�3�4�%��P�eq��r�U��9#e�`Ab���H�C*%�����C��gh~�ךnI�y�<�4�i��B�?��ӦV�D���ؔNY�x ��<_��2B�u��@Ҍdeȩ��x{�hU��D*����8�;~���Up�~�Ӗq�o�����M*����(�-���o�7q����͔)����n��"���
�X�11X��N�
c~�������>�IR
i���5���9��{5��L�#��ַ�4�,/_Jq]�3<
Z��^o��_��w�p����>���0�RJހ��߿�nb��sJ)�s��~�H��� ��^���A%"��kx�4��{����6s��,�� *`*��!�N�	ā�8Ѓѣ�M��`�9j��<���T��x���yԿR�s�<r�u�l���b�9t���@ɗ1oo&�a��5G��8��7t��6�@H���Z�8�;@��1��G[�E�+4HW1O�3��-����U:��|�p�^q�\����+�v��������I ���ڠ��~�7NhM����}��Q��/?���H?�'P&������O��K�P����DH�].�f?��'�Sc��*`F\1�O/W��gn�]�|}>�@�	�����I��RBEŖ3�;�U�`����0��[D�2��pH��X)j���BS�㜼K�L���ؤ�׵��]��uM����:�u�S��q� �ɷ��|r�Wa+ۏ'<����%�Q��$/��t2^�f��X��G��:���p�B�
DV.j�cx��0�^U�i��7S#�)H�\��7��c�\ѻ��^Q�	5(��\ʎ�������oH���� J�Y0�1�vk��Q��n��n��ܯ�f�J��F�HD��+U K}�\>Aߌo�֜�1ٰA��j�c�(��O��/� �Z�?B�oVӈ�H�R�V��n
yܑсDض��Z�e�L'�h�v�I�m"��zE��__��@�W�$�j}��t�#�-cC�Z�Ur� �b������y0�"�O� �Ia�����m12%t6� ��!����_�m�	�|��0i�V'�?_���.���'&��z��.��JN�k�� *�U;�E�j}�sq�C;����7���:��{+[��9 ����� <8!w4w&��$`YA Oys�'��z$�F1|k&�wHD�d�4�5���~���Q����-��*�Rr.���P
E�v��P�;�7�	��ʄZ+69N�;��b�t��Q�R
��.})�85H�.��?0~�����������"߾�A4�肿���4�{EO�����VA8�+��]�
DE[���<�*�p�s��x{1�f������@)l�A.�׾����@�B8���8'���M�	[�x;�~��M��!�ĥ�;��Z##Z�_/��}B��B��_��RxFYL�(��V j�G�t�+>�ӆD��vT��ز!��5 YpPҔ�^9G�O_7�"��ȱ����e\��h����$����z@j�&�vy�F�� 6f$ڰﶇ����D�����C___�Jq���6�����$�t4�R�ki�&Q̌-���Q�l�T�~ʢ��Z�j��:(W������|�~W\sB����\�)�㸽�W�����SF���7Ho�nL��ʅp}���v���kFM�nN$Q�lح�6����Br%�.#�'�3D	��rj��J���(g�ڑd�3���/�L$/e[rQ"�R��94-��bqmv�����jG����=�@S>1!%#�Y��}g���ȵ~��:G�����td�[#S%��ꍈ��Y��3T}���<Z�[a����g��c�I�
u%1D�n m2���D�
���;N��G����(cn���ye�˶�5#�@X��`�&��<�E� X�II�];�-rȄ�^�g���֦=�l|;1���X���`����{Mzԡ�4�f����3�@HN 5��������5�F}*���1H��V�<�bvg�9&�7�$$�<�/��%�4DҭS\t=l(ܩrIM�֯��SZ�ZjV�n���ێ������-������>}~���Պ�^���	(t�U �,��}��+/WV�\�VEp|�N��2�8�����5
��/_�HKz.�iD�fV��蔆#9RgK�%�[)���ڼn�Ѡ�[AVkt�5��>�V��5kۛ�۾h�ι�4S�L�,�h S��X�X��yڤw���!�����~�`��U#$�v3h��^B�n���;��jא����ur��}�A	V�O�����>)�T��dA�*���qR%��Ο�I*K)vл����+H�ʎe�+�-�������x}����^œ2����;Y6�#v�7�s�w�xP�X���m%�w�S���m?��%�V�/_�*LL��*�9;dvv�2D�7��:����xee����oի��$�hiN���Gvc;0�pB����zt�i'wMH��C@�Qa�R6�b���h0v���R�}W�z��ێ�!���@l�uB+%�䄐�&W`�Q'<i@' -�pOd�����L����a����Eg�5�<t�NƟ�����Q�Q�Jr)gC�W�	�w��R�ɊWژ��B�r)�̙���@C�2�q_kd��nM��*�Y1������X��@��C�L�h���-'�%#_����.mD�v��/��E-t̩�Nv��W<u����io�n"(N||"A�&'�Fo����9ä�k)��� r�#�����]a\,�����A"��+��u�:�����'Hk�>��ޭ�H�qF�*4�_Xq*�#������0���!��:��P��	�;�W��i�&{��Џ�:~?���9�v`���[��w�_xC+�C֣]�!εi��ʐ����*��_�Q�����no��!BhG�nhج���X�e���:�+����b�*wt+!��t+�NG;^O�a�G�Ct���>85$���i_��=�h��%Oi�#��-���?S��u�]����K9��^�s�3��R�ؐ�H��g7;$�[E�����=�����?����������ׂJ�g@��|ɞ�'���YZ�U���@W��>ٻ���Ul_uEw}.Ɉ���l6稛�T��:���Dg��׺�� 4^Y��jC!5ң������N��P1a����0/%$��������֎�l�甠�(0򥰋�X~	�`d�6�* ��n���_���UJ�dRS�{�n�2c�2r�Q�0�m"unPr! V���&�oZ�mh�Qg�֎InB5���`i?|���t�#�S��=x���Cӳ8e,"UE�<��x����ɛ58�޻"zjdb��m�S��ݥ�GI�u'�!g�*f^M}9���Of��o����|ٰ].��W�{�qO�.IƬb�q��d�X��3Ns|��{V
1"�|��q�W�#�kg��,m�hT2s���Q����r�GD�H�粒��[%{���mlR2��wK�Ql]$QsZ'��	*����.9=����^�<�#}4���P�ɮ/��
�Q
Wk=���V�>�?��ũ"��������+R���ЎN��OW_�L
�
��=w�����m�m
	�;�c�H�YF��wr��⬐W�;Hڜe�а��L	[[���������t�9�lK`�?���Ѕh���'B�l6�$-D_��$!� wq�$��pКF�ŝFf �j��j�E����Rz@���NJ�/���tD�t�_4��B��gFm�VP��=9�UP;Pk�M��kԓ�uƗ�}�����?~����p}��=���"6~� �����%!ӆ�������_��+Ralϟ�~��k��59��q)c+��;v��y���~�z��@�>�G�A:�<G�	ˢ|�Xc���G]<%6Mq�!'����>���x�c�{�j�20[�[���)[��!Q���& �p޸�U����Z|'�ӴI�,(%��C����T���n�òH���%  �¦�6'���vTS���.tS1������tl0�8�h��~0�G��ē�~�	�l��s�.���n2�MƲ�b���4Xsw@�O�r���p������`�B��#��tf�a�TU�����C/ <�[�b-.�*���������cs�`v�}���}�֛�k	�(Pjf�mD���H��QG��A��P�H��&rR������U���:"^{�1_7pD�0o�G�?F�M'��b�/�#"Pɰ�C�L�{vܳ�l�M���KWψ;��#Yo�X��&>t4]�?#�A:��%�X�~ԄR.#z#��0N�d����
��i��"�D� �7�'�!"U�3�S �
��rV�^ ��	��=�T4D����{Jfs_�h��4	�W��M�����e�N!�4A����tM(�e�٧���a�2�w���Q["�۽/��X@t�S`����v�5d��;���\	�}%Tj��u��%� V����S��s��R=���t�=�{GZ�$|w-�ׯ������u�������G��������5{I�m���`�	�M�	9[�����/���ϟL`��$ŻK�gs<,MN�z��A[����L~~�th���=��e� �X܃��8��qI���v�B���M����КX{�����g�(϶`/��`�QMHLE1S�38w?��o��[�G���¸n	�-��-Q�+��|�ã�Y�b JJ['�~1T��M~J�����(*�>�4Q�l W�ƈ]�������<�D�����H,~�@�����q1� H���1���@OV��<��LАMUjkh2�L�+�}��W�8yJ#j��K���'���eÿ�"�c�H+���Hv�����E��wD� �!0�-N(T����Q���tk(��(g|�� �͌��9D@�G�    IDAT����q�;%1T�WTj@�Z�y���Z���ώ��$M��~��p���֞�*�_���Y������ޛ�o��*�0f� 	RA�� �35Xnw˭������#��n�����%Q��E�4e�@ A��\�B�oμ���?�so���DTTፙ'��g��Z����%d�����f���++E�<��@���e��ΙJ�N	��x�(�-����H��b��(�D<�"�C11���si"����$o���=�U�7��RbYK�w(�l��#�8Ė��ere��5�������-I1Ns�=��qU�F!�7�Ij�#뙒/���_I���z����~Q�Ȯ���g�����9G׉ki][����k������X��F8:C��.��|�b�$v���j��ҩS�Nˌ� ��)$NNjC��W�`�4�oٔ���� @*3��d�Jb	�Q0�E��Ya��=��񐉃��TN���IeB�O�d��M��y�%�%7O����xsE?|�U)�^�_��,D{���Ɛ����9�@/���\x!f)�r.��cL�Q�s2k{�'��G��k�`�}d�{Z���*���I䌳���j7���*��J,		J��i%L�`�H��2/�D�c��Rb�9I%����5���MJy�k��R.mY��Y	���ȧ��Ju@?V�h���@�$�2�aб�7A?eY�5��M9c�*ci˔+�����]	��\���e�ð�Fȕ:er�D%)��W��"�*r����5r�����VT���v%Q\MІ�D9��=���4�H���"Hv�u�ʾ�=!�T�2d�ҧA�h�p�4gxV���uA��_�V��yK]�����]��}+Iu�H����L-���șZ��-���?�\����+}�qK#�
�Q����	��(W���Ң�����,�򸏼/�v�fRa�jm�@���.�&���Ƣ�Њd��^���*M��d�T�2�����o\���9$��A��9�2vs��n�.�T�ͪ�x(�w�c�Ab(D�jo��@���S�^�w�������[�G�z�cK��j��"��ȹ��=��f
��fA�Ȟ�GT�9b�xϨ$�&i�*���e,m?[#�ؗ�01���<<T�x��H9�"g#�v�$��ϱS���:���]���b�jl������Ry��AQF�u��q�6�Ƅ��A�N�\�
U��9��9�����!E]�I0�ދ������:�q����~z����S	�Y���Z�Q#��Qi%z�<f�r�+k�V�Au��� ����!����s8�	�b�z�P��q��L,��X-=�a����(pD�5o��U	j�3��a_]�d2�J%����`(�F�e�voP��#X����u7��q�k�[>��ɱ�~���Ҕ�RnF]d�F��L��i �!���ɒs�hg%����s$dI�T��	��^�	��ԋ#b�!�:Qa(�$�i�ƩY�@6KxsHb��I&,�e�� J�D�ܽ��)��\R�$=��8�E�{�x�4���;�Y&BZe���,�W�+Axx���P�$ic��)1F�V����YUܳ"k�Eo�AO�@[*��NK�_E�R��ɑ�[c.ܙA�b��K�	�f6�-}顂���Ј�Tͱ׿���8$��JK7%���;���K^Id(m�j|�$����-4a��&hBIb2g�*��p����9���P1��ҚL)��K�*��.B҈��P�etц��a!$ű��h]�,�H��jxoƌ� �f8�Y���D�0F\=��#�	�):��R�"q�j��S�mK��
AȆ�TP8(r.�EjJ�"NY�
eN��c!�j��	~Qΐ�:[.�}���LLU҆0)(]Kԑz}����=*����ȽQ���r)Y��'��Ѱ6�h;M�R�*m�1qx8'z���W�,�S�|B�٣�������6_n�(w�$��J~�[��%2|o�I�p	�T��b ��
�Y�3B.+a �iip��@����R��D�F��-~ޞ\�'uU	�Bi�����1ȥTY��m�p�	^�i�{S�)���)�l�M5��F�y�QG�jhdH{����\�:\d�(����*"Y��TW��qEv��Y�9f��r,y%��a�[Y���Ѓ-`�@�I���<��d�+�����SGf
�F���/�䘢����*�3YI`WrX2k硣q�h�c¤�5�"���F%�DiP�#1&��*�i��d�)��,?g��VL���@z)�d��>�ՊE�cQ��`�Nk��ֲ�]𘪆����S�!'|�0N�![Ȇ6w����P�PAz���$����"�6���>�HtN���7�*J^��A������I3S5��a����(dWg,:+RL8���E��⍭ѵ�hs��iTJ�{�F��T�(�&��GbH�TV䏊�"U!�TAI`����%{�<u�D�Ӓ�1٠�.L� ɷI(-��dxN
��8Q9�xmK�>}^��S��N���P�8^�a�&'�DL��G�����l�o��]���YK;�IJ���2��g�$�iI�M��K�ܡHڢ��ԩ��J��1N�m��3���1�
K�%�I.zce�b,4mI��� �t�R�B
���LLF����Z�X;Gi�h-}���&��YE-S�]*Ð�i���Z&I^w�jAnb�,�sы'd��jLt��F�@� �۞*��e���wDև��PV��i�O���p�{�����n:u�X\����*1�-��a�yْp�A��C6�d5�]P���Y�!֐z! V��$����j�pDB�+{�8��1�l��8�Q�'@I���"y�r����m��b�=,����>����I5��E�Xs��a��.=��Ά��@!j���JĤ�}�-Cob)tU����dg���稲0���jP�%�e�����-�2��3�ɥ�Υ�Py�ͬ����죫�[�j��1Xw8�P*���J
��2�	}��UHYL���Z6g�^�g�$0�a��rAyO�����laŖD"��i��c���Tr��i�l�D��(����eA?t�Ţ��f|�F�XG�V*cH	B��s5�L��zR��
)�i�5���/<'6Nsxx�I�3��[*�)�&*m0��͑�"n�r�[�q��:E�z&MC�,��9B�1g��:қ:�BB{�tNdjWs"F���]���|$j�:F�2$�`+A<���곐��PY3�,3]Ѧ��T ZS7		�Yn.Z�U`ZA�ʲ�=�d�,	����.���zzd��*[��%`��G�s���ڢ���~��΂�D	JF+�0Q���Y����@Ohm�j*�6��(}ie��i���b{�3��6�U��eV9�L�C��Jҥ��Ŵ.���S��H�K���(_�A"8�2o��@��\QJߎ�V��-��8&�S;�w�0�]Ɵ1)=g
�\��L�Lf��q�G�:]8��AR�=�d#�<�Y�|L!�*�l��<�c�fA�ք�`6�uA8�b�QH2s�T�B�D1�q�,S�Xt��	�(e͍�;(�9uz��j��gZUԕe_�24%�1��֎�������L�
�,9Gv��\����N��~����D5$ʜ(�d�pJbf1�	Q��i�i�tpi-��g��mm.NhÛ;�"n����Z�����2�L�#��K/0�ю{94�en���J�*�_��0�� ��e�Gq�*>�0e����q��RY�N�@IIHXՑ�K�?+m*re	!� +ĭ#�2(WC�K�~��]������,�{��}��<�6o=��9X��+!��oXl�s�%[!�iB�mЌ�G'�����E.'=*����,�n|=ZK�u�u�A��L�+?hx}
�Q$���H��{b��P���_�"�]B�	>���)��)b襟����zʹ��!�$]��	�j�޵���&��^ ��`�Hw�SO�D��-�G*�p(*}e��4_�%$	:�����F�$�:c+�.Ěd�B�] $/h�#mچ.J�`G,]�醘h��m',줒�+A�Z��iO� ��s�O�]��AA�b��!�H���vt}�s#��g;��C,գHR�2����++����*T��l7Ɗ�%
��\��Qs�} ��YN�q���%�q�I�=�I�ƪ��\���0��pPC���3�u&e)8bX��r+���F��}����l5�S��Zk��۟����@��E��2,�5�^�]fpO9���K�@����27^~�� %�TB+�yzx��:��g�Ť�R� �t\������l�rZ�QZ�2�:ĕ�^�:�U����E=|L^�Z)��6��隐"��SUM�ɩB���`Q8�kWn�S��֌��M��}B��f5:Ɉiqf4�3h��*�,8�ޓ�e�c��F-��fss"�LJ�$i��s��"�T(9kr�1�L�h����#�5˻euM(�(�\\y����hc��F�����pІ9K*Fbg+A_zE:�q�)�)��*��ˍ:�ڇ�/��\�]߳�C2!,���7	�d�N]i��8/����k�4Ρ�!$�<��~�=6z�F\���@r&�Rqr�辕+���@�&g�@��-a&Y��v���PW�`U򨦙�m�&�	J[�N��u5���G�gmdʞ���x�)
�8�1��8G��E�&ɖx&�uuU��y�K�Qz�37�$˚�(������MQ�eIHjm���!3�s��O�IE���8��>���
׈�ݼ�HYa�
���)��g��(e����꘭M�bb>?B�$�A�̰�õ���p�[�"���>2k6�8�ӊ.{b�Ljl/���
�=�H2���<Ejנ�@�*�a��{�ʠtE��[�4��0&|��$���h�9�(�X�HJ$)VF��h����'����u��*�!2	GC�BP�.F��ւ�h$8�{��:�2KR���".��T"r)h��8�����^z��J���D�0�E�Q�)J�L����yKNYZC��a�,�>�9��z�qHj����Y�>�c�+c1	���Z�@&EAܪ��>T�G�$n�Xi�(%��z��X�q��=�]�R"9�+D�,kd�Y��'���^���T���
�V>�!�&1Y����h1�,���-c\&�޲��h���%�T�#��"K�m�c�X'�R��t�.Vq�x��j���<�Q�T��9&���2kJR�9J��g*�y��+7�����&}��`~�lcJ���:EP�Ȝ�EY[�7�T�g�h�}�R���"\��O�l�LfT�r��O�=�3e�\�H�b/?H�T��iuݤ�A�� 'Q�x�9S�c*6��)�.�2Xu_+�x�d4o~Ĕ�!���V.��ʳ�PYq�S��?0����Hde�Y���ۀ��&���<�,��Jklm�j[�+,�e*�Tj�fJ�����yϢM�w���t*�Y�X�_�����WMntF�6G��
��0��м2��u�47��]�z�i�(��dڊ��4MK�~|���+,ڀs	�K\Q��sɑ�GR��.3�&�1���!�Z)*�n��D$I�Q��LT��2M�N,6��&0��'�&'��-1���`�[V���f2�d��1��
U�:��ts�ߜ�K�k��4�&��o[��'�ln�I+�T��vi��Y�ƹ[n�M����۞M�Z��	&�)&f�B4}�$����Cb3���GsrJl�X��Pƞ�v���uE�p��������N�>��.Y�%��r�jp�Js�=�4���~A���k���o�`'uaF;�^��ڊi�������dĩ��={�P�ơkCT�Eb`��:�D!��"_j����"tR%ZC"�A�B�Vӻ
��,�!0�I?#�L���Ge�I�k�@1ʢ��1Y��q��E��9�3��H��� �-Ҧ��9[TR��_ι$�r㌭	[W(BNYZ~9/��>-��K��%28�D�q�������~ �^v:v�k`���v��~�����|�mE�̊N��CI�
�W�i�]����T�I'ȕ\�c�8ĶRh2�^٠$ ���-�՜W�F%�ə���Ue�T5ދ߂Q����S'�qLfR|KH�J�]�l2�Ϟk�n`9���غb�pe�g�3��5��й�jI�
��ZGD�Л�lolP[��jFjgI�F�CAŴ�2 ��f�` q�{5�Y����a�/̅ݧe���f���^L�fơ!��m�̌�F�c ���
�O�@��N�9K
Yz`9���"Ӷ��7��#�J8�d�����ZAAHe-:[��/z�">$���)�g��Cb~�`~�-3�Ĩ2�h�`�mJ�RU'bX�W�	SPK2��V�ח�B��.��a΄4@w+��4���"��9�e�1��q���� �#C��V��B�Qe�]�n�r �Pt���4���=�k$E_�u��-�QPk��8eXsR���#��*Ƅ3�T��ӷ���Eߓ+K3m�)�|`�5��@<�Ռ���˾���`v�,=���K8���2�uSr�Z���a�AEΎ�F�ͫ���mS3�pp���)�ٔ8kH���&��h�F������H4��ֈ�Ȯ��ɔ�Ye&�|A�.Xs���k��ޠ�7�.�X�i���t6����� k]�`�6'k��U���d���6�����T�#���!����2�\�$#�`�W����1���!K�=�=g�ħ��Z3�08SIB%!���ʚ�����V�W����,�������κh�k!4� -��\(%��2�e������J��#h�I�=vR肶h���x�}�Z���4gq΃"5-��#){���!���P1+��vz99r��1J�g�j����Z򕆷�V2!T�Y�V+���"UČ��`BAw�R��r��I�8H����0@�C[v�������)��%�:�qU���c�dF��>D���\�T�_����X�+��k5m9��դ���h���՛��Y�7O�+C7�IeN!,A)��%��۴�8c9�<]{H����h{n�=�MŤ24�	��	��䈮�"��T!,k�ǹ0yl�jr�; �c���氲A�a(�/#�S���7k+e�5)�6H����]yon��j���B�JJ,C�
6C�˨ٶ̈́\�t(AJE��"��$(e�>�"�(},�DTRx�Yt��6���0���R
8%�R��Qo��W�J�ó
y��i���������.���1�*�M��J��p��{��-3@熬/@F��c����i�<W5؏&9H����#���l�=��?9k���9JGX��(�G�>[�֠�����G�
j�YK0��.�z�b���v!6�1���ٴ������{4�[�z�N+���8�^���-���l��³3�x��>ŝ�}/�j�?��=�].��I�y��;`������_��C�R7kh���e^����������r�ּ��1����n9C{x���'�˫�>�y������d����9GJ'�}�	��^fۛ��\�e^��wY\��&�^��[�������3?�}�"�e�y�[Ǿ��b�>���s?��9�k\z�2��/���+ldM�u��!Lj���Fۊ:�)�aV�a�9ʙX9���!01�Y-R�6��8��wc��s�iÚ�h����<F;��x4��HCơ�*�v��*c�C ��9�L�5"+~�.��Q=���\N�1@֠E�)�����*-U@�TV��{d���5��E�ŭ."oeRA7��A�E�Ҕ���H��z���C}1�)2�Q���k�IA�2z5���n�_>Hㄸ�����e%hj�Ę*J�+�����K'���g
O*%�72�+�*!,EN��5�_��"Y__�6�)I�UZ�H�mo~�o�f~����M��&',�5!fQ|�J�Zi�ʒQt����Y����/_c��&ӵMZ��HE�,��jhk+�3ð�^fH��/"��ɳ�Ym%q��!��50ʎ�$Q�?�"rH"����l�x�%F�����7�m*,�qqWu���|�2�1�Vn@[p�z��     IDATଘ���6���{��,�e�=�6�{�65Y��ٖ�hT�n,��ᜥ+��R�rN�8�e4�4}�8j{��21�~����we�i,�T$���ҫ�Ky�ƌ�;s����� k��ZO�b��G��<^��v�T�*�!��Fӕʊ���^���a��禜�aQ����X2�㩉*WB�D�JKBB�(��S_*��r1�����d��*˦��c��c?f�j����O|�殻�M�;�0W�s�k�`���qz}5���&���N�Wg��2��4n���<�7�^C���9s����>��'���W^�|�W_��~]��눽�N�����U��6:+v/\�c��~v�{������=�m�?�#_��>�~�����H���~��������+׸�����4�|�#����������������(g��S�ж-n{�{{w}�K���,vsFUk��>?��,O�ٟr�W9m[g���/�����ޜ�^|���Xw{)b��<��'�����ؓg�?�c�������^z��[O}�$k��f��yt�p�S�l��������O��ݣr?i��&�m�.^�?��ێv�9�Ʈ�ѬO9T���5��e~pH����11IU����Ja�60V$Q9x��z*�;G�#� .@ѿI�`��$cTS[kce�h��H� �G�5�D�^�Q��Zx}���(*�&E��Xt=��(�H�2�������n�s$����Ȥ�@ʕ�J'r�a)���=���ἧ�8h��o���'���+�ᒔ��3�Wk��d�(�;�{�E��Ȝ���^x�\~W��*ÀR����Qf9gp4�1�����V7�,��XGU�+j�Tc�0@g9b�Th���ؘM�8}�����>)D�6��z1l2���S��̦5��c��7�a����Ţ���[�>q���ڣ#j%fl¼T�h%{�6O�
m�iC�2k@"����*W4��T�2��D�o���8��	�X�/?�J[ehK{��� �:fB��WK�WIzLZ)��M�/(r��Z�Ԯ�{����D'��/�TMS�5�2��d�]��ؑTBP����|�w��@;Hi��n}�S;�lRaj��d�І�BU�X�-��`����Q+z|�$�I�}�6f�x��C�*2i49�K��У*ɏN�)�h٥�&0I�*r�%�q�
#~��Qe��1z�e���c�R�v���J�P!D��$��8�bMqk*�G)��y��	��r؄F�d�+O��:ҕ��=�T�z��ҵl��<�?����9C�����)w<}�y���?`著�=���ſ����iU�w7�ؚ�#�����C����k���O��~�jcK�*>�x������������ g�|���w��S����O�N�վa��q���n�s��ѳ-~���py��� r��f�>�={�Ǿ�.��qt�=�y6��(�_z���_�ԩӬ����x��z�������OXo���ɩ#LZҽ��¯�/�q�n^e~�2}��4���A�7�����W��'>��<��������Ѥ.�hNq�]��;>�[�Zw�������y�_�ǿ���N��_彏}�����y�V�t:E��>�������Wh����r?�����<�/��7|���-�{�����0rE5���/���/鋸8a�n�Y�ܳ�����X{�
�eK�m��5�}❟�,���J��0ϥ�7���7�ug�Nk�p�{>��O?�l}�~����n��3^���p��9�j~|��>���YO~�����f��R@�6W�6���ȭ��g�&;��v�v�e��_c�{�E7[�z��S��q��â_���S?��]�o4\ٿ��n���G؊��kv�`��s��	B?e�G�g��� Ѩb�]n�	#�]K� f`��@�z0^�Is�{"#v�>9g|7k���W/ڷ!���ּYY%?/��"-�֍AlEʚ.dj�i4F��I���p�e8$19ʰ���bņ{�*�l���AZH�)Z�|��f���>���6�����1�
3]��KR��"F�Ɂ�Z��.��ZZ�֠7�� �Slo���ឨz�H����Z̼�{�5L�
���ӶN�>F;�89mF�$@G�*f�J�Z;����9Cb!"k��Q+q\�$���)����E���2K��X͗�������x��j�suɲJO����h�V��t�3Z��L���	1ѵ��zOR1c��9�VL��I�+-��x)��Ӣ'���6�M�|H�)rW�����B<Js�5�d��r8V�������B&FGJp$��稵f�eX�l�$,�T����׏�@1)	iU�ddE��qP7�J��]���������������ս�٘������w�/�:�.�ŋ�=�ͯ��3��wr��>��m��K�'w?�0w��Q�þ���J�:Au�=l�y������p�:�m����������ₓ'α}��}�q��_���\{���ml�{isµ~�S��|�96���}�]���&��2v���ғ�������?¶��W<���	�}�W`�ŝ�?���.w}���r�"������g�C�?���;�#Ln=���6�JI�}"�}�<���7��?������E�����[��?�x�������Oos���hgIܹf�yl�y�'T���w}��4�-���п�
a_��������'>ƅ�a�%z��l�;�����]~��8����4O|��|��_������<���Μ�p���)j�BŊ�l���>�c_�5�ٜ�'o��	{�-��<�;{�f�x�������T�浝=���'��o���n�7۞~�q˹[��y�O��4�x�W~�G�k︇S[�\������2�V>��_~�x�Q��?����.q��3����(v�Z��^]f���㷹�}�&�L�3S�y��g����0���h�{��}�㗸�����{��}&���k?���O��ty������'��s�g���f��l�q����C��W��Sf��0f@�2Bz.@k�۞����/��%���z���1���!�UH�{A@sc܈((�Dm�	
�T���8���RXS�?��20h`�(����#A�Ǟ��A6��9� ,��A+�����v�9o��y���X��2�F-����9����*1�)�G�2���@�/��;w���:}���Pi�t:���t�B�N9�G�X��8:���깪"��������&T͔~�
�^+|AG\U��Od/[���#&sL,\�7u5Ɗ~x#J��f�j쭶�)F����^.�߆X���IIU%�\r��`Tq�+>�F�1�3�7�}�me�m�r	̔I�Tuʹ��+a$'�8P��d���b(6��`�1�Gay��眄)Y;f�H¬Vh#�C�����&�6���+LZ%�����2�v	�����/��(NhC�5)I߭�/룸��2h���8zd�co�� ��+�A��׼�VoV�N�5����kx��'ư��[γy��tNsp�?�����W�n�A��u����� �[l{��g���^ϓ������u�N���������lms���\{�"��/��+����9���<{/�~��������;9}���t�2'�	��	t�0�V4G;lܼJn�x��_��o}{c�I�G�������ĠiXu��[y��e.��0]K\?<��]w��Q���K/s��U�\���}���8GU�Ʊ�JYL]�]���w����^������0�
�}Y��f�/=Kz��ŝ���}�)��Y��cq�2���܅;�c��^z��=�t�]�'��X���<��ٻ�`��5��_�/}�[�Վ���s�|��oq��)n{�!rS�XAH�Um�^k��� �������y��'_�
���S6N���2��?��'~���~���78�<�<�(���/1��vvo�Ć�+���v�{~�O��?�������Я~��|�K�/b�w������!��u'���܌K���W����5���}�Ҧ����S
�>D��w��|��?�k*v~�2��4����G>�Gw�����A�j>��g��N�5�"z�>��gxn�g���'��=����6�ﻗ���#'N���S�c�ow�5��x��Β��,�Y���^
�6�Q��J�]���]��c�RǾw��cQT1_�M:"���B4�C����C��&�J�
rz%b�#ypPr)%�+�JP̡�P*R17%�q_�b�%� #n��y�k�^��[O�6���}K�rkP	�0��E�����8��4zJh��ve�|z���'QJ1�ۧ�QEq,��Xm�
��2�����c�%g��|�(��r��E߯WTK*��i�
+ne�xl$�����!}���I�h���Y�Il)%�/������/= W�����:bH��t�G�0��ã^��A�U�Rt�fb�M*�J��~@ ��b�S�~�2�lh�@�fI�"WN��Sh�65�IMe�}+H^t��C�2�?~�
�����e����,g��68j��膍8F��Z����H�3�e�Ġ�l�t��N {y��ؔO;���������0f��8H�A����m�'��8��6��1s{p�N��޸�w�Ϳ��S����%f��~�c���7������:�5�G�̻}n�	}����U^��7���bqu�L�t�)���p�/��S�'��r4.�U��Q��U5a�4�՜�4��c�s��l���6�����qb�);�S���Or��>D}j�+��/=�c��»1ʲ�>c}�!��������т��#eKek�6�.��C����mm&���@=es3p�[�7�M��`� �_|��]wS���ȡ���2��/?��g���p?�������ǆ���}�p��wC=ag� ;��6��L޻I�z��2?�^����xe����Por��1=y��SSf�O���8p���n����l���&�lϘ��8�x��~�=6���w�No;Bw@�����}�;��Nnܸ�s��?��W^c�[q���<p���u��W�ek��W~�w��G��^���L���?��y���}�[�=|�s�����U�EO��Dc�Y�miN*�.���cV+���7��_}��y`��{y��>���� ���-^}�w\�����<�wNz�u�AOw�9ο�ݜ���?�0;����?ȉS���w�/����	7x�s�x�<�^��k<������W�\3��Փ4�,��\Y/��۟ͷ;�ow鏿{%f-�D
0*�+-

(V�����M���Nȸ�]�]�0zH�Ń ��4�di?�2�	,�O^�v@�c�Ru���$��H(��s�Ir}���Mn=���t��L�%��Y��|)�,�g4j*E�|��M�lbg�s���9���	���-��RkKO�	�k���O]�Q�|�Ĭ0vJ֙�E�W�[��8:أ��X��`��T��T�V��eT�T���Շ5�(��#��6ƱgH>��>F�V���:aM6MEU[������$px(��C����,:]z5j9w=G,��f2�����������w�y���Bf>o�;Fs;Ȃr��DS[f��YUl?���.d�����[�V���N��!��?�o�Y�v�2�Ojb�8���e��Le�ϴ)J\BI҆��#gF�~�"�+����ҁj�up<��b2�6jPTȘY�*|���w�N@c];�G1ٞ��W��)��gNlspc��+�4vJ���['x�3���;�2���5�Wa�*}��Ln� 7��=����g8ur��~ʥ�_ �hei}�J�%�J�c:�������2lO�i��*�����~��[���3��G��ثװ�CE`��͏8�-���}��l�3��Z�*HZ�����P�s���^z5�����{g��/����~�Z�D	��*E��˯<�O��m�w�A>��g�:֫)zn�d�p���looR'E���3�ºs�����<C����3������!�x�cd9�T�ӧ9q�}�{�mx���/��4g��]_�"��;y��6�>�։m��_�۽�Վ�+&�T�5^�9?��W�^�9�̯��S��e~�������ȳ�ٹq��g���Ϲy����ǰ�3�6gp��E����dr�^�/�#qlt��8w�}�A�{6�i���2���?d��"�)��}N�o�s߃0��R{\z�ܸ�S.}�����P�μ���_�v�>-�jA�����}����?`q�i^�����e>\Mx��'x��x�k�uc[�/��{#��3��~��/"�cj��E�@�[��Qn���c��3F-.�*�C��e{]�N�ur���5&��������Rp���KH���\|BB��H2sbq��8ƛ!v#yS�hS���e�r�{Az�Nkn��k봋׮g�uM�:bޖL�Ћb?��؃O��-�DH�E�\͢;�׮r��&�Mt=e�&Z	�<��̙,�]��Ȋ���.II_�������u����D�2(�R�p%a��	J��7_�ח� .�hC��Z/�h��J���v�D,��q��t�1���[ ���-�m�98��z
y`�Kժvm����¦M��a�T��4��4����-9�Pi�hS��$�ڰ6�ehM쎙����&��ck3.����}�8Ō�
K���h�ٹF�(5ZM��fIZ�*���ب)�AI$��x�����5E^���ˡ�{���[���[�vx� !q��������4kL�#�[��WMH��!������g��]�3q�j�Ƒ6��x���>�9&�f����+~��L�&lmv�ܟ�7;ǝ������y?���������{�v���6�4��!�9:vl�m��ȼح��+M�n�p�'?��O|���S�7�`��|��o��M*�V��9��3QS��r�R�W���g�j,����Me"W����H�����U;6�<��3;/^�9�B�l�l����K��G�}��67*M[5�p�|�eۜ_�96��e֔äHT���b֧�����דd�y����1��u�o��	K�Z��(�Ԉ�fF�������^�^n�^�_�&&b6bcCژI�D/�I�
$Cx�э������NfU7�ܘ�MDG���N�9�3�����<d2��ң�wo��2o�Hi8u��;����a���E���q���(��y�Ǩl�7(Q�a륟"����B�O��ǻ��+eK��j]3��3��f\����k��XN*�<�G�~���1�Yר_��_���O|���s7kGNp)/�ن2+�JSAA�$�ر?����ð�Y[r��u^�OK�}�."�����Qm_d�U�R�Z�]��0�O�MTs�d�^��?�������;��'N�������S�N�*K4m�[��u*B�~Ym}�Z$�2�ņz8(8��M�^��%���ɔ}/J!�RċHT�� ��戲�̧�L��x�24}�˲,@�Sp�����`�@�N2�~�%Ow�a�hh;�����01.�<1��6��y�'2���L2�!���AD�2&%">!J�4�E�(à��ڈ.�#)I�x���Ǩu�׆��3��B��I���:)b�p!i/���Y�hmC$u%ضek{�c'��z�8{7��V3����W��m;?��:1#�A+�-M�������m�:AW�H����b��5B&("��c����)hm2��k��*��u��R$�z�ѣ��@�����:F�ka�x�5����b�e�΂H�|��BR"�$P jRݨݠ�N-'�ቹ����@�xW2�X�5D��N�)��}����=S��2!��pGt	� �_�r�ʎp�N��V� �[�����K6�_����u����~����7�M�\#K���6��͈IS3�0�"�9E��W%7&5[k=�����o�.������/��~��9GQ�X�pa��cO�������ٻr�����s��C�J�K7E�@	l�״1c�r\e���9v�}��=�7��+�UN}��|����ͣ윿�O���\}�_Ѻ������\�d�Ĭ��~�\+����ꏿG}�<*�o�)3C/S��)�%�    IDAT��Uv�}��}�ɹ���8��l�*囖#f@�*��vV�\ ��	2玻��>�U��|�4W/sdx���S���cl_��{���H]WT�);;;�֒�
jgP����
E���錙ќߺL[(��S^��yn{�z?�x��[��;X�\?��9u����a>����1B��i�����ٜ�Q>bV��"8��F��?����|��tɻ��#��>�訂gP�X=}�<�A�y�;�/_�H���r� �{��gSJS�"Զfg�K�4�8�lf�Lc�7}��R��3�#g������(�7��.~���B5e(3��~������c�\r��y�����e��J��Z����.��ͼ��'�5����T�;��ە�k�-��.�;���z<'��}����B�����}�,ce8�5-�;�E~)�ە���p�[x�,aɖ�²ĸDM�l|��+y�@�-k���ܳ�?'I�� �E�DB�LC[M����򵌝iW�F(�E�ܪZO����BPf6�l��EhA4º)��������5Pj�I
^�@Y&Ѳi�Ҷ"M5o�ٛ�2C9\EI�uU2t��im�1.;����^'h�����f	�gq���2E*>�TI_�3� ��Ki6���%F|T՜ɬaȲm;?�Qˤv����6޳�8L2IpQr��ז�������|gɈx�5�,Ɍ xK��"���V���$��'�AT�%���6T�B�39tJ�0��t��^�պd>C��4:��]�WFỚ��R�A�Y�.�Ӂ�Bt��� =qK�p���b��0������{���E;�~o�2������! +Olי�d<�r�ͷ���E�;�v�G>�;<����_2�x�7��%���_r&dȨ6���я�����g���w/�ӿ�[^���8�$�l�����{�i@�s�^��LkN|�I>������g��z��>�1>����ޑ�.^��~��^�)�j�scn�ݛ�7�����3�C^X;r����X-�E����%�s�Q ��|�W�W��;l��)F�����x������.�.�'&�5��&r�4�R[�0SLww9"r�?s|��q͍W�������V�X=�����	3g��F��B��M�d
���h��3���4�<f�&n�ǭ8.�r}%c���a4ൟ}���e����������;�k%���fG@��l0����O��O=�D�L\�Ɛ��628~����?c��ӬyŹo|�_|���{�U�Wf{3z�����Nb���nl'�ƒG����1�Nq�3��R̥C���Y`��pUdhrz�ǎ��18�ß�S���X[Y���>�[�U�;7X=����j���+o1��,�T)8���{d1�C��T:�p��"Yf�˵�vs.�n��o������`��Yܽ����]��7c�_����T�3hj��-%���A9Uk�4j��K)p~��Jv�A��o%S�(�,�Ӊ9�*�Z����u��	Q�X��d&g}m�d��6^H�Ҍ����"ǶslӢ"I,Iij�L�xv�%P:#˓��t�R�%v�bH���g\���Qs�����7mP�Ӧ���{��D���єf3KU�7�^���M�V�y�	�&�e9$�S�~\�&>����?t�<�|!���C�۷�	@�1Q|H.tZw&2��P-74�H�ؕ2&����N� �&i]�P��p�()��W��t� ��q�E�㜣u	RiI5o����j��RG�4�݌�0E�VI�2�Ā�>b[(�N�Z�O=��mZd7��1H!��u���L'}Ҹ^ԧ�k?��$;U�Ұ\��(���[W�	�hA�
'"�ZA�`f��!m�"�������@�䒬He�� ���9�7C8���e�qA�\�OZd�`��� � 6`t�!������|����|���}�3��3�����	����x�>NcV��{����_��s?dqm@5o�r@��Gx賿ý���ƅ7��_�5��=�}�S��
�+(����!�N����{����3�_����u�(4�ʇ�C������Y&9���8s�Ѱǻo�����Cx�'�O?���ɿ���;��_�p幟v�Հ�A�5j"�����1*�)�����}���w�i��g���<���r��D錓~
1��=�w��w�s���y�����_���=I��W�q�!|�d~ieŉu��#�y�)^����׮`O�e�c�p��q�/0��A�	��2[�ݺ���Y�>�R5�U>����uvϿ������;o]�诒ݤ8�ct�O��{!G�/�1����;�1~�:���h��ezҒ�	�e{"�ￗ������&����������9��g2���ML�g�d�j~���Kh2�8%�uͺR�9�j�KJ�v\
jE�#{�ǂ����i>�����������o|�k�a�6�5����0�����L^�f��Ӝ��Gat7����k�_:�	���X���l^,��˵bcs��pSV������Þ"]ORB�Ę-PĐ�ޣ� T�䬭�`-v��2�b����%F��H������@p.I#��բER���#c�]�wF:Gͮ���
GV���P�Q�A�A�֢��Zk�M�
A�[q��ʉ�GX;z���v>�(�u�	�x��$>@�`�y�U;�IE49Aj4���޾���,�J+����`C�+p
g#���z, 4dRs�����C)� /��ʹ+��L	lt��I�k�j�,6��;���5�D:EO���ypܺ�� ��H��Lm�5�E���4>t��ݐ�!`�$W9Z��:�W�6 O�"�e�Y���jh�K��*�tJ@�iz2i���,v�������]})q�Tx�P�@�=���;�n�y�o�:�1]m閶��"���"��J)l̓U�NѠk�#��`�"&��(�C�Ut�7��B
���?~�=�/}$��������
T�tw��7��3�s�SO�3����rG�('?�Iځd����'��x���	�V����\����󱏡�Ǳ�����^����<�?�kN<p[x�����Cw>�@¥�os����&�ɔW��m�p���ڧ�8}7a��\�8ݗL�|�W��#����O��z8�9�#h��ǎ#T��9{�1������S��=}�>�����3��u~�����~L�ִ�E��2/(2���[���*g����z?/�\f.��Ư���R�}��y���G���N5Z���G����=|��?��ƻ�틼�����Ü���E�S���9�so����G�z����E~�4�?�4�hح���#�'�c8��b�E.�q���Rek�j����|5�}�x��j��eǑ+s���_z�^���ǟ���1ۺ�؃�)`��1�n�8}�~�3<�=����9r�,��������?���+�'x�c����?���}�~���@�U��
� �&gV\#��,ֵ�K&�#�k�:x��5eV��k�Ռ�ǟ��s�l���N��(��n�v���o?Kq|��>��<���f�?�Ͼ�U��Ɨ�7�����8Ǖ���yUl2ۺBo2��_�"��*�=��ާǜ=��͓L޹�0������k���?~�M���9�!���D���d��Z�Cn4���|b�w�wr]���.%�}�� �:ą��b]J|��~!E�K?� ��v`�[�֦�-Q��EP:yH����ltc�9���%��K�,'��?\c��tF�g��g��β�yc\�e��@�6�q��9��+��JV%���{;�&��{�nj�0�D�H�i�,co:���8��,^G�N��[co���rz-;���nW�}������>�W�����z���q��Ԉ�;=�j�A��
�IJwBdg�(��EO m�.¬n��
�I.."XB2�)3CiR���ӻ����H�̓b�R��>N�ŀ�졵X/�kC�(y�t�̒}��/�XE.n&�F�sԺǩG�g�\��N��6�<����Ow���e�$�ɂ_�P�pHR�ts���&��޿x�&��n,"[W�g�z���{z�p߇�౧��ޏ|��n�~&P�m^��W����x���1���?���G2�s��W����c�s�c����n��w���am��4wU3~�9^��78���x�����.�?���m�i�����R��&�������or����L��eF6,A�4[W�Wށ틼���"L��a�ƩS(�ع�åg���_�*��-D&�yF1��)7�݋\���Y�n>p�(�GE�}y�aV�^�����k�Ǐ�#,>2	1/Y[[a����d����͓<�G��V�Bè'�v�M^�������'[]'��Ͻ~�{����cLWK���e���y�0�������;���I>��Ğ.x�{_�]����~��^Q�y�4�=���:G��u�2o���4�;de��l��� ���q����w�,�޸���q����ńW��	��I��o���$�J��kW�����W2|����W޼�y��}w��T�U�y����W���2�����HE�rFN���������T�>+�Gy��ft4����=��]��دq����\�t��׮0��!��u�z���E��O|
�������f���ѣȞDk���ZO�\��~�<Zn|�d�����[�����s�����69�dBB(�ܯ�:}R�1��$g:�d���@�>Y`��	]��*]>���Ε>8�N�-�T�R��1
�@��9�CȄF�ح�)I��:%!z���ŪgW��r��*����4մ����!x�j�<�H(iX� PH����΄P;2-)����,FH\�I����J�uc@���Z�#�e��-^����e��x�[��$��ѩ��zn\�d��!�:�D�7s�85��dަ������ɡ'zTd��0�̨���1�S9��e�w81y����tF�x�W��tr�s%�3Ead��7�\J,j�s�����IŬ	 f(��z�i/6�Ä�,$S�bRFZ��w����� (����f^��>b���޵�x��z6#f�c^謄#�HR�z:�e��N�u<L��ݽ��y77A���O@SL����'��{��+?et�,�Vȧ�v�����ϲ:�e��p^�'hL�r�P��r._�m(����M�2L�T�)�d/��ۥ�j�а�	ra�z�"?��/|�o(����:�'c�$!�~��p�^D1���mKP]P�PM�_��ݣ�٘K?�.��,G�6�{%��m��^C�Ǭ��l�'%r� d�^%{���ş�g�<��i��̷97m��_�����Y^ܹ���`�W�bϝc��d���˕�������:�� �o���7�ig��=^��_0�E�����>r}����+�x�l��s�ڈ��_0��u�F�o#�_�޾��NX��k��u�k��ά�V�X��$W����w��W������MDL[���"�~�����q��6����sV������|�����#k���C�kU�Rl��o�8�z�9sL����3����?�棏�lE6,y�#d~�]~���!1e���q�����s��iN>�+���	HrY���gy�~����'>�������a�'��T�:���]�����w=�w>��d�l@��Sg�i�]��~���fTt]<ݺ��r��ݺ��͹[��[������a���cZS����e��MG�f�=�O�J�]Y����-�:ޑ�&�[w�̙x`Ig?E�IZ"���M�Q��u؎�'�zz��Q�dD��Zcb'+�Mk��Μ>Ju�t�R�X* �N^��7(i��.�i�٤���8�~c����+�X3��LS��" 
1(Ba�!�@�ò�Ae=�� �A
�!URqh�����q��=J���gq�⡃^�0tǸ��\�5WU�n����O'�E�)���&�����:�ۮ�@(��yU1�-ŹE����^�\���K����t�zK�}�O�Z˼�Ts�s"�Us��O�ч� !�.zY��1�c�)!i|�ib��6�@���<��qd�S���3���/7��.�(R��A$3��HB�a]�u���HBD�{z�(n����	ᇮ&���{R��	��)�M͍w^����q~�@�̮�plu3:�k?{�K�R������`t���);�7�8������E$f��Sh����+H�Bbc����Usƻ���'k#Z!qY2�d@֖����F(D���H��EF��\��i;��4f��ULQ2�<�^�K;�\3��Lg���ڥm&��fV�DÍ��m����OPd������].�kb�έi�Ⱥ�T�K��_˰՘���+T�H*	��a�h��K��+��uLV Q��eG�W�I��{���/�fC��u��V�쌾p��l���M�܏�/T�̈YW���r��y�����e�Onp����7_bw=�~d��s˵�y&/�ȫ��&��g����>���(r�hif3���r����z���K��y�8"�yD:���MIpMp�L3_�܏�`c������#�v\~�%~������s��èKWpo�X���Q0���6��f����<��O~�_ŷ*����������O?f4k)�����@��f�X�o%�����[3`��OH�!%��=:���"|��Qu���Hi���6���@$����`4(�
��AL����*)��l�� 	<���~�.Q���ʈ!$h2r`T����c��X�r2�ڰd<o�Ca2�\����jA�����U�ˠej�^:�ʀ �iŰ4h����[��,�i���k���<��+�����ԁ%����%J�����d�%��%P�dJvm�cq��D+����˒��?���dw�ڶ�m�S��2ս���C+�ںao�؆B(>e�RRf&�ಂ;U;6$��(E�d4���*yHx��IhGDK�)����Ԋ�M��b�>��e��m��a^Y\�]�P8@�eM=Ƹ��ٽ1�Sj��}6�#ګ�6�Ó0ƈ��~r2�ŝgϐi�t��Q
k'hq`e��_GJM�8&�y�Q&G=!:.�A��c"�,zdo]L?�$�{�M� �;��ةv��E��2��p��G��LI<9hC-NX�V`��3�z���ϙ�C_���!�|��
CSh�c��'<!�0�60�P�C�ȲO�"!N���i�(%�vBe[�h�.o�����7�D�}��Ɔ��*v���$�9�+.\�L�/�cu�Dz������\�)M�W._�k�9q���յ5��c��:F�w��Yb?GJ�����LYt�S�9�6��������;��e7��u$�!u�h�V%�LȰdTƓ�^�ՄJv�v�i�)�7�{(eI)5s;#���ѻ3LkX��qq���26}�݋��SZiY�ټ�ꕋdF�8O�#�\��C��^_�w����}��+�{�!i�A�l��+VVi���Vpe"!��g��^������ѻ�d4\%jh�}��|�p}�̶����2��ów3<u��G��ؖ�n���+T��(B�h���qF�7Y?q��cD3fP%�3��Wx�՟�����#�c�|�qVB�π믾΍�z�3E����D%X�/e!�2�b���ub1�n�~��Xw�lX։�S���\K�%��!S
y�չ6;,֜���S�X顳]��JEZ�;Y����n�vM���)�\~�.Ql�c�"]*�Lc��[��J.p1սC�(�R_�F��iei�B(�u-�ln��:�1�ߣ�N�"���\��]��&>H�cV[Z�L�>��ύ���uF�a6���I��c
@D�kHL�DBe�(��-�M"tenȌ�^H�eM��Z!i���1y�w�������k[��(���e�!���=�|9X�t��'X�"Y)z���tQ\ ���2�����r�_���E���p�к@�VL�5!�12F�L��J	�"��5����Ò� ����C/������*��:�E����'�jI~�J&����RE*���c�    IDAT,����c:ܪB(�q�\@���45W.]�؉#�׷�����;�d��Q2�I^(���~:�s�d6��k��.�}�����M~qj�n��O����/ ��z����dVb�ŋ���*r�������>+�����k�*����|NN�P��	-^�1f�C��$�y�� /���؆�(���fc�7�\�!/{77h;���l��1�2��PBSh�x<���8z�=���[[����J"}dE�\ٽ��k�<ʑ�5���a��Bpm�CJ�DЕM��R���x�X�#t4L}�ۗ.�/{�	2����SE���Ļ����(�ƵM�v��I*��P;�PM
�^NP��?a�ƌA�$
��#��aqVB�y��96�)<� ׷v��szs���*ާ�i$u[S��{�ʈ�ic�����OV�(!ٛi⊡�g�X}��<hW1ߟ�6��z?E��ub:�CoЧ_j)�H�x^1�fTr��h�O����o�3�����f��jw�/,ż6O���; ���7�~����'9�����hn\f�4�ķ�����U��[�s����J����M?'A���<JAQj�<C������z�bAN)�K�`�7'���s*��A�d��m7�䮦�;ݐ_�aP��tJh"��YYY������ ;@Ŀ��yVuZ��K�c��������Nk�Vxپ>���0�!1
�lBm[�(-@| A� ���:MѴ��%4um�ٞ �F�������.�A�L^%"�V�E{{�09v�B�[eK����
��>ny���nya��+Į%��`]dk7���f�hqC�,�Z)$�H�\�u����bR��ZO�>I��d�I��B`���������~QP�i!w�%��Fw�а��xZ�X�P����Gl� "h}����tׁ��B�:�1K�I�A�X�,Q.n��׷
�"�eU]su�*��68s���^M��	!T��ʼkj�T�ƋԶ�]׫�.�{Z%����m�J������q��v��ƀ��ck�F��6XʬA�{�5C�GT-���L�X��52W̚9�h�¡T���h�SJ�R��'��	�'%5���8�Bm�f���ƾ�ݵ�֨���2�j�49nޢ�3�3�� �g��D#���g4ȹt��<�SE�h�|�<�љa<�"�cU�r���Ԯ��Z���,g�;!�)�b�H�M ���Z�ld�]�d9�%}m�'�`Xп�$�����h��xoq�3S�����e>`�J���\"C��-�������qOTk�6����YIa��uK^#�)��1�W��;f�#��R�����6�GD��MCF�T���)�l5M��V�s������5efPmƶ#sI�b�4���MYE�N׾�92ϨD�Ui������P�T�R!�E�mXk%���_�3�r)]��!��IPl�
���.%�W��.cw����ȩ2�+������׿ʕ��G�~������Z"]̥ï��5������~q�	wA'��� L��D@���%�43R��=��I�],
��8��R���I
�Y(�N�_~�*�,m��B����T�Ъs�s�!	��EDܸ�ƩM����n�W��2�TW���y��a2E�_P�>%HB�˥�[�9y�յ�=g�*]�z��j������&n��%�2C(A%�ji�*q~���	���q�)�+��X0��(�t<.��S#��X绽%��y޿�9tQ�]t:$�io:|�տ�����Љ���h� Z�%B�L�D,�D'��\��Z<,���������r�Q�;^�I�BtJz-ѻ�V`�~�3�5�jK�2�bDň��j�B�+R�Ԫ �Q
�X�J�bLǏ��WLf�Yd������AEH>�%�"
�|M�D:	���"��G�$,E�*':rL\�X����!$H��yb�d�Ϩ��=Z�M}��.p�� �MH}��%�X"��XH슮�>�dj�[(�(����5��������N�BC�D�RۍP
�$^D�Y�Χ���}�c{V��Z�u���(�a�@J��t�fqu��c�B�A���R8|փ���J���jK�f���>����1�R�MulJ3�׬F�(i��5�h�U6uB�@h[���F��9��,mh�*b���2Tۢe�*G-�k�B�G�D��
��"�F��\�D/�tIQ�Fz��޳����FG���,�*궡���M0h��i�W���L�bh%�d����'�&[m)��m@*I���t��✦�`��y�
�B�	I�޵T�/s}g�>&��2���bҐ�M���&�Zh�������Ϻ��h�3lc�Qqm��<�8穛
;����� Uƞm���N�9�����.R�9u�`�}�B�o�U���	�)�6���A�!4�U�Ԉ��IAkF��eNi�~�y��B\^b��b������sf;c֥"�kB)���32%����E�ۑ)"J���HXh��vZ�j�2=�� e��;���<K>JF�K.$"ʔ��ź�=F�>�ʠQ���	ε��"��dC�F��]c�&*��s��i��RР�B�P]v���?)P2��h�6�$&Q�ӾשlidDZK�7F��<u�w�@Y	�fE�ґ�����QA��D������PW� ��)�>8�udQ�����v�3J D �&�u$)�|R���e���`m��"�o!�lۡ�
#X��@^�~���C��2 2�V��d2*��
A=����8�k����$Vʔ�/"(ՙ�I.�����"����ڼZlL7E� BGIu�[T����B%V&
$D�t>�j,6�4p�χ��
my���!HF	]�A*E�}ڬLN 	�4���.3���([�%�u�&��`�۵����0�X*�Ԟ����|>���&+p61cM�#8Ǽ���|�#���L��Ȉp��N�Ȍ�vDb	J!p������#t%�e��a�������Npe��<A��(M�Λ�]٢V��.:�N�"X�I���5D]���5�����JCM��C6@�-r�N���S�r���&C*�H�>�/�[�x�����9�O�u��dX������s�R $�h�#a00�L0J`�<�Y�P75���H��S����15�LFM��#>�r�>���*�	�y����ֻWY�(h����>�V����z�A�Vx|��C�m�޲Q(4�j2'/��k�K�sDY^� ��7h<jZ�a)�����!D�;���1�:F�G(�ّ!�xt��H���3��Xߠ|$J��\�!��Yݰ�w���8�v��"�&����"�@?�r�LڐH��9L/GZ���A����f�Rb�'$f&�e��;2�Z��Ċ@j�o��䤣`]llQVSG���]��kL�e�4�,K�8/Y`Z�љ"��$��du����6�E��X�^�߅���S*'bD�ĳ*L��"Į�� QJ��ă�mC��,Q3�L����-��K5�[N�Y�������;%r�B��u���!�U<r�4����[VQ��3�V*zBe׻N2�)�$�>ou[c���x�N�<2b0\aj���+V�=�X&ލ���^"�� A�.@��y��e�߹@�5�LQt-{ ;~�Z;c\ �,�T�k"D���x�=�p�ub�Y\�[����;`�K���P�a1�E=HH�\8����IJ���>�8��ۮ���-jInW`rE�i2m�R�Г��+@$�#!#Zfx�U5U풘��%'v�_zs�C�2��˖n���e��*2������Zl�׮��䙓佒�x�=�#��nҺWZ �"��8i��&y��4#�A�B�{)��G�����Z�r�����"BL�.2�edH��-~���p�{�E�QXPe��3�I���l2��}��D������dN�����\D�@�G�14���x��_�?DA����ơ����o���!��2�]�xh��!�u�P7T�VB%���mkb�􊌀$���O��&�����ݤmR��n�?��c����b$�5u=��잭s����VXy�&�!�oj&U�d2��WX��j�n�ĖC6}�쮻h���-���MÍk�_�N�M��m�{n��=�õ'��FH�a�ø*@h[�{�l�la}do2F�9��=���Xkѧ��ɍ�"*2a�Z"B$�K���;�����&� mK�#.�q��Y�h�g�4�l=�=Y��wʘ���1g�"j�)hG��w��cL����Ƴu�<�x�#E-}_tk�"��j�s7M��y��2�^��dW��o�0�]��T�X��ۨ��#u �A��B��F�@�Ԑ4-50�4M6�*�UY�;.̶z��{3�8Q���;b�o}�[H)q���E�W��m[�����$�m��ZZ�`R�XO��%�Ih�h��c�m+��_�~g?����փ�4��5K�0ą�T��^(+��ޓ��s@�ʛ���T�\�Q���#xEYL����n��o���=�}��<��T�����k-'ݽ���p���$��Lrs2���5�H���GDG��o[޾��&��7Lt�)O6��4(�*cryTʌ"�>�����i.y��ܳ��T�P� Sj�y�AJ��K�}az1��#��m�#����^o�l!��y#�j|<���]F��ֲ��M)E��'������	d�\����=Mg�����z�WDL!(��(E�伏��x&<��u���l;������S�I1�$� ��q<�,y�v��cp4��w�|�UbϞ������_/�X-������Y᭥>w���8AR`�Pz7̼nB��CJ)�"I�c$>�.�Mn5���>�v�"e&*J����3�A��R���eڬ8�jT�#�	�u�A���NPj�q�s{ͤ$(���f��x~LY���WC�;�AU*�n��%E��Lf���b���b �u�k~��G|����д-Zk��9릥��ԓ9��!�C�<R�v"x�`{R�T�@�4Qp�������O&7�R��"�=/~�|�7��y���i��B���b2E���|�E�\D �v����ڎ��5]r��E�U8�6�~v�>d��'��b+2�!c���������� BOFl����!dA2,Hʀ)��b0B�u=��-]��mÝ�O��D��%M�R�j��PMJ�ȃ����C���?��?rB�#�B�O%B+�o;ʲĔS�����3wa 3�NL*���؄���11�k���}���V��������-��Kd� ��*��~(W����p�(rm��Q�E]!e�B�m��+�������?�o���]�(�����S��ѵH!�E��bR�C�C�F/��v��m>�����c�we��=I䚹�b �%��D;�8�K��1⑨� �h:O�9��`?n&1��������;2�`�¨��?��K>џ2?=�9iY-W���:I:%��4����\���P���ͳ磜�m;��%��3Y�Z^��pŎ{�C��mr+�H�F E��	.��sL�"�="�qx��j�E���2  �~� r�T���`߂��>�n;����xcBD�k;\�<�F!�:p����R�z�C�6�t��F�� 2g��Y��T��,$z(�D>�i �L𝨀P�����FbR(=d��{�В�;�?��۴��4pv����~<����[.���1�"�㤞qyyM�zN8:c{u��=�1�<d5�p̑��de�Bb�'OD��(���R	n��ygwd��:��n8�[7��RRY
SD�x'�li�EIYh
��RVS���j�ѓ�����Ft�a�\�����_���Ĵ�QV��5��i�p�3S�R�VP4�gZ��F���"N��K��g���,f����<9%\����1.��p�� ����%�m!Y&e�ݻwY[A�N6>1��#s[j��D������@��3�{�u��!г2
&���Ͽ��?�{uɳ����'.�u�NG�,LI��\���� R"�]��IY���?���0/KB��ڨp��Q^dq��O���x��9�7��
1�9�&��0)&xj�H����5��xg��Q��0Qc3�W(�6�xK�+DY��=�h��z5Ԕ#� �y2ü�|�)(��!13YDj���U"T&��H]��%݋�2�>��9�� �2P��%	�ZI����6h���w��ʜo[j$�2���]ܣ�P�(�)"<�g3�l�5��.x��m,��v�L���޷�	�ƄU޴5�-g�K�.s9d�!#_g���B��]�i-ރR��"�v;�����~��#�:�<)%b�5�B� ����~�[��{�}|���\���!�EA�ە!|�=B䎯$`bJ�۞��������uw�ك�h/�i�)�����p�l�� �x+��2��u>b�E��Ȁ�d�Y����vZ
rB�1��$�uwn��������)=�`%�jo�'�8�� ���ɳ�3+O+�	��e�A�hč��!E��N����B�Ā�B
*-(�>z$���^L�2>%U�CR�@\Dk�˚���KƎA��x�9<�} ���m���፨	hVW[�O<y|����,���v-Z�,��k$EFIf���}
��-�A�i ø[������+h�����cWk��ei���LgS֭�b����5�TS66�d����_�7L��	�:���_?cu~�zy�.�a��L�)Gu�駟�v+Jey��_�=�w[D�smE,	A�Y��ň(Kdi(JI*�\y�����������Q�����o��}O��.I��lY^��}�$��-o_C�k��t��	�� �#f��$�c}@y�	��S)MkĪ"M�S}|�O?�g<��3��Z���Q�3)��5������ӿ���xd�Ւ����NtM����G�ٟdb��+C�umR�$Qi.�)���㏙����	�,(s���<Yoy��K~��_���?P$��2e���bJ��Bi4.9"�թ@�4�R�q:��F�ɂ.r��.�ޱ��
��+Tt�Q�����prv�R��mpݖ3aI����c�4�8�R&KpAG���DV9�]����=FNJ�P�͆�v��15�j6�L�5k�x�	�$q�qG+U��B��P`�g}~ΉOL��h.�;G�J��q!Qb?�:���^{)�s۔ܮy��s��0H~K0J����[�F�VL?N��VHD2�����N����Z�p47��a�wm��E�����O�ō��Ӳb�o9}δ,xp�/S����o-�V$��l�Ȅ�3�03f���Ds��m-W-��rt�1��+l�����c�-������!
�Ȋx"�k�I�hߝ|����:�$��
��'��$+���J�����B7�7!!�6�۵����o��n��[���>I��z��1�6�$G.�T%U��*��#:zW�7�<,'&1�':��N}TlK�A߶�QdC9Fڷ��ߌ����я����k�sR�R�5���+s͝�ǘzB<*��@ȁd�"_HZ)�bp�v$U���j�Ӹ�c�o,������.�"3��I�m�)!���$m��c:��-ت�u�S���3�{�I�1��L�������I����⚫�u]3��f�t~�aK�Ͼy����)�d-)ee+L	1K&{�5�	w?�������S�L`��.Y2d������k�WW�޼��Oؾ���Ւ���A���J�,�+�3��I	�������>�������/�e��uH��I�����~��3���gǄg�������?���9��|��7Do3���\V��($R�и$R��=�ɟ�����<�-d
�!"�a�:�r��9��S~����o�}�o~��/-���'������6����6��)B��;��C�\1���ÿ��������%��
I��\.W�It�Rj�q!����Wt��m��d�O����Q%i?齣�Q��#�����?��_S(��;.߼�ճ߲�8'�	�Ԋ�rE���u���#�	��o���?c}�5V�sn�i�    IDATW�V	�Ȭ�<�r��SSNj�'��������R�1�n;�� 5�I�6�+9�v)���6xj�	� �DJ�"�<u�z:�m2BN2 ��>�1�Cۖ������>��e���(��K�B��t�m^?{�}��-���i��<�mW�չ�9�:yN�<ǋ��t\-��Ri�m�W_����=�<:)��#EJۻ�Ih�(��|B.���zt΁=���ho��B�{��.�\~�9=�n:z1�^���r�F��=�2�#��o���z������|�R��h��D�!���1	���Rj&�:�JچJdd
y�"��R�C��@o.�!���!�i	3��Rb��E�f��ٓ>C����G=�o�>D�	GZk�͖B̧s�W+�n���c�N�h޾�5��<%$q�#	����4 >��!d�E&&���鮞����f�����1N9"@HI��������u���=�Ŕy/���7/^���[�<¥@�%���v"��#�$Y�V\l�1*���rr$���L�*&%���Y*��y
�"i*US��mHF�./�lVL���@���2yK����k�tm��j�b�o���n���s��-G�r,{j�&H�TEn+R�")E���;Rs�<���.)gdY��Z&�A��h;ʺ 	����b��)�T��d�gϸ{�1o����%U5��m.��GZ�����t8�.hI%��ǜ޹��߷�JR	.P(K��;��b��>�����cI�{��o�ί��!(�'��c����h-U�)鈺§����Ϲ��?&	��j�7��~sN�mI�񑋠5]ױ�n�wv�lZr}�����"7�ʣ#����Y
[:!&�(�}bnf袠I��������	��q��g|��n��Y-�}�,'��-�d���9�(U��� �9�߾"YC(��e�]?:����V4L'�-z2ɶj�x��e������v��v8h+���;(I
-�r�u�3'H�s��6_"뼇�h��0�n@<3�J�Q��:�=����}�u�m�~��~P���-ᜄHb����Q���g���=}�G���xC8?�NQ�]2�bD�0&ϊ���3�r�Ń�z�˷�|��J�WK�H�mo�2YL!��
�@���m�(�F℈0ia���AnB��!~�w���)4�t. �Άy ��b>z�ȣc��RB���r��#l�C�|�Yj՘<&�0$$�!j���Y�D*f��K?d��Y�HSȈ��g֨��\��R!�����i4���;�.������������
!ax�p����v����DDD�0<v�"d�Zr�u�u8I���Z���)�4�E]�j���C�W�P!�E���c{E$�<)��
U�lm�������͜��!���)��KA�����O�P�ѶR�� %)cO2��&&.�Yƣ#ZUp��.R�Zx~�w�=�p��w�J�Z�(U喲�����;��]�����|���W�sG/f���,i����
��h7���P'������-��0I�r�%3~��o��'� R`ZN�6�At�z:��;D�'G\�K�4�=:��
��*���҅?���"-�P���.��� ����0;�<Y���5ǖZ$*�UDJY"D�N%R��\���7oIuIk�*h;�QU�Bз=����(g�'IU����g��,^��;�=��]����h%1�����5�+̤�~�=���5���Har���d=��LkC�m�T)�-�y�W���r2�	�������<���Cd�X�[֛+�m��-u9g�z�3l\D��ݒ�C	M;�!����P8b�;Q�d�uH똜�����_����bc-������k��h�}��v\�~���۞��^��,sڵ�6P���+Y҆��<*�(�H�5�����(�cJ����M���B�Y3���P!�A9-���c��%R���{OiJ&Rh(fU�O� M��%:����`��@bk;BLHS��m����;� Hd&�Ò�� ���ۊî�[�1��r�H��b�<@�S#��)��� 	�BԱ���%6<��g	��c)j��h�d−ii�����{<��t���BOX}sͯב�O�����~�5εԅ��,E�5R�	���*bt�%r� ""��C�p��rI0�('�#���@�@�d�ܫ�[�{�u�D��,��	�D��{�(v'���� �����Å3��k�c�`�`�C�	-c��W����c���Ū(5f *�4(�%����c�J��c!mL��߹�>�Q�mH�3p�v�K;h~�s�C˯U�]	��S���ۿ�&ӌPθ_ZgM���k&A3���\_�[���MӰ��p|z��M�o�dh�LȘ1\���ǝ�ᚾ��{����ˢF)�����0�w�r^O 6;�Ч�����]�8{xð�jWw����F���)�������dB
۷���rw�*~���x��ZD��
�%E]�3
r[�6�4���c �<)���	��f1�q����.d����AcU�)ɟ�ٟ�(���9_��>��v㌳��>�a^�}Ӣ� �<cT����\��Z^t�3���`ѪF��)3�����XKY�D"j`��c$�h�uD�~?vy�Nc��!���("���g=t� %��/�~6���3�� ��	�d�l^��畆���㻎iY�6=W��SЛ���I*�:C�z�t�TQx��!�������rͯ��'���?�(
Br�!X��̄ �]*��+�?N�ZS*�����k�ٔm�!��c��Sp�8F�%FJ��Y��m�=\��{�Iɶ�6��B
��$��-ۻ�'rh�REFLb@h�TYs]*I5�P���M���a��.��C�(��w����0f��ux`�RN#7�����v;���%���!r͞�DD�">$6�o���'�������E�SA<Hh��"d�3��dTb�M���򊢔|��N�NY�}Eg{����p$���r�͵�;;:&Epӿ��R�A�蠇>�]�N�{6��>C��ln?v�����b��}� �����Ic1b�Ç�JٰB�ɇ<�@J&e�G؊uŰ?I
5��r�PX/i�〚xc�/����,��9�<q�9�P��Ϗ��}��p=�L��$��v�fuq�����	zRq�l1RO*|�fH��3tB�HYj#��zSZ�9���;�w���~�����V����ݽ�(��i�ێ�uĶ��^�˟�� �S� ��(�A堇�׬�T,3�u�&��w���R�Z����W�W��l�֚�O����Xm�\_]f�y���)D겢�sf=_�8;;&i��J�H�Ȋ"
��3��9hN8�}�s�-������(�����Wר���2�I8�p����G��⚖�i��C$�=��p����r�X99f:;E�	R(YF(rqq��_}��jw�B���m&�f��a��!+!�GL	;�s��Xkw�)e�l2�k[�..y��%Z*@дĈ6��(X�fܽs���ɰEQP�3�lʝO?��GO(�D5%ױ���kX]������.�$.߼�?�{��5��EQ�;Bh@�`z�����<�{�RI���~��fF���m	}���R(�s��͖�oRX��� ��9{t�{O!
MY�7�!�w�ڡ��wZ'R�)�싲.s@@n�;xS?��c�M�x���%��Vߴoc87�ﶝx�?��m}��9����#)���L)��f����._�eq���.��G��cIO`h?�߀R���Fbd@F������o�����:����c;��w�N��sr��U�����	��-�j��#�~Hp3�9�qg~�A��3�sVW�5�,�|��ټ�*׸� �(�Q3�M�� Dv�r62
)��7-�mO1|��>n��y���Lt13�%H%��[����=<?�[��=7.b!K������8����O鼧���S����(�k��ZG*(�@�1J��Z;G�k�L����~F��Q�z<���)Q*���ܪ�m�ۆ�.�\^�6�m*�>�EBi��F%��є���{���uȘXTN�����*0�c��`�-�8Y,8>>bq�������_ `82���$��8�|Vqz�����$�"��SL��sp�o����
)�ُ���ϙ���+��� 8�����"��S۶tmK��ҵ-��aF<�p+RQMg��"�2E�vKL��z���k���k�qͳ��RC�w����+���{ 	�$h=��3"�X��ƴ�-�e�ʟ��3TT�d�>���z��b�R���0����Gs�s6�����v���B���:E�m9)$G���0_Ly��	'�)��)�,J$2�C¹�S��u���5�v�!���|��WІ�oi6��͊�K����>�Z���-�6�"��:|Hh���O�>壏��R��R�RZ:\��#���?���x��Z0�M���8t$�DFBc@���D�,�((�
g�M���ɏ���(�ly�۶���;�W��c�I ���
z���` YJc�F%m�7��-�O�=z���}Z!�b�І�4��׹��t¨Di�("2yf�
��_���۷���=oD���������g���}(���}�q��E<��Cȡ�^AP w�����������v�u�:�R�$&�ط*�^�E'n���<�]fG���!
NBJ	$���s�}&�	%A���}�vJb��9e��C#}��t;H���m��>�^`p��}I1�nFk��4���/�`]�΃��bմ�� ���C�-���FE�Bb�0J%z�0Nq�.�Cp�Û~���2A"z�
BRO��E��n9�O3�9F�͚��,�m򻵑0@l�H�)'H�ض6�	�uD�2ۘ��tƴ��]����,�oQ�SO
�fó��z��C�v8�e��88w2O6L)���}��z�횮Yg(;�GJJ�	�.�VJ�v��j�������5�1\^^Y�'t�d����hZ�2���Np)OIL��K	)9Rr�ǔ��m�!K�]��cZOX^]Fgi�[���"��x�Ѭ7�	��#�1�R�i_�{5�3A�ZKi���jKsu�S�$E|��UI�ni7[�1���4R��9ǅB\���xM�a.I��N)95�ޒ����R+��6̎�|��G����������uv�)	�B猽w4M��޻���%�z�k;���eH y��;���z�p�� ʒb1er4G�{���=���@�˟��_��g�R3�j8�2�ޑ���f̳D�*e�KN���V���EJ�8�$H�ǯ�=]�H1��ލ�=�u~8X�]{v[|�]�������r��|�f�F���(��I�䫟��|���''\�����w})�@> Sv����'%r�5�Ɍ��s�m�S�o���)�'�{(�@s��o�>��p��08w�h��_i���w��bh��g��?�[N�m���ُ�ޜs�.��$���d&20�!��&�t#J!�0�G���{z�lDHM������È��!@>Y�'?�'�	���#���A{�a���;n��m���};�g(�`�S���uù<|x�ӳ���,�*]  c�R�]Ғ����z�bȣvo�/��:��fT���ٱg1��HC��)�B#b�Ԇ�ݢN�a8����RF	i/�f�
�u=�u��6Ȯ%G!:	RH4��zu�st|�Z����1���C�e��a�zK�;�l�tyr�NU��#�����"!$�ϝ�}ߣG�r�G�"&R���Qx
)�#c�.�fn�T���x�cV��$Z]������
�3�r�����$p�%Ȕ���%u�VtJ�vH���<�Q!�F�T�}��;��΅!,N�8��3	w�n-�Z!�P+RVg��c�f1����k>:;&�G���v�v�$�!$>�sYMi6+қs�;O��,j����_p��0�'\.��|Kg��ח�c}}��/_pr�>E5=hN� ��r�2xCr���5���m)w|&��.+��	��w�>�4��YD($
c�R�Nۡ���D�"�1R�-oe���-� zXʺ�,2�d�>￼�5"g]�к�����x�KB�]S�m�	�t���}���]�ۈْ�6�}��}�q�EH1LY=��?J)�fë/���b��!�h֯�0�rR��#�U�ȃv�Q�!�h$5�S|ʭ��CƄ@#�H���m$�}�)��Y梉�Ba�W��ރ�|���������j4.��pH����݄'���� ��l$ E�ഄX�(L��a4�z�m���d�� �3@�Ch飠�z�A�n�o�!�X��&�.�MG-���nrv�,�%�ݮ�v�����(j�q�og�q?�QJI�j�����7<|r���)W�m��3Lk�$�����4O�o	z)�d��C��|��}Mc������X�0�%��1RC�Uɫ՚��C|�Tu��(�R�g�H��O��έD�bq��蘵�XR��ozʔP�������7��:�M8ټ~�-�`��u
�53��ڎD���Kp�~pmC�Y��훖�uTJ�i�6%�,�����R ���k-�Z��hY�]o0m�qa�R�wB+
m�6����'�h]Ć�]P��ೞ�(#P6�ҡNC6�j ��h����-��cJcr��qXQq��R�D���[���Fda�}x">8���ux��*�i�{.�r����z=vr��A	޼}����(�"ؑ�Yo&e�f�aڵL$��������ÿ�P�
�}�wR� �������%b�i���Čݦ)�'��"�]�ؘ!R#�'j�p*C��PH	ۦ�K��q��ﱸ{ƫ翡�l��#�B�S@��Y�mD����x��F��,%Z*J���]�)L5���՘�t��|Ht���I(�t#b�^�{?�(9��(��>�
�w
�A҇l���!2��[���`@�w�����$o9==e�v���s>��NO�rѶX�bb��>)č3��ZKdXk�&�����k��f�י+!n��b��DN^��8���[���Iʛ������UɧC}�y\����܂Q���j*;�!��J_<�	;�=Ȯ-��2��ߵp�7~O���N�Ć��i炜�Q2R�����Ma�ß��;!ҍ�rB������y;|����]��̢ۤF���%���2j����Ͷ���,N��y�v�$���9XP�H��(%F�!ɜ���~��ǃ��qw���򽏂2&C\b��zuj!�h�t�ủl��O���]g�Vr��4�d7IPO�ܹ\�E״l6�x@-��hN�M� �!�	-IIl̰������ч<��(ݖh=M�ж-�v���[��)��~{N}E�=��%�u��!R@Ę���׳4����ftmK�u�bʝ;g��(�!�Y����E����v�D]TP��.d��ii�H��Cq*䠅�;Tz�ج�\_^q�{�)��8��5)�����n��(P��}�z�u���-%�l ḘT��BӇt�<2��ȃ�r��ry���c^>�����	�,��P̎�	�5��)�A���_=�ُ~N�$Rz>��ӂ���YR�
����L&8kѦ�����L|LtQ����c�D�%U��	M38�@�w�q����;�횯^���L�Ɛ���jP�|檤@+"Y�@Hq�Jc��H��dF�
�k��SփWJ��'C�R��тmے�Қ0�T�QN{g�>�����[�A`�H����~�v�I��{�{�������-����>���ݻ���|���hJ�Ӕ�K��h�����p����Y�>΁��e����}�o�2ȉV��Y�)"Y�̆t���W�A=mX2u��_��2�{.fr]�h���)	�'&�4Y�6Az���uL��f����l۞���"�J%x�}"&� R&�)��O���T�Q�Y�B�ʭ1>�u]�p�Ph�3���;��c�2F���/���o�[n;dT�"��$%	:k�'5��8|>N)�nz�+�����W�h��V|IV���$��L��b    IDATd�Թ��ؑy$*kR�Z�BH���Ie�b@�P��`S@�@�JKZ+�������۷T�N�@�X����놯���/������1���O>�;g,�|FstD��K��>���������S����5�m����+��t��\��K��j��	W>Ҭ�h�@���d�ݳ;|���|��g<z����Z��!�>&T6�5��mRe����&tE�.A:���v$�fbWy����mt��3LQ@'���m0fʀ(�f'�r��1jv����)�r=O��m�O�.Ydt-�È<+��=1X���Ϟ��^RΠm8�tĤp.z
��E������"
Xy�� qi�"���$")�r��z֛+"���r�+f��׫f>ϓ��۞�r�O~�3^�|MksO����(4!v�&R�D������"��2�v+b!H:"cC��.0iʝ�ߥ�
S������c�\.�h��T��Bj������$%22��Qx/�'���L���+��U�O��dZ����E�*80뭵�2��A���0*�%��p��!����aQ+�"Z-J@�&J�����@W5C�����́�I	3��;�02ە �L\�;�8���0s�#�)# ��C�����1d�	�y�1����@�m���LHR���"�����_�|uű��ꊠ%^F�� �\0�4�*5A�u ?@��ID\ $*E)�ޤ�L������G������8?�y�p
�|F�\��yA"�BN^����v I�ah[��[��ZLh�P�!�����y�XPv����f��sۡ���v�|�)�vБY���co;Xd�v�B&�;&�'���r-s_O�ؾFr�χY���o������o�7C�z�n�6��3?cv�p�4�~����svvF����-����2�)]�>O�����#����51L�I"S��H��� �A��λ�Ze6��[\ہI&�@�����)(�F ��K����jŋ/x�����jE�4���<��������/'S�Ն�:t�v�Rc���;.^�]�*']�J�����js�1��1�`(Y�1z��X�6l��T��9��?�C�N�s��_�r�K��9gc��ƛ�9����.�	�{�j]�|Oe� ��a�ZE�dRq||��-9��x{��K��Y�N�y1�l,��I	eJ֭E��==A�Vr�@�pY'��ϑc�a.uY��� �9�L��a�7xGg[B�TU�y���ꊙ8���w?壏���4?�я��|���Ȥ��ȨKӵY	OJ&��������1�������Z c�]OF�����c���k�$�)sBr\�=�_|A��;������;��]ǫ����g�MGH���"��(*�
��j�WW+�|������?��w��	�7k�ߒDĤ�kW�mƿC uVv��"�;Li�͐���>"�CYgxc����:1ח��g��-Ю����{M���{/|��8@�����6�}����BbL�$�s}yI�\3�̐^�w�v�u��:���Jc9f,�J!d\f�ܔ�AI�ᑥ��;�����xB��sT̏�\]]��@uim�?uxl�3��{|2WI���q�!E��v�=$|���bpD�P���+��H9
�ffo%�n���͟�IA��v�ޮ;�7�~����C��s���q���6���w*QJ�u��CEx��.���/i��P��r�H	)�!_6"	4Q�(��bh9i`�Ɣ���s�ܷ�ŘKB��Q>d�Zo���%G�W�<G߉L�36H���?h����d��	k-���3����w���~�O~�K�vÝɜ���ѭ�\O���Q�����b~J*g,��GǜM�D)��������eCIdzV�5���˫s���q��$-�Js��#�?z���=8���Gތ�q�rpҩ	!s�4U��j�,�9[�)�!�!ͤ����iX��xow(�f{��z��*��3_|��i$�n�d��]�%�����7�%����=�p�̼y�*VY�H��D�(���ڍF����@��0�����n�b��*S�HYŢ�Xwʛ�7�Þ�aGĉs�䭲�(d��8q"v�ر�w��.�lږm[���	Yn�l�l*�XhĚ���uӰ\.Y.��3����������M��>����K�7���"�-:�~�hf�)m4�M���|u�������y%�����яy��E�=����Y>!Ӛ�(���!��&F��seB�t�;���p>�r�Do^p����>C��l�8�l욯����4�%.颤n>��'|��߲���ưX���+?|ȣ'_AZ���?'f%�E���n[�4d�%�u��l�l+��?��ι9D�c��Q��������i3u�LD8��]h�i��6��%��r`�qt�9�p>��6�H�d�]�K�
�s6R[s�5xD"�ܛ��1#�pߡ�;��?�R�R"�!��M�02!���%��XF��{���U7��q�HD@ң=��][���5���Ĺ�Yua/�{���a(1��؏9��� n/�n`_Y���iP�����[�v��MR�w�1��:C��J�kv�xB�A#���u̲;����7��@�c�U]�tx�c�h��{uq�҂�LY��:�)+Z��t���QRPf��$ p"y�1*�JFH�:�G(d
�R�s)��=� S��Pp:�"�K�2�Ŷe�6��Qw��E�3�LY��ԛ-JJl�R������eL�k�^	2fbmj�iC�"�Yɬ��N朝ާ8�ǫf����C^��/�y�⤜�����8�q>rqu�v�AH�7dA��Y&~��R)�^'�օDIk�F�Ny�-�����d�)+븾x�˧����K���"��j�a�޲��4Mӭ˴~����i�O��ڣG�gPe��3lt�F�w�C)�?&fD]�(�Ѻ�|����_c�4/��H]5�#�n����YK���r�w��u��W5,�.AF���.���:�4�m[jo�F��O�~��|�BAuˏ�c>��246l�e��Po�e�1r2/89��MB�a���ж�f���$ţ�L�z���P��IA�|RT`~:#���7/>�?��G|�˿E���MU%���C�S̓I�÷�e��S��-1(���j*�&CǄl�|�Ͽ�/y���bM19�!��Y�O�O^��:i�#S�TtL�%�I����چ<��Y�P��xJ�;��%����L��(6���c%�����m_$��s��/:�s�������J�J�F�P,)��L�c�~8o��eg�����B@��ف[j�����4*Igv�K�����[|E"9��Q*�~� ��AG1��w�Tr�6V�T�b<NĀ�@�׻.�(j��~o �Y�PQ�qW*1�a�{�u�D�cA�`e&D�3�1���s�l�Z�Ǭ���~;�&��E��;|6:vl�Ǯ�ZJI�5�0�W�.i\Óws����k|S3��8R\W2H�J��B+S�#��0��4v�#�5F���̤�p�Sh�4dENP��#���M�rM;=Ad9���QUV�,�R�v�f��2�L �[Ke-�����s����F�5�����nȳD^p�Z�}��	O�ݰ��|�=|1��T,�	Z�F�#A���3���� �ٌ��׼ڪ�WU�pP/#J
\W����BL�p�łZ>C=z{�O�է|~u�G��v�_"��'T�G(Mk=U�e�F:�α�EvkAt�ф���l�H2�j�j�B�	�(E��6)g�:|�ȏ����e��X�ߠmCX����iۚ�l�2k�@�-ѧ���fC4LJ|S���?��1�����>��r:ek#H�rP�Mے�"q��T�S����OɊ���l�'3
#^��ɦ%�ed�)�r����O�����5�bC���:�/j���L5M��5�f������cb�T�E)E�e0��4���3>��c�k�;��NOR�h�Q1�[O�%C(ʣސ���(
�ɼ$S��i	�v���`�%�{�S������ܫK8N�(�Z쮻�Ab�ý�ۏ�.��'�������
��{J>&�C�>�;���{�kғ��0�w�c8�o���	1t�=*�}:=��%Do����>�O��{H�	�H��v9�!бi)��cu�BO��{����F��$����n� {Xe���ev�L���ޫ"q��7��g�o��Z�����[�����`J��l�c�x<'�^�]�cǏ��.xjoW���{C����C�^@�39�+�
��b�Қ��~Ľ�OX�\��n0"�|
)�rW%��|�:�%1&�8�y���yچ�����=�s)�Nk��("�k��-��Z��5��9.WXkɵ�78�w��r�����)%��H��Y�-����v�^5LN��Īa4��)�G|/onX7-�����@�x���wp��U�^��U3��&�3�優C���	Ֆ�nh*��`\D6n�b(Bg$��h���!7�����i����Yf���Ƿ^.��x#�(��N��t�]pm�5h=Å�ń�|`�15ֈ�$izrB~rB�ג��z�6-�zդ7O�4��s�;'{���ϯ�.`72�1>����R*�&t�LD&ڠ���%5�I���5W}���klUS�L�����r���L���M��(6J�ԕdBP���f�馢i,S�y��]%�2)���4��������g/Y_���j�ܔ�(�23��Mǅ !��A)���9EYRw�􄴾��lZR�KL�@F\���L�6V�G�����&�u�n�d��ͤ�ZG�KN�r#��ں!Ӻ[rp�B";��m]R�A!7I��{��NEBVw�hO��!�Zq�����y� ���\���vw �	%��U`o���C^��i�wv��B�;�(�HY�C�C��QY�L%�Cǿ�P�����������<��,��a�+�8�קb���Gb9��.��{�R)5B���/&Cv$."y)c�A��튘2���O(�:��W^��F5�����w􊵟�c����w-����F�x~w�V�q���\;O~<����y����� y�+�(�g�l�9zf]-��.�A.}�i��tp]jH�A���|�"%���Q��G8𭥩S��sZ��'%���o�Je�zq�</��Yܿ��<m�%��4���������k��Эg&����]y��g�^���ez�Zb�'7=U�ٜ�,ȍF+sBY�I��<`:����l6�t~�f񚥵�\]�o��*5�S@�@�)J�#6W��U���=�����*Qk�˖i9#@ph��g�</��Ȳ��҉E)�m����U�g"d�1x��H�	����1���? /Jd���:	
��&4�x���կǉ*~I}�%�5��SNfsژ*1�Q��mKS���FI��z�u`]"�i[V��o��缼��ZI�sN�N���m�P�53����Ֆ��k^^\�`������(���U��WW4�W���ۆ�e�|�=���X�%mk��kT��1�%�����	m
�����Tb�J�CCnJd&���FK�f�rI+*L(Uö^`Q�T��8v��2�;2)rC���m�mcǵ�1�I�<�æ�<~���ߞ�vLN��*���|;��}�����><(��w��kd8t(�(y\tl|J��١�1�xS�Y�1&߳�a����p��N/���	��.DJpD�K�;fpDF��봚�3��fE6)�*����\�܆���C�N���R����z�cKR��ir�	��!����q�xb��?�h�FHM���>��{����1����˫�� i�АhI��s(�1i����������[�<��[oᯮ:�� 1t/�B��@H��V#Rݽ�R�ҋ!|����E� $:&>o�RM�V�LiTH�MUD��������l��ų?��-QFj`�^#�����E1�L��r��}�1�j�Dg7�T����Bi]�g��B�.
|k�e�TGTtDA0�
L�Y�T;�X�m=�>�y�ki���4e�%��ۊ�jö��&%a��9G�G�.I�dYk�ֱ٬�������|�O�~Φ��'o!LN���1���sTR UA����(d`�Z�Y��G�9Zv`�lB��w�E�.QgB��M����V]�d�(-�:�s)iS%H]60�	����VK��Q)�tFM��m�i��Ȕ��-�՚ɓGܸ��d���qZk�<y���^E��ε�7�_/��H]�x���1&!�1�M���򊋋�"*I����Q��>2�L��-2j�������\G�ct�1������S
�:�a�֊,��%_f���*�<��X	N<*7�m��dG��ؿC�ՔeA�i\��چ<�PBSW�F���+���^>4MK��JZ��ܧ���Bo�����>�ǹR���ɺ#���q۸9�}J:la��1�z���S���I��� ,�D����=������Q��z��x��ј��m1 �R�􌀾L1�H�a��&v�9��ίk�2�9mW�!y�=�o�!��M�[���<8ߒE*Q���I�D�ZQQ%O=8�R(����J�@"���Q��%iZG�$6ơ�R��!;�g����F��H��O;F��=L�~�S��cJ��&����LG�c�t��6�4~0Z�@;�;�]1��8��x�&Ϻ֍m�6)�\-y^{�߿��M�.W�()�I�Tf�K�LsJE��
Ik1�7M�]��)F "P��9����|����:���'|�'BY��cW�T���%��Ͳ8�,7X���lZ�y��(Dǉ0�8  ՜"Zdgӌ��E���Xoh�S�ʱ!��^N�ْjY#���P8�Pq���-�O�4V�8IU׈��qR*�c$TJ�+M6��P��'�-m�����p��cB�i�B���ׯp�3�́U�Ӓ���;���w�Fݬ�<�`�$QE�:y�!zZ���DC���"'/��9r�b�n&�f���	���ٮ���2��l,˟o5���
VFb��8%�G�;C�%)�kJ��Nz�R�-Mf�Q���ak�2�Ef"k�F�H^��l�(�tL�@�$O���lj�?9��3�UŢ]Rdڶe��R�5ֶ�M�vQq-+��kB�D�|RrY5�	:x����S)9���e� ��8�b��G�N����tJ�gSW�uŢu(-�����m����u[D�`"TkNf3|nX�����4d�!�9	ѬYǈbFnQ'�,ˈ1�Chߵ��T��'���t�o#.ڄ��5�
�B(�����
�"�D��V�J�H��X^2�)(y@{UvIbc�­�d`/�����ϳ��O�}�<��$"xB�!-$GE��,�Z��mED��M��#�j��z�h)"���"�Ó(	
�� �2�:J$���ɘh�{#�CJeb��c����Sސ�g4ZQ�����M�-��{��&'����}�����҅�m�?���[������{�`�C�c+�.x�������	���K�Lc���q|_��m;<���4���<x뜓��^�����
���u��N��+ A�h��2�&v���5��DE�]����_��3��_��=>��������7-�"��Oy��!�W�M���R×���DB"�>ŝ��N}�Uj43՚�sl?�����=�����O���{��l=�?�3��W<��ԫ%:7��z˛�HBa��R�̠����3Ĺ�A(���i1��dN���g|�o��-"��ϯy��{\-.�ş�9~��D�hچ�R����ſe�z�,+P&�:v(W��UGb��'E�
-�Θ���g|����=��q��	r[���3�j�p�ZO�����2	Ā&t9.N�"u�Ӑ��|�Z����B���Z�<��b:czZ"g%Z*~��&f��wߢ~����0:ps}��������
�'���D(SUuSB�(M�Fih�4y"7��d��'<</yx��i0��������Z��I�T���
U�M�:Z��Bmq�u��>e�^�� ��    IDATDT�,�k�2gu�����������/��k�T(bg$��c�*�R�,7Hqm���I�Sd�#p�v�3}��(bbI<!!�d��ZfO���{�ۗ�Qǎ�q��0�a�)�����9�������[���/��@*M�������R�H���^�������D�c��c�~��=s!����]춢�K��'n�7��F���bA�R00���sS����;hl<���z�:X7"Iq��E��z�֏�и8���ݺ�����H��S�{�J����)�`�ZB���a�p�ի��ӕ,jV��A�d@w%�.@����.vI!RDN����������Gq�ל�����e
2�������%���9W�6qo���<DW���Os��h	y�'p��r�ӟ�/�'���xu}���}N�S^=��|��O�"c��heM�h�0�(0Ju4�b(���χ0F`ʌ̗�k��-&������o��!���/��}�f}Ë�~�Z�FwIQy��u�O������ɻ_�[����EA���.�Z��us!��,EG�.QLu�������ɇ�P].y��-|ky���kf�$�Q{ANK��&;@�=ƀ$
BD_]�t(�J��8��i#�����'����?'�{��Bj�^]�\/U��rA��Y/	ŌLJ�I��V\��`[D�>Z�����9T���&È�}����	�~���92;��-��
�|�q��H}�Cŀ��"��RۆƷ� 9�\jT��C��90��,JJXHI&=/>���O�����FI>��_��?�K��F>4�RDRV����'�&*A���hA^�`���}흢�}rL�"���B���(�S�����;�&����"�
�샇}��v\��w�y��;��2�M�u��T�����Xq�QỶ\��>v1IY�����v�(JЕ,���T����ޅ�8C<�u⸖�e����m���]��a_���}l�!.�Q(��N�1��.��y�d�.�c����_����:'��|�6���x-!8�b�l���y��U�ｧ^�\\\3?���'�;�-�K���]�A��-�4�؂�b"FY� �킓�s�vI�Zs�2#�G�M��kɐ�ơCoz�b��f��[�J+E���-궩��V��B3/&�H�����͊)
�]��jCY�<*�Ę�@8Op�=�K4k�L�:~���nw�gd�Y�.3�JU��9�����������zAn�Kd�&S�*�*gY�=�uLL�,2P�YJ�� �LLto��Вe�#*�t:e"����◄mâ�Q�5�U<:�a�b�mqD�X,���Ti�ϭIJp�F=1&/�8R���B1��抧?�2D�I�N$_��o��xu�@�����,n��>)ܼ�1�h-�uC%*tH����G�1$jT)&sb`X��ŏ?��O�!3��3��nyCV��jE"��#0R��NpkL9VJ�(����	��OJ�Q��&55ɔ$����?Z<�g%���`a����Pyt�6�x�֑i�tR��@��#����
%p�ln�DŶq4�A�&(��(S�����j����׍'v���8 vyE�Cv�"����ߴ,�o�
B܃�s�?T�DG,���;����5���u���5��>R���^�*���!g�0H���s�zJ�~��6��؃��з��8$��C��������1��K�8������A0�Q��$��`��������5�nV��.���>���?��/��!1q��=8ϗ�<�4�/
-�����u��R�����%۪��WQ�9��X�(���#=G�e�֗ 
I���� x:�� $��加5�yI�u]�Ʒ�Z����9�2h���Zk�XL�S���]����a�Kr����d�:l��eDx�4�6LT�6��R2)��&yJB��3�y+�����������ʇ�9ND�"7��iIlk�匛����"�WWiz��l��S��V)l)�'ejHԽ���wDJ,�]s"RK������m��e�tY����[��1Y�r5��H��yB��"�sR0ƈ4��REDh����im�(x�4Lb�m�4�M���2���@w<ݵk�N@��,A������JƦ ����`c@��4���lj�ߢ��][r�RQ�(�;D�萤�Z*�L�7�4�c�ޑpU�q��n�%�lB���P�z�j�����sN�f�=�[+
	]3E����~e�d��L�#d2,;�)�cF�7#"5^r�<�F�]?yѵ������[rr�C����)��N����;�.�����і�c=��]��y�n=*O��������>�.�g9t;�b����}�0�c{�a����3&z�Ůڭ�njw�nV�T���G�758�PP ��uTw?�<�;���|��������qb�Vt4�2e�
��R�� ��ԝ���u���/�I�=Xo��Kw����>c3�⾵�������>�n�Yj���X!GQ8�X\/89�`�)�S|�����=*��Gr) �K/CD�c"Px�⤱+��.���"'&5Ԑѧ��R&ӂf��[{Z�ߛw$B���Dl4�ac@�"���Ȑ(����?D��c��v�����:5[���y�1�Zk�N�7����d$j��
雔!m�B�H�۪E	IUUH-Si��̦
���A�Ԓ��ydc�[�����ij���5X_SxK���� �L�c�jjB$�!ĈRI�)���d)�q�y��#��r�JcLa8�	�T��-�@��6�ˌ�/�B����\^�����\�T��ݟ�mAz�����F��O�^��8�P���y0(�w!k9�
d����Y�PGA��N�#���n���8�y6��ic�%�m<�j�L"��LsEK�]/Qn�=3�Y/�R:V_�k�r�|2%�"��������"�����_/MF��ԍ#�� �9b�8�&�9,�}rL.�)�o�ɏ�+�H%����~'٥��_E���A��돢��������y�S֏rt��{��њ�!�#����#����M �����(pJiD��.RJ�L�!�[��.��>��b�c���$����1{7"Q�+���,���<\��!=�n�{f��|�#F���/=N2^D�����uxܱ�1��У������5ֻ��eb���Q�;�1JѶ���KB<����I���LI�PB�@LW�S�9-Ơ4>?AvlyR!���+T�1F�4��\e����	��;��&��c����P�*	!��A!�EI�1�V�1d°�cr���%�v�Z��B�h��1�p�"�[����R�ZKvR&�}��s��l�׌wh!>:΀���d
a��5���iBde�}����zb)A�^lȤ��4��8��C���y��BK����V�J�V�u?��1��LkX�{���"E���=6's�%�����r6a�=��ݯ�������Tֳ�Td��	"�PY�}���+	S"��y*�:��9�4x'R#U -�O�*�QX�֨��4%�!>FHbDEʦ�J��Bh!НG�t��تAKM0>5=:+q�!m�a��b��	�2#����m�����ݻ:~������ZX��5��z;�j,;���v����ݱg +c�;h|��1ǹ��<�=G+��B<r�� 9v��(�NǇ[̥�y�b�Ӈ��Ů������L?v��k�Dj2�T�'b =�6�?�	y�|Kq�Ѥ����{�J;�7�Ĩ�aS�z��8;6 ��=E�{##����{�ͭ�s�~�c{hl��I9_��-���ޤ˿�Acb��'������7TUŴ�Q�)������9����c*�]xG���C��I��}�OL�T�I�l2O�W���٤d��DK
/e���jj|�)�!�@�c��tvs��оAi�$�X1!` ����2x�wg)sM^NX�6�̌`��q�4���1`�D@��H�1�=h���f�S�u�TL��LHp�IVR�nyB3�Ld�=���"������M��t!6Ij��T$ ��HyD�V�<BPSOsE@ɈV:�w��BI\��@�ƃ�2x�GF9$q�%~=���$���!b$�K��z�V�QeLb��)|b��^��+N�)�vd�lP��{P%^$tE�r':�R���#�@Y�iв@��!��"C�i�}E��9��\��PM�H�f��:�#Z�{�����׵��D���l�y��L��H$A�!:;���.%
���ӓ	1:���d��]����	�B`��RB�P':D�A����ҏ�ʨ�X��eS_��[<x�c��:��+�-+��|;���s9������Ȏ�-��~�{�J��8ܿs����1!����>�oD��zSj�"��*�$4�Ӈ�i=�I�*���w�i��PbG~3xx��(DJ���u� �d!E��|4�F��.PB�D���.��H4Z�ă:�A)3��إ@h��>�ej4	�uaR� 	�%��v�K�Cҝt�[~�p�1!A�,V+�P��Tr��� 0�.��p���{�iğ�%��Jއ�?rZ(I�wٺ]�|.'�<�\��,/��&r~~o=f���y
!���z:IM9����TĔi<��4>�x�2���lM]�0��vI���)|��+�lNn2��%��e[�n�A��.��?O��QG���f��^�����2z�*�1�6��ȶ�"2��5�e�L*�T:�2A"2��I�QvU]$D*'N%���H���<��L�M��y�^T�L5H�-���x6I���.9}����҈D�����(�ᢃ̠�[! �ilˤ�t�Ll��[b�h�m@��Vj�Q�˹�-y���W�%JC��X�z�TIF�Jn�g�)l[V7�xv��M� "k���� =eVR����/VL��v5�Ո�)y�DO�6�6�6��8Kf&@@��Z��&��!"|Hmg��SE���������O"S��CNr6���|�j<4.VĶA�	����k�&���w8!P��V��$�f3\m�L5NoQ����׋�m����7�bRҶ-�PXg)�%FT����iȤA뮕n "Bk�h�#*�V��F����]�M�|&*A�p��p�h\]6>;��vhꡂ~�HN[�9���H�aܡ
K���n�L��١���$���v���D��H;F�����D�ߡFr6t5�R*Z_���xD�h��z&�A
1��O���B9��� O��Tw)9)q��h�gB��`�۴��F�4	]"%&�ΰ2H��>�>w�D�1��ᡱo�ܵ ޴�ù#�,�@�2��踳Pb�����[>=
Ez�����-Ҋ�Ф=�B�p�������oh6q$���?�'}x���6x�_pLo��c��on8�͙��Q]��m���p������SDߋ@KEa��*��EE5�ȓ{�D�T�,BV���ٔ�������
��u�Wk���K�V�q��J"uɫ��DךVA�D�+��HM1�qM*y;�ϰۚ�h��\y�[ǩ�h#,������0'֦�����5�1�-����$\���Bf�Ep^��)�T��<+p�Ѵ�G�Q��b�$�-�k_g�6��LJE������f����u�@h9ӆ��m�Tf#&D�!���\E���2�������g֒�&�M�4
+,>��9��.Rd9��K�a�E�o�Qi#�mɄ&��&��D@ʖB(��)����.�dŔ��i�&q�M]o��Ln�FI�6������'�
E�����	�����B#
dVb��Tf
������F���|��-���q�M�p2+(���xV�b~:EIC��2U�:khs�|2Aw� *z�&��,���h�y�>�	��hˈ�I�)�Zムi,��%�¾=�y��ʠZG�6�⨛��p�l;4
��:���G����E���|������4��F٘��wc���#�>���Sw�C�?�]�+!}��!Rpk��Hzp0��@7�(S�T�	v��C����H�� uq[����I1(e{���E�{½U6<�>i�﹜�	�ւƋ�]��xBc�,ܚ���{��_��,��p�n���ۡ��w�g�Ѐ94T`Gpa�e�Z���޽S�	\_�d�l�j�4]ן��� S�q�=�7����÷��?D��X^\��O�����@��N5[�6�O�����V5:���(%�ۦi�1R5ujz�-���r��b �)��8y����D��a�4�OY}�&mLge)f3N��BrysC;�3=?���dʼ F���Uk��u�C5*֗��5�jhaXf9"��Ea&��Q�9�fCռ�8<s9�r]1y�-����kϺ���9h��g��ڵ�X�S�)�����5eY�I�k+�6A�.׬E��Z"��]�7�|���eK��ט��/�K�B�"%;�!b�*%oFOӤ2.D@��
�)"jj�d��͒lr�kk2��(��-�	|�Fi�uͣ�@���F�Uæ�	Z�],������%u�R��dдL�r�I�#V�l�g�6
�da%�s����D���q��Y�&U#�j���i�V+�\�L�H�����}��fL����z*0u`�x&�����cJ���V�%��e�!���)�Gt]�b�C�9��*f��4�������3�A���~�{�g��<�/��u��c���Կ��IQ����_Ӷ���$]ö�<�bJ��a�����F���0�w�X����w����x��񶗝1(�;�6	]�h��0�&1߉a��1$ �I	/����:�(��D�ؕ~����*�o�ЍW�M^С�vh�zӇ��g�hٷ^��w6Gr��s�uoo����B<�V�s�h^��狋������9y���������儺�'H��		Fu�]N������|�����X9~�k~���(�1�Q[������۬_/?�a2���o���Ǐ999I�V�\^^��石Z����z����)Mki�%�w��η��ߥ9?#WW���a���o�5W�����,6��	*�R�����o�=�҈n9�*�Gm���P�������ǟ�]Z^˗��	[+��������\����(g�ُ������(�[��t������]����?�����o_�b���Pf9�z�bq�B�ԉ�TY��s �M��놪����ۼ��;��̦%�5���'\��'��|dmk������x�ۿ�����WV�5RG��x��?��M���?�O�7[...p�b�5~Y�-��P��p�_��w�����w�����X�|���g��%gyN�&P��#��m�&#��Y���`=����dT)�p��d�,K��j�JcC�v0��Wy��� mT��UR�����f��T+ں!�(�Ӵ��lm�mS��J+�u�UZDB�b����z��%��(����op������5:[Q(��Z�m�Le�SY*!u]�\ph�C��K=DWR"8�v-��H�`�]˛����,�������x�9Ys�ܓ�cy�w�az��1;����܍Hz���c]A�Jy�Z=S �����;��?:.��]���_c�%2vN�و�[mkǛ&� �v�ߥhn)�/�S�	s�Q����@�S�ARL���S�Oߔv앻#�(wy��;���)ރ�{⇞����=����.�����y�I�Q}2	;�l���Ѐ�As��٤�o�ǽ������l떲���8D$��#�wz��[Oń��[2y|��x6�"�e9��f����,�!...��S��5�����<����<e��iZ�uJ�")&�t����w�ż�U9*�d��n8}�.��%/?���>|�j[S��K�bUb{S>Bp�(�F��v�by�����Ʉ:��֣�	g�3=?g��|��������V���M@���b�U��Wה��Q*>}uɳ�BV$�������������"��i�%3AH��5m���'��٧O�^�U��7~�o��wx��D=�G�%�i��d�է?�����Y�4�    IDATa�Z��//�˂�����S��mXm7�Ր$۴-mS�X,�뚸j8�j&�	n~�[��]~���/(�<"�ȃ��_٬X�|�G��?��?����!3�gO�nZZ��������9���d��L�:��)4�m�����n�x6�5�z���Lq턳��M��O�������J���?��+^��!lM��b�%��V[����{�ɍ!��S0��pu}�r�d�ڰ^V�@��8eP�$��P|�]�����_��f�l��g\�xJvr½bJt-�h똙$up�h���н�]�Q�ZOӴ8Q"��G�`��s����|e#�pE�+�	���Wcgo������}����٩�7��!4ٍg��%��#��Õ��1R�q����c��T�ػ���vc�{T�q������}�[���t�Cƺ[DW��I�#�[!e�S�	vJNqU��مR�����p�.�@�4"e֧r��a���^��xW���+�/�����T��`W/?��oǷ��G�`���!�E�]�#t�ָ+aO�k�aK^��9�͊G��9;{@usM�<�[G=�A��������dK��~ǅKW���w,�3$G�j�AX�����A�A  PZp��pgvܵ�\����É��̮���+3��	���5�P#4�i��YF�h	MG���d]`����)�5e��YJ�e���u��g�^l��u���^4��0������r����Z	�M >@����%e�\C1�p�;�e|r���hf1i4OH'#�R��w�����$I�(EY��8;g�Zl�(-(��:<e6UHb�L��+/eK[YZ/Hs���������S��1�bf���9/~��s��J�Sܻ���v��t8��֭H�ί��ox���\�W� �}��F��	~v�҆�y�|���mR)�:��.&4�������G��S�����9�?z�x4���W��k��IS�cH��Y
8�}�,U��C����8~�y�1�ME6;������/Y��OI�5��RA�#T�Z���eSsU��ʐ���h�m]dl۸�jI�j�r�Ã{d��YF�x89&}��d%0:�Ν��.�9���p�Yf�|�U5e]!t�����l�x\pxrLZ�X\]r(b�rkS�P��-)Fb4�,͸g|�?��?�s�����6�O������ڎ��A�Q*�	��QUkTV���P���RH�	R��������k��9���rh#/zE�-��>l{��/{_H�&��F�aoΛ���~i�x�[���P�0����-�0�m�z��j[A��U^�@������A��4�� ��Q?z���!l6��#�<�����^��W\�}�{��c������Qb���vH��.����!C��k��ii�qm�lǧ�!���o���x�>��kq�|�[�nw����>!D�t$zC�����m�L� ��㾽��5dENhVWKFiƭ�GH�8?{�T���-e���ÂJ�.kή.9�JR)I�&��ѤM�u��Q���ڎy[S������2ҖJ)cC��:��]/��B*Mb2FI��3�YJ"B�o;d�wH�C'9�ܑIM�^Dh4��P�UE<y�aLB&
�"vv�IJ��K��Q��hDs��M���dF���mC
>�L����}���G����5��iR���_�րV,ʊ�����~�ܺu��ш��8{��7o�x����^�ؖ�t��񌃣)�:
��Ф�@�X�T�?�%<��Z��L��8�]��1�crz������"1RUל�������!M@�͚�)����@`F#�ֳ�+�R�5T���Z�4���oKݵ�و�xJ��/����$]Ӣt �&�	E>F�1�\#}���;�	�j���/������	���������� щ�b����<�c#1y�j�B*��l�B#�atPp��!_��w\VK>98���:O(����%y����	�?R�~A�ZECz�E'�o�� ��*m�h��Xd�ї
Y�(���v�7����6aƷ�w�}2sB��Wq���)�ߠ֡ϼa��~P��З��0��'�o��8�������ݞ'Љ:�ygP;��ߧ��m�Om{��� Jw�;bC�҉��B��D��`6ǒ%b3�ᛘ�qC6�������s��o�����og�o�+�.\�?�����C_7�=���p���^�Pi{���s�Fp��Sd#rU���k<��{�)gWx�!|ߩv,�i>��Y�<uW���#�G*��y�L�f�!6?qm��ͪ���e��)%�)Y����5��#&�)��\��%�k���&! �e}y���L2"%L'�ɔ�9�k�u�1����΃{���D$�.+��c>�sqq���3���n��%�Ҥ��5-��U{t�!���jR'2��jn�f�b�S�bĪmhҜV�b�����y�x�s8+P:�Z,Y^�!(��-RNoݡ(2�h�LQhO��,�IBP��Y��qBSu`@u�ų�>�0Is�\'��/~���|�h��u��h���yQP��m�k*��iaP�<��*$'�d���	b���*�����9��f!HlC2��Bu���ylg��{�6)E�Q㴠[k|p���hڦ�0)Zڦ$ӊ�$46�ڀ!ZgcY���b�x\@pX���#F��6@��W�������锬��N&5��.GS���y>��c����ObK�����<��8k�{�Auy{R4��Z|0*A�H�-|���Ç�����c�Cv�������Ok�/�������ٸ���*�~���ΐ�������o%oǏb�rn���rl#$��.��y)v���=�Jz�̳�-nLr�:��G�Ҙ�"��]��(���|���oKI�D�����^��R���V	� 	�F�h�L�x+,���[]JA豪���_8�q��%"�ޭ�߆��D��>�Ș�t5Y�㻈>X� 5�� o���뙭i�|����M~��m%��o�M1y��bc��\k"&�X��'����H��o�����֬.K�m>bI��	VAJ2!ojU3���
C�2�ЬL�r}�hv����͋�����7tA`����bw��hL����5�d�����"�7ۢ�SV��h��C�F��[W,� �3��+N�{(���(�m+xr�>����3BZEW՘4ź�y�%#���=~�Yy��Pԋ�?<�+y�7���\�����5Nu(/IӜ�㔑��Oy�3�M��і%�:T��F#`u���.�Ԋ 
Lb��Ç
I�o2KItF�YT6�3
�3��h���N����j́�!���rx|��*8��C�����y�O�������1�<g~��mU���TU�l6���;�O�����������SJ�f�&:���0*ܕ2��$��!+��st�RjM���;JC�rQ�$
R�P��.X�"��).��\Rsb;f��J��a�'� �')F��c���ǡo�5���\E{uF��q�Ř�4�8�2�Z^�]5�u4]�A2fRL�J�`r���
�ɕ#�L�1��/y��S�b�o.�drFz�!˯^2j*��ۡM�s�G(�2)���e	.V�(yB����S����2h�(7u��*�k�p(��md�>�h_��Ͻ=�e(+�=+�s�-ټ�����^_��5IP��m� �Ï�S�?�;��y���M����Gqe ظ�$UX�#k��M�cC��t`@�=�=� b�,����y���:h�A����@����,��b3�>?#8�1<���,��
��랰����n���u����f]3~�X��O����F4�_\w��Y�pa.^1x��!a��|;u�!!�zOՔ$EF�Z
��u����*�u�)�P<�}V�M/۷���{����y����F'
ږ�,y��9��Md"s�"�霣i[�ԤE�h2"h�zU�'ׇTd�q�q�.�xl�Q�������ׯ.�<yQ0�2�Ƹ�dr�t2�0�q�,y&`�'�&��)I�T
�F:�4=��$�w3yJjr����� Z�Mg[%�lK$W/^�������)9���YZ�:OPn�A�4�'�%��@h�IA�',E �H~"�&�X�2�0&��ey�=2�G3��1F�,e]�i�-#��1�.Ԭז�jI�6h�zG�.!��ږ��Y�n�͘NOx��!���=W�ͻ��!&�	'Ǉq8=!i�\�ר�ùH*�Cbi���b��a\�p>�Js��A��i�g�}F�T\�y��՜�tF�����FcD�����fS��Q6bR�LJ��zB�:�L�B�Q/����46�qr�6i���!�^-,���r��C:'��zSJi�!���׶mo�JF��*>�e]�;A����W_���o��;yx�c�r����jF��s��B����H����}��`;�rO����l�ܶ=ݍ��CK���}y�>ž/'޷���u��������}���� ������u���<�&8{z%��m�M�d����7�]�jq������뺮睈┈0��TK���I����&/@G㰁�w!��Z˷�9���$���nN���]ohH!�J�4"�?ް�빮o$�s�����M�M÷Ef�F3_�1�����%*->8�ۙ��_����yI>4�M�I!6�l�Z}I��`�5��t����sx8#�g�痴e�8���4�o4!^B"󗔒v]�E����I�~���������)���j�H�QU�V+Rm�u�'�w8�4�^�Vd2�Lji�[��}HPBG�	�҂W%ѣY6E���p-��9�����w�fUr��s.�����_�~����1ҚB(��Tt�`#���3���! +r�{wɃg>������%(I��x;NN&��(���$!�s4��(.W��rӒ��e*�>G�,�s=��l[҄�ϟ3�u���!�'?�	����m[f�vdi��<�Ȳ��(��P~����l��R�qTli�4B�H��N��P;�2�$<|�?���Fi���K~��_�X�m���" �:��)GGGt�a��:� �ƴ૞�(�$"%�UUa��� ZI$f|ĝ;�����7}�;�-��_~��=RJ�E���x��%��c�阢(br\�P�)�4�#��C�^�?9"Ԟ\S����ҩ��N���J9�>ziRႠm[����j��]}s���o�ìۊ�CN���ǻ�ҷ	�i��m�`3�{��>#c�ڮ,
��W������u�mG���b����=����u�$��置�WQxE�՗����D��y��l��ఀ��`���ݔf]?4ז�5�sӾo����C����^������T�c����=�UI>��Ԋ��d�!��c�wY��q��A]7[���J�{�>�߽{=���C	�ش��i)�B2��p|z������3\�b:�D�s��Z���,�$�d��	i��q�$��dJ�QJ1��1�1�ȯ���m���$Inݾ���9)��׬�E�\��'�0i��u�0�b�H-bU�ǹ���Eg	f�#L�P�/�ߔ�:�@�H�+�zMU�x��%Ip��Ջ��b���Q�Ѵ]��&���C=��M�L���q�r��z����9U��	(�ٔMU#� K��$ޢmKu~FUW(!���6-��TJ����X�k1ư\���Oʧ��5w'�?�����}���m2ʙ�G\�zI��9a>g�t�h��>M�7b5>I�R�&&��'dYFk;r������{���/�x���){�kIp��t¸�.A�[�g���4J-AF��Tx4-:4� >1��!��SMÁ�ӓ;�������c~���QEq|�1��j��r�X ��3$i���7i���"qz�������0c��1���a6.��pA T$�q^R7-Mm�>��y�o9B ���Q�MW�r�{�D!Ħ�从q�y�a�o�}����Q��y�rX7c�&�m}�{�Q��:��ns=�gd�hu�b;��؄�c|w8d�$9ܯ�BOחd�k�$�����Cֽ��!Ě�}��GȞO�M���؇#�φ>����[nb���XV��$n�چ1��ŷ����{<ܛ�Y�r*���A�*r��3ڳ�o�#z!�~���Kڄ���~o}���s��oR��f�췡�W��i7ﲧ
`��<���/.1��ރ;dE���*[S��xBQh�	M�	�u��|ɱ���1k!����h&�	J).//�s|��p��ׯh//Apxx�d<&O��,ѸeMhB݀�"�� �ƻ(�����KE�ԅ�x�Ak�I�I�Rf���,�Z%�J�!%�K�O|�	YJ2�'5�Z�'6
c�!�H)MCoL�V+^�~��j�R�<-�M���ֻ(I�Z��5�Ʉq1A��c�k�ׯ�(��S�밾#t%��h��$�C�VdZ3�N�ۆ�<��_��|��ܾ}
����C�I���n�ӄɸ`6���u%���v$E�%A��q��]M/�m�.�C�$��*ڳ3n�cu�p||���9W�,�s�VYN�4��e[���	I����s8h�РS��`�E(M����y��9��y̓�O����𽏿����i]�֒��Cf���a�Z��PIL��L^�9<>b:���_R�%o�^����Ȃ�,�8Z���&�q<M�jyE�ed�<e�F�� PR�8�Ơt"�n�Mc{%�u,����濿�r�1��I�۾u����}�!�/��z�Į�a���j�����ro6�}@��J��e˗e�V3^���qa�߄6d�`6,�>"��j]d�"v�(/����^_�#Mm���K��;;(��,������77����4�a';|���[psӖͼb�!��a�&�k|�����h<A[	\T5�'w��������ů��5p�.�zH�K|h}����M!�w݋��~;�&®���\b�!�6��}����%Zk�N�8�}���s^-��F�&ы����!���5i6�0%�4/PAm��m���O��0;�������JJ�V��zQ�)�5f�*�zO�*&���]h��a���� Z_�dh����ݩ�Z��B��:���ض�r���C��c�_
VmK�u���	�#�'����	������4OX.����8�*�EAVL(����moP��K�9F*�"%ϋ���6�^�b��)��W5�J)�Jct
2�&��`Ҍ�jIq�S 2�FH	��������b�0�h!9���\�ueW1�9 ZFr��r��gz:��vtVQ:��k�=���$��s�4!�d:�������/�����X�1�)+��L]��Z��H�
�u$n鼣�,���'�r����[���iJ�����)������_�Fk��&���q�>��(IWV1YJDȽ�֑A�傤�ԩ�IO6�կ:�шP/`<AyC�Z�UKU�@�&)B��ʋw��m��.E��-oc3����mq��ؙ�[z��\2޵����\؜۶ݗ}ۊ~��W[ivʓv�}�5%$ND#�����{&Vٯ���~��Q?�ߗ>�/D�.��j���!"cf�\$�RCΓ���z� ���D���}��A�G3��{�)�l��Ds��ֆ��0�!�-�n���SxL�m�,V]˦��z����������ls������m=���Z�g�!��߇���^�M���OT,��(�QPj�e�����7o�+����d�[\��+�k�:G�y����Y���Aд�oc�#��C�<���	�y��!�''��%uY�Z-��2R�:ҧ*E�q�Ҟ�X�n{!)�ab���2VQHI'T���!MD,�i�N�r�$�1FP�kV˒�9Nf����:�ItB��i�H�3r�IA���	2&쭗+�V!LB��#����/���z���|�x<"˲�Hr����)_�b���T�teM�	�iN1�D�А9��[|5��AQl⋓ɔ�G�4͙�g��3�T���kKڦ�UM4D|@���N�ѹ��u�r�0�:�R��,�:ZӍ�$� ��� MR�ܹC��^�1�U��ʖQkY_^!�E�v���~��Q[�u��v���e��0t�)V�    IDATԫ5��h�d�!Uܿ���?�=�חdY���C����rCۛ�4
4I��a,%
���ǣ��|����`t�˝���8�P5���������9�����P���eK��d���P�Ȁ�z�}����ؗG��o��/�C�3�n���Iᯓ�v�I�v�{k��y݉u�u�>��D:�e���7���uK)A�ػ�{�<�k�P��F�4/�m7e��=��@<tŋIG�eu7��0B\ȵ�K��_罭���mow{�a����1x�7��7B�������m���gehȳ�����0�b�3�m+�ok�nwt��t��}��
�ws"J�;!��HJk�Rt>f^I�7���hi0H.Ηd�C�|����e�!��d�����s$�1���^-���&c���[�o��	u����#l���cͼ�$I�d2�k[ڪ���_��F�pB2��&1S���#�g ��su��:G���b�ib�i)c��Ri�by������g��?|�yLȺZ��Ĭ*�UE������<Az����u�Q��v��#�����H'S~�٧ܽs;��W0�2�7x�Z ��-׸�"E ��{$ڶC�)eL$KS��tm�z1���������k�߿�l6�EHD���۷o3�3�����(MU�8"ݩ2H��@x�4�͂P(m	�c�ǫ�\w��\]]��)�����<R
��:�֜���&��\��$�X���]�)E�e�����:I�2E�$h��|K״4~����ׯh�g6s<;@	&�)�����UUqpp��Zg�	���$f6�ͳ�v�`2��e)��
�%x�G�#F?%9:�6L�9msN��V�[�<1d�$ֶ�����rd��]���~��m���m�s�����W�h�m9�/���X�[sm>�O &v��m�'7I������)�gI��c�և���W���w���R��2`���F���"��������ִ(0I�k�Ϋ]�bk��,A�^ J�V=�gd��(@�MK[D��4fM7.�[G2x|!�B��.��(��@�)��8�1Б��x��Z�!�IA�����Nb�G�\��0�����,Z��w�S�$0Bc����B DB۶[FI�F/r+� v_!^+Z�]kl��β�~!�xݦ\do��M��6�2
����8��},8!h)���^����b��ܯ�=G$��~�CNO)Nf\5�,�t������> �j��s�x޼�w�w�K��EP���u��]�$ϰ�%Uǔz���(�2�w}p���1�q��%xM�& s��c��!�c�ҏ��y�ےW�n���=v
�m;rmh뎟��/���:�^Y
��ghj�j�x|ux��L>"	]t�Z��Y+�?��� ��Oh��5��$��ۏ����ڲ����!��m./ϙLcރJh_�3�,���_}MB d��T�`B�sy:�x��7�ɉ�4^�9�"Q�D�~}ƃ���IA Y��x�2�I�D(�����bI9:��j�v�T�^�!:M�@۴\6�j��A�L�N��\�q8��zh=W)AA�6t��r��cmK:�`���>C/���m�]��%��]B-A{����G8_/��HFb"X5А��V[���c����_��r~�r5'�!�c���8g�'�U���B�UK�Z�M'�㴘R��r���:{�ů����`2;��	֋ i2�1+?�$��������"K/�B�ɐ ��?�=[��1�x�����>gc�H��m>��1~o+�M�����R*6��↡z4W���y7,��ʷU�Q!��+N%�n�	�Z�z)�6�BFpA���B�Q��X�HLA>!�������F����$:�x��#1)�� 2">4��b�c��(�/�����$:��8,JG���asѷ.�N����O�u���v���D�Ǹ�R
#�xZ���mI���A!���m,�0���Kѽ{��Y�nV�)CS��c'aF�y�9	\/]2�����:�"����&Cx�&T�m+�l#�J$R��k0�/QrB�ކF��z(K�T %p���o�Z\1��ǁR�,����ގ����g���P\M�g~!���$d:B�*OhR#1�̕#��z9gu���49���xF�Kj�^�E26$I4�.�5+������#�޼�7��s���!�xʓ�:��ǯ�����ł�����������5a�"xK���o��$JEjR�q5�p�j���3\:e�r΃���+8�*>��'�V���H����)�k��13	�{�U�AQ���Ղ"�qp�@�+P*Aj�&r�+��FaRE��dF�r䣂��QG��,K�D�cE�J"����D�>����	��[$J��1Z��{�+�2��88>�d�`�R�rYKD�h=̒C�O�y-�<�j�S�S$6%t������ф����<��N�Zb�L�@'\��N�L9=:F����\�v$��0s��;"���f|�A1�|JZVh!18�*�/i����'��D�ljF�";:�r�ڣ���*\�c�t��@�7)�?EҾ/D����GA��<�Aan��.�5�e��v��M2x�q�rm��{��l˳�a�����.�PR@耔*"!v'���=�LD�n�j�T����N@gZk\���r��|�]���:�,Ù��\��[b����O��q�f��V��(�6�O;(�
��'$�>o����R\g�{�6 D�9�닼��/\��w�Vl�&(��u�;�J~���m�L�P�����Kn�e\_�w��c0.�w�� �*{��o6���1��	� E�������F�y�%�Qk)il����ӯ��uh)���T%�]����˗�&9�zI��/�8s��>hC:@x�Q}WD��<m]"���.�\�xF��K+Ń�O������q��Y�� ��l�H��>��,�
���Z���3�7g<��JiB�7�g|�������o��Y�H�C�����5�o^��N���D$S�����Z:�w\^]��W_r�J���f���g���$���	E��@��;��*������J�p���/�KD8<Nx��P_u���[P� ��I�h���M4�Y�ݿǽ���]�Z���^�)�y\�b�.6-�,�|��/H�	�(�:.��q3xt��d9��ʁ��5���TٽC�q2��� t. �ݗV�Q��h�I<��_G����r��8�b]@�)F	�b�2)�Y�$� �傧/�~�fqx����;p�OT�>f����Ay���_���K�7g<:fr|D]$X�b�x�Gwi�a��S^]�'Sm8��b9_E�o����>�
l��=Y7�m������a�����C����{[ކ+���m��_>���5���6�\�A)hi�\����=Q�.��l\�>�iv����%b�E�	�o]�������N��<8�/�#D�s��CBƄ� w�C�o�]rw}�Ǽ�ɷ�����>{{(�=\o�ݹ��-���`��oj42����=��x[e_��|dV�6^��F�vH�x˰�Y��/˶A�������ێ1�ܶ1�>�����⎽轈IzC=�(���漫�-�{C(J��`�d\5U����g<���mp�X2��*�x��MB�h-)˒�e��r�V	��IV��m*ʫ�ؓ]+$1�C+u]R��;Fi��r�.k�r��?�1��c~������S�S��	!����w�S�g�x����
S@Y̊)6�S��ri�
d��H�� �h*T2�����������#����J�X7�F{f�B�R/+.__p�:���oh..������!DB�4M	A�G)M6*(�1�;�X:7���>��	���m��C�"�B���&�9Y2��k��Ƶ\�yC+5�IQ���V�,�� 2f�7MË�8�KLș�?J1�	����IB�Ev��M���"(^X�\�eN�Y�6EH��r�ղ�2c�ke���(�X��Q�9�r���U1��ŏ���gt�>¸(�E�
��`��s�^a�*Aw�juA�����_���k��.m���6H!�������Z�Le��Ws�5���[��O�Y�>�NӇ����Fҝ��kdo[�2`[�_�A���<��6*	���2���{�2&��A�D�Im]���-�8*�Xn3�=B�I���bXV���P�o��P4����s���s�<�*&n��qЛR��⾨�Z����]���ch7��{�����~l
��2�ݲ��������>�\��|�����޷�Z6�l=�C�ǘT�	B��9i����.�k������U������!��o�_+�}s?>��x����$z�Ѫ�C�����r+��J≙�^t()1Jcm�RO@'�b<�K��Ҡg#~�=���#:JZ
��P�"���,��eUR�5A
NO�T��+tخ�[.��CH�!�� 
!�&.J��Ʈ-���j���gT]ë�/�{�_K���tB^��U����tM���lY]\2^���#1���=�k��KKp6z���,?����c����p�/?�F"��D*TPdF#�buuI�\��W�W�늯���,�,���m�� H0$��N�&-��bmZ���������b<���Ճ��u��DH�x�x�ik�m�ǚn�P�F�ۆ��JHo�{AH�,I)d�/r��|���ܻs$te�CJ����A"B��CIhR���[Z!b����Β����8���5��Qׁ���== {�1w~Ř���r��jR��M@A�Z���+�<}���g̿�=����W/�0�4�9�����/��ٿ�56�;�%�w�W�I��v��Hڲ��+��;���o���˙�Go��~8s8�FF������S�?<\��#�QYú�v�nR�Q6��	Bzֺ��,���$*x���<%D�'�T�8$�$
b�F��
ѷڎK�Gd��7o��PK?���g�����O��=P����!*�l���(b��З���^/�9G��Dl����>n�[oǠ�%��gȜ�6��񶡯mE+y��4K�1��d�h���e���7s�]$b[y��܇����7����>6�^ ��n��sܰM3�"6B��H\�!�@IA��]��<���u��}��\b�g������equ�o8��3�W�y�U�d<��~�gT�W|A��X����J��1Hs����LF�3-9g��}��g_r7�|z��k��5YH&9��Ԧc�l#����V���[_aۊq�EOZ��;�+vT�#�F"�B����������G?��Lh�uM�z�UU�|�~���!��
�>��]��~��Q��\�$:h�M��Y,iu�5T��;�DRpt���Zk� I�(��d:��Mf��.�㜲}�W
JU[ruu��i�o�6�]pU�^.i����l���f|�/���d�] -Ftx�շ�EƊ!$h�+�0̲��>yW˘��@�%A������W�&��0��g?���T��`�FB���i-	��4̯.隆�|���9m�p"c��,�9�uˤ�1���(�KV�^�t�%ڃ��H������ڣ�����^.�w���:&�N�f�7��������}�>7)q����`�����Hg[��@�����0�ӈ߄�"v;�:b���bֻ}�9z��9�-b�!�hG��E�#�X>K�9L�]�%�b�0��b�~n�)ۊ��q���ܞHY����AV��������p۪���� ׍߅��<@��Ћs��b��7)��I�9�'�_|��Aoy�.�&��&w3���oo��V�ֱ!K�tΡd,�X�VTU�v~�BD���ʆw@����a���f����/�ݚo i`s�����\�>��"]�M�E��;���1}�uZ��46��%b[R!J*L�m-�ƫ@W��������3��9�B�Xpvy�N3&E�����I�U�z:�ʯi�|ó��j���22�]Y����BNF}�d�)���l%$!8D��z�9wR����t����$���P�	��j�(W��c�n�$�i[b}��&!�	ע~Ou.%^x��zq�ٯ��'�IY��_��˧�pUGf<�rAu�[��I���P)�)��V_Isy�)��9&��M�ID[���Q2���&>��g4�g�_"ˊz�R��qԈ��bEY�H�0;>���]�ƅ��Wg��7���
�z�"�@����"&P���tMK�e$t�U���/�� �u���b}�d�^���L�(�r�(7L2Iv:����+LU!��6�ѥ�gw>�]���*v-���q*He������Y��ʒ������[�y���tm�J3yx��G�G��_S��y1b:9@%� �ф���Y+Ȕbv4�]W����i{�I��<�[+"����gf�}yHI�E�K�ӂ�����l=0$A"��_��I�DQ<����twUfF��Ê�Yݛ�scvWUf�eEĺ_)I����������lm)��l���5��.�-�ն�]��|�E;i��N���^ͻ��јJ�m���j�EBX�����q�㠨�Z�N�ι�̈e�f��̗d	sZZ���=���"m��]� 7F3(��y5������3��Kf�N)@�/�r��W��	13kq�%�2uJ��k7`�R���8oCA��HsS�������i���w�#I;j��q�)���o��_��wk]�W��$jި��V�����۾)i��2v��O��	7��$I�{�Ȃ�Ւ���D�����0����x������wࠎ~��fN����;��s\�������D����*�����7r��02#L�eL�O;�m�rf=E���'�?���?�W�x�G\�Y�'��cY4� K���7�w8O���gx	�cN���x7b�ϕ������� ,������?���g���CD0}|�џ������9?��8 ,�9�1޿Eb�?��-dN��x�#E��*{<���"�A 
�y�=�̈��ӟ���?��ӟ����'\�y��9 ���������k��޿���Aw�8���/0���8�`�.ϏZ���c�4��FHN��٩#0"��?��7��~	�o~�3,��7O�1aI7�q<8=�Ϗ����q�s.�r�4:�yz�0
�O3��� |�?���w��3�������>���8� I���#>�;�>=�-	�޽���=><}����_�~�[��w���i������ރO�?A�Rw8�pw-�$�WBߩ����N�iͤ���%���7�i�k���-��I�1\%HC�NWm�ў�f���K�=��L�@T��J�[�'5���eL� �V�t9oFJH�ih��.˘�w?7�Kq���G��쨽�)���CHO8����U_K�z�Ym^�]'�:�,@�:0@ `n@�* K fD$L�x��R�	S�wf*y�	g0�� ��(�	�$�s� �9ǵ;�4�$'@�֫��b6=0�5��s�C6s��U:8����Q���!��=A����&r�Jz�v|m!�k�!��2�eYmj{'A�Á�M�};@�L�u�(s�1.+Θ�a	2�>�5	�b��p�gZ�vLZ\��i���;�|�<��A!�sҜqHH��:���;i"�9��~ƴ���������4����?`81���Π%!� v�������Sē����p:b�#�9���]���!'���㟞��t�p�HS���CX�oO\R���4�����x>c�R��?�K	��~�-DwI@4kd�'KL���Oa�s�i9c	xx�����~��,�'~���Ņ���Y��F�8`>���՗��_�SD�fa<�z�+��sHKB�ɗx�����Y"�G<?���ޛ<x�7�5^��x��������8L_�������q�`�    IDATDhiV7b`�DSڊ``��2���$ͧ�\p7:�w�8c�܇� ������-N!!�n�Ñ��#Nw���3����������$|���a1d/|>��b�3�$|L	?�iuO�K���xT�9�-M8,���c:�śOO`D��xϸ����������t�������[�+u����֒=��P�&.W�Y;���/d��9薄�F$�I]��i�T�ݴD���ύ��c>���\�j:��L#IE��v��89,�e��s 7d�z�Ï�4��Ai!{�c�PN�j�#��8<��K1K'��3:����iZ X�v	&��\�1%$h� �c���hIHf �� ~��19uQ+� K뒈����:��^`L��B��0<��gl����e��d�!sU�M)�(l�v�	�]ac�^ٙP����J����bT�8c]�ɤ�-i{���߷��&�)0�c�~�40[��.�q�����*���NE�^����= ��y���=��?�ܽ��4�\"����r��(�u�dH�i�����#.���<����;\>}���.>��{N�� �0�.x���3��#�����✃�pw| �d	2C�X����8@�#���g�ő2��<�/���0�0�>�X�`qG��a�'�55�HJ�S�)8�$�!H΃�4!�l���z5h��N1��3<{0�a�cF�' &�������gE��I0x��#�5ϐ`	#jH'� �D|��{���㋿�| .@ѿw��>��go�$a�	�'xbܟ�d$M"X��)@b��y��a��S�gwGE��7�H���HQ��e�8L#<? qD�K��O.��x���(#�|����x Ma�T��g�lr����Y����;8:"��^0a�	�c�������Ai�u蜢��)���>-�y�u�R����\�&��~�*̌��qǖ�U����E���ϫ�6-�d:`�/�
�[�PՄ�˾����I,TLF��1��	�&F��r

3dJ+�8nјg�A �b �����z�� $!�0@YIMPb�@�io�����sNP7>���}VگC��y�W_,²═�P�j���U�-2�r��T�Wpm��-��0��Ll%������*�Ԡe֙���6P�#���qa�SZ�p7�<��xA�$��w�>~���&.��)��1_&�I9��4��"�����w�0,���	�_�>��5�޿�7q�#�?j(V���#������t��y����X4T0-bvF��`�\ 1�#$�8�p9k��{���oqa���A3qyvHN�����x����� ~���&I���5]!x^���Q�R^JP�R�|8�oޜ��Q�����f�0R��#c�>.	��3\x�Ek�NC�8��0��P��zG,H���y���	�� 8?�qw<�SX���>�/X�q�h��� �Ys�3g�d*Z5?�C��,$,DX&ͯt.�Y0���8_f�%�$=~BDB�DD�x
�}�xN��3bx�p������J��|���>̇D��)��Ì�̘p�0���j9jFQC�j�$�М��b����j}�&�k"c*��\[��ιή��X��U�������{�3�KW��K_� �������c�ڄr�{D�!R���#�9����le�}�V����(}��m������%P���R3���^�� e6&{H�3s.,����aU8�WB�۷��Ò8bH#U�Pi�6Χ�"��|�D�2�7��櫍׎��`���r����HW�����F��گ�{ێI���o�ֵw@�X��ŞwW5�2G�R�$��<�,)j��x8|�/�������hiN�y� ��b�7ˇLhU�9 �K֜Di���9�xAJ.��B�����1\��c ��7~�������s5&K���A�2/i��zYT���AD�.��@�	��gSB�פB\� :��[�w����7p'��˥�}n�"�eA��r]��c�c D��#$A �}"|�뿎�8""�NX(��p�w��⯽{ ŀ��3ށ�V�\.�������"��1�~y��|�a�4�����w������O�����	�S�H���[x|��iZ@�L�l~���劈������3�qħ�!�8�N��7�b��p��_��8|��  �Gw���	o�#���� O�L�0��r���/0�s�pv>��Is��/�<ň���iSU�#�8��GXH@�^4�_�,��N\�۪�۳�2�A�_��W��$��}���3�l1 Tx%�>HY�k��U���2��"ش�7r����	ժ6YVE�PyĴ^Z��(f�%M,V��\��_��Qq��n�c�κ�5�n�FW���IɌ�7�w�!��Ad7�H�	Q8���d))f��Aĥ�}J14S����T-Յ�q���s#68_?s�'����_���K�&��s_UK���'�n�v��*��Gw	�e��#�a Q&���o 
!�wmo�[�n��L��?S���J��y��������S�8vx��i���%V�ȌA%����}��d�D�"��#�p8`�G9���q��O���>;y�ww �~	���|(c�8b�8%����)%8O �/¤y��q3���#�b,)���9������{?���BH'�{�r�yݗeAX4<Q���T	 ���{,1�H���	���������]���;ڇ �0�!�� �bv ���PB��R(ɟ\`i�8��o���'�1�9j5@����?��?��p�D<�q�f�x�p8 .$�D�iA��1��{�^ɉ���3�e��t��p@�Q��1><����G�@ q<@x���~���M��H���7x��q����1���A��B�tƒ��XLV�j����_��/�B���Q��R�C�@�!�����"�"��'坥_�9Xd�wW��j|)��{�����8�����;g�ջ�@!%t1������W�%9�H��آwL3R5�V���J8�d�hW�L������57KբR_Kc	)]�:��e[zu��R���l�f�5�Ħ3�8TG�ZuҪ�׋U)Z�A����WV�|�}e6pC�l���!Q�m��J<��{V'�F�o��~×�H�Z�J�\k�J�G�G��_��wZn�J5���;�I?�0����~�����o�M|�i����c�9�2�_E�VM��0�
��\f�n��b�?�8&����8���$��4��9� V;����D9G 	�1�˄�P���|�5�����x��=���k��woqd-Y�< �3FfĴ`�1����I& �(:~����u�i=�� %#�r ��N'Lˌ���˄�<iXZX���'���p�w9�w F�ڡĚ&�	C>���X;E�2<\�\��̔f�֯�i�='�8#� Y�����pt-W�a�?��I�٦�3�`�� ���a�����q7�7��!x�{�� �����sZ��㞀a�0f��흞_�z��)�K�jSi!�O�7�p�,x��"�c���.%p.nb��$��$�p#U��{޼�;Z֟�V�����9�
�������}ۮ搫��]�����o��綮�1آ���<�����ibr���\m�dH}3\�d�Z�R}ۻ��iVW�CB��ojO$㍬y���>�A$��n�Z�+���YK�B*�,�}�Y���#CJ-dfn��׶-QkMkTj���K���R�r>��a����4�]P��[l�q�__��)�#��z�8s����V4����NvP{M@�����k�DQ$��AmET r�ԶZB��8�������_�����,�p'���' Ha �SQr��I�0e8�	�8*r)��t|�D�8p!A"p�D"�� sN|���0�!K	�!o���3������e�hy����b�|�����{�C"D8�#FD�(x;j.��7""b^���a��+D�j���!���E�B�~f�?�#�3fGHiƈ�Ӊ � vS�G��#�( �H���h�����i���0�	�D���9�y��0F/1!,3N<`$ ������XsM$�H ��/�!�v�` ���a>gs��w�)������91с'���B��A�o0��g͎�� ��t $��E���k�$�pT��Xv�3A�g$��wpiFHO�:p�=\�`����!��ֺ��< ���Z�`�n��Y滭��֜�����o\[c��5�t�v�6��hoi�9��WB���5sa~!�t�c$�����*�S�
{�9y��B�63{�����E�Иo3SVF& ��*^��_#R	� k
�g^���1B��ږy�lR���R�z��gh] M���"���w��I��r{H�Epz�^&�WDX����xW| Ri#%e_t���s�)l�X�!���Mء�R��V3����������^RwY�!������զn�(pl���m� ��ob9��^?cܖ���������O~�ʂww���Og�O�hl��A��$�%'��t�UER6���p�D�p�����ǀ)��W����0b�k7z�-Q��P9�v�����ԓ��g|��=bZ���#��?��9����a�>xC�	�OF?������	A<������ו�J�<5�*jIi�!<�� J���x�;�0�wAp-l4�Q��,X��K����z�� ό�g�g^Wa�#>L����#��OO�@1�Q��5���p�q�a8��;\VS[?�����|? ��o�q��yƃA�D`�9^ ��9��~����IB��8#��1Og�Q�M@4����Dn�Y>]h�Q���`6�d�"'���������ǿ�{@�@�LR��nђ1�v��؎n��W�g�Mś�� rMo]/᭾o�_��K*�7#u�����䃴;j��D��HylY�`3l��(�ˏ9�L��	̔����YFJ1��6�LL_k`}v*�=�)��A)3#��)Ja��ˎ?��a�!R%~]܀�|�\�euc$0i�h����\��b*�[s ������y�TH3F ��!|@
�q�w���Sop��F1��I�\��:\/�f�X�9��)"I $��")�%?�r
ږs�$����j~ƅ��x�nQ�)�u��۸�ҎC����E��Q�� [�-�M�,QՖ��0�}f����rZcfh�W-������|z��陰����$Eu|��5�44�,�rݞ�y�1C@�!x�sX� �>�x(s"�:��$���3�M%��?��N��W��go0=?��O
?A.J�Dc�L7+��13�-�o58˜�Ú����y	 x�\
�p���m��t���uȒ�ؾ $Ԫ�����Hf�ؐ��Ybe��;,Q%u�=�9$� ��˂�B��9��3~u�x�>��f�����ph�nR��.dfD	ڧ��.���y� $�uO�E3g���8�y���ii�^����p8տ�T�c��q��c�ڳ2��8�/�,G���������ÿ�g�3��C @�<��pQ��)
�U��ӖY��'��}�[Y�6 4�C�R�t'9�{�����54mE���$0&]6�e��iR o��%1�����	'�oW&�6���b�|-�$���N�x{u��$���	�)���C��;@��hjmA��DBк�<��F��6u �UQ�I�L���B�A ���&B`e��%�=a�ꎫ�����}��s"�B<��DŦ�.x���5^Ir�qe`�"FJ�T7#�a��$�vfCH %���g�s���kmq@Äp�6�`�LغzUP�h}��k_��2Q[;�ݶ��%���k��+8����1���߾-�~Cn�f��K�T�L���V���!�3�s�h^琰��Q@(�"���t;Ĥ�����p�"��x*�&�Wr� �9=��s�I?����� �S.���M.e髅�jv�QI�0�V"9_r\�ռCZ�Br���o`VLbU�ί��y�j|)&B5h�L�pCYԁN�CX2��4Z�������=e��$�2�LlNK,�.�7��9��PP&��#��}.�	���Ã{����'�SO�����8G�шgfHK���sZ����!(���dE�%(2�B��q\���>G��,��BEJr�!�KY��w�h�Αp8��D���a�\�x;ϐ�P�Lp5|2��	��%�ר���W+o�����wKh��o}���K�-�F�u�`�,�o��!q9����Si����|�*�g;*x֚-F��?jL�[}y�9��)��%�=qi�ը"�T�w�R@�P� �B4�!d��4��Bݰ�1��iӍ
����b9�m��v��Y�v������b*{���@����i^�N>��s�����_�iR��oȫ#�/�}���y��[�)����Ś�DR�Az�V̀dv��)?� �����\H4�>s\ $�<���# ��bx�V��
A5-�=�kZ�&�3���̣:eZ�'@b�9�z�F�bO��Q^q@��Ț'.p`��\�BA�4!8�!Þ��,�ř���Q��Zå0O�sn�JXT�-<�us�_Զ�"�S�����G�o����ő��3=��x@r��:�Y���L��i�PR�ƨ�"?9Cg���(�I5n/`���Л� a�P^+��ܥJ��6ˮ� pxRU뜫$
0Bs7Lw�b{�3v#����".�!=1�zcOD�p���p������O�<��T�j����f/ `�P�_M� @�I��I���ā��>�aulkx������t�zԐJ�'	��t�1zf�T��%B[��k�`�[ KE9�PUm�:9����`V"���^�hr	MV�@����Z"����Eƍg�靺�[ꩭ{�C�=7ߑd.��C]�v�]�9D~�_~�=��E�/Kq�j���xw�VB���ܸ̇���~ccD:Dj�)E�٦2��H�*�uc:�Tǃ�;�|\�J�N��'l�OR����Tj��KcG��Q�*Xg�L�,(ڰ���tJ1_E��f @�<��Z��R&|ɘ�kC��T�ȹjH�A	�\���1��nad���s�xí$�!��#PZ0���S �4a F�O?�	bx���	�o/Z8. '8Re���%'�����H	�K�nQ���9fPPXIDJ�ĕ.�t�����Id���UƸ���HH�D�13�Z��9�f��c+
�'��}��VJ�>/]/I�mx�k��^�eBO?�"�r���Zl�?Be������+l
�"4���Z���p����EF ��6���4S�����4����i�.�Z׆����lC4�7� {�#�T�j��:6K��S���,\�k={>f������!�V����e��j�7��S�f;����9��>��+ ��s�C�x��5�Yeg^{��'�E{�s��)��2u�& �ĤU��k"\�l{C��F��ڣ�Ӱ�����-�<��*b �g5d�,�Ըn#$3̨���ٺ��SL(���'��%Rg�b� @q.�)����d����N�l:�$�X3 L����r�8���l�sv����H�:�v�4�f٧ X>����2���<~���<�D9duI�� ��&숨a��ƅ��L�
J�!;�Ңf
Q�fE��<2(�c�1ER�]��8�#L�џm%$�FP�F�i��4�TM	(D��VDr8��Z�g��7�h���*�;S{����~[���B�>}���r~_��ָ{&��{��[8�]�L�Yi�]��7�(�9Dj�눊I���/o�@�.pQ'6d?�W,� ���Ku�q��� !��1@�kr�_�Fs���5x    IDAT�8���Tg4�D��iI>�x(��H ��kg�������o\��T}���2��;=���pK ��e	`�������D��ժ��q��@7|9��vTb&�T$��!�,�F�H���$ i"q$G�vξ%ˌ(#�Q5�ˁr
��$߱���V?e�E��jNpy ��"�,9'm�H�MU�g�WJ �\�ф���'U��8�f���؛^��q~. vSB�Wn�v %�H�iQ6|2(��<:uh�.m��12D<�0;P���RD �&��A��9�X���qɪr3�^i5���MG]���dF�%���E��j�W�&�3�݁�GBŅ@k�8�t^���"��@59�P޻F
Q7M�}��ք�W�e}�_:�{����%�{8�}�׌��W���m�jx�m /|�6 ��+h�w�tM��g+�����zCu>[��>q��j���
5ھ&��^�m-C��I��'��R�]���*��,\]�J���+
&#x)��i1E�ޙ}Dm�		QD���E�*�(	H��HM����X4D������^���9�����n��&�\��;]N�|	�9��s���`�t}�Z��U�m3�ת������X2|Km�XL� Nӿ�'�;�����Cv'.3�I���
s��q�`�1��iF�¹�,+�1�*�&�I�4�xe�%�� �!��ڢMIZ$��2�\���&�����3�vO��}����{�,��By%�Hꉀ(��� �+g�l�@� q��(a<�ڒE�~ Y���%b��c��i �)"�F�d�:��٬�L��1u� ZF��2H��l�ET��hx Wy pf L]o̺'(#�0h�������e�I��Ĉ�|�j�;�F�AXI�7��^����J���}�0�_����J�߹z|�]�u����ȁ�F1�s�e��w���zC3j4e:�m�8A�4��p^'@3g�����楓-}J	LL�яW���'Z½B��ip�S�4����4}��;�č�3�`U"�II%8?ZdTJ6��4���D 	B�L�c_q��el��ݷ�ګ�Ѫ�,b!�<�NѸ��$"��{t�w'8",�F	����=�x���K\�K�e.l>��&��~C�!�K�$�=�;N��K{��TG\��/�|���X�w��XҲF&��F�旒��$ ��S��H�L_��TZN��Q��S����<��@Prl;Pv&������,hf��HMe.�L�3�L�D9����P?��m��wS�Em�G���� �T���!�0��cD
����%���xG�	���'N�K��\�r�s
c���K n�/�K	��	V� ��A`�%��LZ��l���^��$��=H΋�A�#fx�u<�h!$J#N4��N� ��c�,���#�{gvS��X�n�<�U7�g n�{�֙~���.��U�л[��f8�p�e?]�+\�~+�W���|W��+��-A�g��s�D]	n0V ���0 1���8Y���
1yD���}�� �8 ��9
QՀ�ޘZ�I�D�#(&��D���		3Z�R����S�Lu�� �W�v��:�0 �?F�J�"m�R�:iT�ysǸT)I8#��{�jv4[,�  '�Q�z|�-Q	�m���ڈ�E/%�[h��fm����"�	Tl�>3Vŉ/ŢY�%M��*KH����L���@����Y����ps�cM�z<B��eZ0����oచe"**ͷ�la���S]o���{!��|B��y՝��_&A�KS%�l"�o��LfyL�5��m8f���J�s�u�Ga0Jl0ҊL`�$��#�0�qY�<��h�8iA"DH�c��	2xܿ��{f��7p��#<{�G��a���$"�>��f�+�$A�w�+.՘����ȅiQ�y&29 k���`MÛQb�H�97f@��x)��x.kvZ0'�����H^��c�#0�mJ��#��fUhi~ܹ��Ê�#�2^)U�)�[ʛH]8jq��f�.l��A"��Y�v>D%ĸ7!�U�Ͷ	�\a�L�XZ�D"��f�y�-�H���IK�OXb���$A5�M+]�sZZ���M	D'�����(F '/1�'�iZf$��e��o;\�����C��J�U����j{bh��k�e�s��^Tb�֜S��k�wb�����%�#[	:��U��mmq��}��������Rvz��kg,�bi�@���k.֐2e.2�&�q�����uj�RI�
��\[��y����s��0��j���M��4;��`���	r1ǀ���Ln~8��?!F�9j����)X:�~?��+t9Jt3�]��vm����_���7��U��u�}4�����.[E/y(�+������hf��k��{�E+������랬�O[�k�GQ�+8�%�����7�T�V��Y�i^;.�?��S�^ڨ�ߒƍ��ڴ�?]������B�-�@X���+M���iH۷}ޢ+e}�^�\S֢����o�kFo�#�+���_kFU"��gk���m�ýkS�׉)�ȕeK2�H6�[�9��5�I,���сe]֯�d��������~��L�J�mۻbl:ΐp{�(U�`T�Lh�5���3���v��1,��'fo\?ۏ�x��P���9��n�`�}�>i��X�Yq ��K�Su\���Èӻ|��[�% ��%�kג�V G��^DU����௉�6�k%����}����${8o��&#P���9��ؚ��N��X��c�Kf�H�k����sLӄ���
�	?`ȹ��3P�Iq"��k����/��3�<Gk�[t���3:��(;{�Jf+���M�������5�����:fƎ�mٶi�;0}��=�l���7�o�[�o����#�z��>�h�Ιٺo����Z�����}u�}���bBnk�1�٘Yv��}&j5�ܕ1ƪ)�"�&K)��/���{U�DU	U��JͼT���^�_]��Vm�8n�-P對�����9�~��[��o�T�#B�S��}��.�H��ڻ.�� iU�X����,�عv�nu&�!����=���!�.'lR��.���[22"}'���È),��5}���<� <s�j���T\K �I��HsS"�L���H�[�ے8���uf�zM���N�*��c��P<���{��M����g�vA�q�b����epG<��p�,n��J���-6���I���F7�+�^�{�j��U�{C�w����:��Dޮv�Z�so��˵'���=<�
^=��q�Ӹ��~K�oѨ[���ku�2�жH�a��c� u� ��E�T������}Z��,�a��^e��x�WV"���mr[7�fR����Y�.g���ت0�ƒ���ڴ���I������BNˏ�ͭmC������{!\à<��ƍ��F�n|�G�v���Ԇ�m�1��OY��r.�^�=�ǭ�='9�DJA�`�4�Hyw���X��O�<������\�8g!F�G$�C@��6o�_���dV�%�C��
һ�^�s��ZPh_�aha�kr������s-��M����(#�w�R�
q�J�B�騱Z3=�빰�������N~(`Z�f��"x�w\�m�L��o�1=�0�彊����m��XkF���l���ګ85���Y�1ۻ��J;�wy���[=��
����������D��k���i}��͒����C��gk����3���d�\��Ld&�W�~�=3���H�93���n|�̶d����ѵ����,�;����֡��[�l�=B��U�j����7�B�
.�Ն�\�"JE86vf@R���p) ����y�ﶙ��݌!�p%"pu�k�oj����s�-���T/�~�)�˭�\M:0cń��x������*2���qIu���b�������ie��!���>�um!Z�K�kR�#0)�n�lKVq�0�5ξ�������Y�kgW�c����N�3�Ow8�'��ݟ=L��������V���|��Zn�����yl���%8l���w-�e�\��o��/3�~{��_߻��2���|K8�jk�^���=5k%�3�!���* ��}#��F��tQ�� EP!��rBd*ɚ4\t�J�{�Sܼ�K�&sl7g�6��[ m%ւ\VR�@P������Ԏ�SZvD�����Yy {�鶆G�t�j�Vۀnn1D=�Jcڿ�	�<����]&0�M68A�l��4�J�^:�����.�Je����	snzm����M��v�I��ͯ!�Z�^D���y $HԪ�K?$��lk��G;�-��w�f��koo�[�`�
DZ�Ɍ$����&{���7]I�2%/f����E��͞X�	�@��͗�`>Ϻ��c�V\�qu���S� ��$�J.���X��/�^q�>3��)�x'K�VҴ�@��$�Nx8���]�Α���B��FKS�\��=ؘ�`�/[{z/Eo?���--JO��ƱG����c��^Y	g9�={��$6����a��/F����&�+p�Գ�u�o�ؘWkVj/o�0S���"����x��z�#n�m>k�WC������oἊ�^C4d��t�k�܎�Vϴ�����ځ��AN��^s�h1�c-u&̡`%��dD2�K�ÔD08��ϱ�T��(n�@t��#P��;��Yѱ&�Ii��׽���̼��$�/L���	X"���!r��n��؟W��״�A*��5��UU�ۚ1����=ig���we�j
\4�b�ۏ�~:з��� 	J6K;���<���wP"-HC��,J-���OU�b�R&ژl�W~C+����������y��ڙV6֠�_��
��'|ݰ&�J�K��It�\aZ�i������oO���c^��n��N��oMh��o�έ���D^D�O�[��V�o�P��� *Ny��J�:|����Ll���� >��!�N^Koq�tPX8C����$ $H�;�:�3�h�A(�*QI�h&BHN�H�Ej�*�N���sv�
�����f9�8��@���c.��ݷ�/�k1bL��t��1�=k%ܔR��E��m�bXԣֱ֪��#:>���Vps������J
97�,y���fVϱ�N�vX��T�ܳDF���J-&{R���}~�!�I�c���5���Ro�� �)��t
 q8�˰< �2">����]��2��c��k�<5}�u�o���!m+�bɣ�܊0�k�BVpk%Z
�"9�	�5$��~�{��h	�(�����*i`�X=o���0R]�#�pp^c��oa�98�%&|��xxx���>~�-��EM^�Br'@
)���Z��ے�^ ?1fDeB\�KN#[�
f�)yxLP)�{�3�U��?��T5/J1)*Bc� ����~*�� �Kj[��E?���&�ϖY����9�;�}x�-}��Pqzśh�'��fk�WnK�-� �Ť���3КÖk)�h�Jr���@�}(�V�̕+�i�ҧ�12�jt�T�"@�\�<�Z�>iN��I�Dps�%E{���0���UPN�镝&��	-UN�8��y+����I9a]�:��� -0�r���Ό�K�mF6A��aG�[k���b�M)僢)o9%�H��n?��M���Z��!��o�+x�7<��A��a�^���֖�����4
OJr�gH�H\%!��f��TYې��Tí��]:�t���e�7�l\�TiE9Z�M %;��|�;8à��Z͌���H���- }"�kK�nc�{�C���4��Ͼ��-���Uٻ^�خ$���G�0 P�*i{*��4�QJ	�˲"�$]ͭ�C����o΀Fh\�<���Q�ֶ�Pc�W�,���2��_����T�a~"�KP%���U�/�g?�-�_3����	y^��`�����Z�M���9��[I�z�-fhFŗ`~�~�i�K�ę�������RI�tm��/�r}����_�6���նs�mb������̶G�K_l�Y�{N՞i�fwn!���*�bN��l��l���/7�Pm�6��"�1�-���Y �*�[֤�gտ���ڜ��|��"���ۂ��j����>��5�)"�Jv)	b�����W�^�U�긚�9p'����"��q��������Q&��	.�Ĺq�!�m�8����e^"����~N���%��00aI	a�!9���Y/���~Dd��e{ƊM1k%� d��\�0�D0���] �+%K�H]��1ݬ��z�De��cD+���k@r��m�-S���w�a��k�y�8�1�ڻ[�e���OsSo�/���pd&%=oL��*�����TA\_�䶰]��-ӳ	�/�̕D����F0�~�hg���A�I�e�DEz�#��gC~�� ���~^��IϿ�~���yi�zK@��b�� ��5Q�Y�z[i*6kQ���ML� 6��AH��%85�Q[}ֿyV�R�E��9޺ZI��L)���Z�Q�]I�1	�*I��o\-���=��}m35m;���i�CL���ja�w�m���{[���b��j]���F����WTO�'��N@����r�v�l��Ǚ(��
k�gu|������+/����\��=%�k�X���j�E��i�Ԥ��׼S~k�
3�A���Kc{�Y�%���.���_��%h޺�=\M��<Z[��W�>6��^�K���%�)e�jm��J9�]�U��:�'��Bx�:3a_�hm�+�$�}���ZB 2U����
���&�jŒz���<Cr�M}�nJ2߅X���TY��⻧כ:��L�����J"G�`�c�����"O�=<�]���YP��v��� ��g�	U�6k"��U����deo>I���kf�|Շ�1��x�5U�=8�}ӂLt��~Kԁ�_�Dv/����ڿ6q�u�kA����#ZU�k��KgB�f)��ێA�R�1�'���)�*�L�(����iu��7���Tr+��U���6����]m�r�ޞ$eJlo:<cN5g�,��;Y�C5x]�Aa�# 0��6Mvc���޵��^sV�p�����{�k}o<[��-��?��Po��u���_�4۳)�D�r]�[�L��@�i��u�dᦥ�6�9�����)%חoqv��D�� 5g���F�-������k����%!�]C�54'tAF ;ia�T�}K��z��ey�$��kM{h_��.��-�-G����~����Hin�<D$�
+�f��%c�s��t�_8P{�`f$!P.FR�H�����w����KL��<�ᜇD�������o+T���aj۳�[��g{��ڷW����n����-��~^=���"��	0�:#�EH\.����J�ք[5?�3�)��Q�r�"D�$�*	>[�$�b,ZkA�:�[s�}���*�u��n?o	@��仌�}��L}������1m��vn���ψ�ë~n"?
O^ӎ)>X��qB"���w�5M�=s�R��x�=�n��0)nT�B��3Y��+���,	@�W ��B�0���]Y^"�g�0U��G־������;q�[Ȳo���_b6Jj[�lKD��µ��>Za3Kcv��-�Ҿ�&��g�eLO��9/���k�pK��w�q�=����=ưxKfR����Ͼ���3��5R �� �DO���q��/-�鋱��[�|��陃~/���1s�ߥJ�FN�v�[��y��FK?�\6@�@Tc����(Tdc��\�?���Im���b��q�A�|2�Dj!R�V�\MA��5�SG(^�o�=��z������{�ݗ��-�ն�������2�ޔ�����1�=�mkL{���q~A 4_(&�L�y��4����h|�x�o��:�3vw^�߷�R��JK�A8f�sp�R˥��`l@���O�%��%�Ԇ�u}�=ΰ=���yYJĚX���{���ܶޫ�P����u@�H����-Z����`�^�h<�E �i��6�R�T�v?W�]V|A^�k�{}�b���c4%��    IDAT�.h��6ʣ�Mu8����$�?��?�����	"�y�x<���l�PC�{����B�/!��Hǯ���O��-�.�h��_�o��u��Kr\�f�c$aY�_�#x��M�<��ߛ�La³���c����V�Z��I��b�P4g��<��'v/]��&^���Dq﹭w�q�bF_�S�W�C��^l�}�q��{篟�1s[W�=C��-)��*E�i˄_�����K�(�w�T�%͌(��DTߘ��{�`���w	a	 ��|G\m]Q<� ��	vaz^@1�tdHr�%��\ɱ����r� ���S���ℑ5n4�.�ΐ9�!-�?�4�yPլ$�@.��xP��M) ���s���UPl���Zը�iG�3
�m�ў'+C�`��	���g���~����%�=�&� �N��2 �Sӧ��-�]#��`g�&i{&Y��y�����^�;��6��\�V�' W�:�jw�vMO�H ;���G}��U5�N���-DJD�60���������""%�=�p5'#�-#�"�{��g|x����;�C��=��k>��
9��S���cj+�;�����Ƹ�D�'�q���e濓�@1y�KOM����r�;}�WK�â��� f���oNT��F
	�����1��l�9�p�*�)�[���%7߭~K]ۍ�M����WKd�p�V"5b��,�!H�i`k�r�ߞ�ԄX-�^Q�qk�֖s���L�4��WpIR�uN�DU;T���z,��sq�e8Va�3�0#ffQK��bZ�l�*� %@ڿ�1�P]9x\N�cf�*�iH�z��6
�s?JU�AA��߃G���o1��I�V�RJR bj��f�N'��Pu�6�8�j7DĤ�
�N�t����}׍S�P���ڔ��q��y��F'{o���[�z����+N�m�guZ��im�51J�.�����&��Lq�����.�#�s�W�;�!sҨj��0`"�>U��-U�i�[	�Zտ���M�n��i4?6��'�0��'x̸��|�~��'��9k<�����%�i��<�k�(�� "r�w�>4iU�m��v?�G;���1m��&3~���I�&��:�m���v�r��=����]+uB�q�/18���?��D �Ľx����3��d��x	V-�(���p�m&;Id�⚑�z�վ�a'�4s^�ʗݍ1b�3��6�Ƭ8��` �b��Hиk�����X��afx��2�NtI�bF��<א����y�o���o��z�w����Y�>��j��z��hF��l�9�����s�-�i	}oϵ�����ת���6�V9�.����Zpoy>[���O���R�Ǿ��U����P��B�D�*5Z�=���#�mΆ[��a"��e�͂f;���/�����b'�$H� Aj!%��HQ6MJ�$R��c�g"&b�m^�>�3�'q����MK2EI\$��&�;�\\�w���>�*硶�:uN��X7���g��ʪʭ�2�2�U�Fwh�BO���֐ǲ�[�R� ���#>&5��e�\�%R�W�������aL��Ǆ��k�w� P~ϙf�����^�)[�׍Rua1�SN�gJ8C6�m��׫x8(�����<"�m#�ԯ��(��P��h@��3SL�&XEe7c�=*�xCȺ����=ٖg�>�"�7
�
��.��HO^�?ƀQ�)͚�F�L�Ơ�3@��e�9O�hD���
�x��aAk��Ʈ�3�����u[D�3T0
�(x���mr&6e�%j�1����̮$0C�����R�f�`J��lR"Y'�q��"�𻜸�`gD>&l��A�u��F�|��Cn1�*%魉s'�s/��TB2�����n���;,�����&@e� ��S�s�6��*΅��(i�Q��5��]�\���mCX��0W-�L���#Cޖ�[E�Ko��ǖݳ#L3%"*&���4�q�������'rL�y,��)_y�ȅ ��/�8�I�r�l��d%��T��%���~�1�)&��8��,���:�~�hbM�-���y���8΃j�|�6_e�����g�
gՠ�Pڪsq@d��(-ǿDΪN<\�3_�������j �Y$�j!��j�CK�@	�;� Xk`�Y{�x	�{P�!������(� �܄��|���?���n|����u�+�q4��2
�%d����BD k{�c�,�3��a<��瞏��C�Hg+֙鞈\ly��,��p���fkZ|�ݬ_��rAFX�|��  �0�X���� X
XM��ƙ�}�y�%>C)Q���W;�::9��t��ك�ܭ�}�Ӷ�;3��H&��Bayd=#���=+���3�<i�068{��&�H/��.�c�*�Xj�;���[�b"� K�vz$�*��a��7V���q!��w*)X��`�g9fDy��?��:�J^�����R��L�ż+?�|
}����̫����#l�*NZ�  B��i����EtIH$ @� �w�1l���:U�	��[|b���J���� ����fAe�p &_{f���⦷Lg�Z5��f�vٿA_
���=0  ޘ�袋���{��(h�q��CrE�:�av�i�Q|����ӐgЁD�%¿����W>""��$�p�=�s�;������L���eG:�֖:��t(�0��ָ~�4}ۏ����;O���mx��Z�Q(в�r.c8���ق��s�9i��� Q�vF:��Z���YBJِ$��-�8��טz���R� .>��]~����s7[Ƙ�d�G�
4����$Uzzc�e��7�'9�3��݉i��uȺ��ֽ�K:��z�¼�sb�I�`Od�钁D\!��6 j�\�.��V-�;��H#j%L�ˠg���d&�82	���e������Lk�f{'���7��J�4�=�g�!ʉ;�N/��P��aJYj��4��z�Ǥ�%�Nz�O����-�MM������賶b��
ls�⧵�LsDp���u�F�����c\@��b�D;)t��:��,�]��1�c��v*p�|B�2��̂Q>#	o1^D�Z�x폿���	|�?���>����V-vN���x�pD�6L ��'V9�w����-��f�������q$$\H��koJ�ZcI�����	}��!1��4��d�2& l�^�WS���~�]y������98�=n�/�-����P����{KQ߄��	'^�5"��ܗ���ڝ2E����;��$I��Y�I�u8����o�U�� ��`;��]m����K�tG�� n�0��Xk�i�X����]�!q��rl���R�n[2"$����ϗ���!�T��� �H��͗B���F0$���D�ҟMN��iĳׂ��Gw ���h�&4	��"4Ґ�K�7i�����W;\�� ���Q�u@8G�M�IQ�4CYd��Lk� �,n���x��~W�/\��bv�r��jp)N���f�)a;50֏)mH�#��$Pv/#�����zD��r~�1,y}, V�c�]�!_ӹ0�����ύ)
���Y�rJ��]��5�v<F�o%�낃��vk��l߽3Nz����Q>���1Z��@��yX7����i�^ܤȆ80�SIdG�"��WXə��]�wAKᎪKX�R%�8�IOh�	l�kJ;b� i���J.�N18(���Rm��������X@����mcZ�_y
�!@�4�0kZXk� �V��)��s\v��VXG��FH���R��&�gT5�&�of�ǈ���*�!�n��ո�jt!�80��Yk�2���� Z7 � ]���%f���Awr�Z��W�����	fD"�Jc�K�  ��+r�8F毤�d�ȳp��������Zk�V��N2P�C`��ȟ_j�Ov�1E-�g��	F�1`k���y�?7'b�r�����*�w闃�J�%X����ǿ����}�; ��ѮF��'3�M�<&,w���*�z��%O\3���J)�n��8s�� $d} �n�5m����~�����Qx��y��s�襣�%L��\����]�h�.؋�A0`�� b H�9����DGƚ�.�����p�
3ǭS�v=MU
��X��m\:T�4[�~��B+��a���Pn,xH�"�W�H&��,�䏩%�"�&�	��Ht;%;�<�G��������'>�:�Y�[�ԍb|�����P �`k�Ф4N!���2�4�kf����#1`Rq=6�k�Z�=f�f3�c�@0������cŬD��i�Ƨ����+�D��vg�w2Y���5P���\�Y�H��h�U
x
�X���yU�4q9���� S�e��PY�+�,b�їZEx�.{h��� �p�:�R=�m��[�����i|���{h�3caO��)�E����}t��K|�_.�\yT�����~J�)9���
�<K���1��M֋�^F���>#:�� �QO�T�9�*���%�����3K�Zƕ�7�����p��:*�^�'� �F���^k ?��uE ��N��h������+�3�tH�쉣��o�(k�\�y�;�V�`*Ic��7Q�L���B�8��ٲ�=iytrg�\-`ǚ�� �c�f8YZ�z���Y]E��(JTD��|)P�@
+�wI����Q6YZ�u���1�v��i=[��Q���4u77%�Jj��B`�^���4r����T6������ȡ�8��Փ�Gj��r4��B���&Kq!1�#"[΁���w�^2���.L���L�a�ëy*F�Oe����^�� �RB�<�u������H X��z�����i�,v��k��5v�wpp|��
������7��}�}����p���X1�p^]:���&��H�^���x�i/=�g�V΢�ﱢ([ԶhJ3^y]��BZ����~	�1{ ێ�֏�CBμ�$�3���]���3F�����π�����C"`�h+�^�2:!T�WY�Q��!T0o�7Pß4BX�٤�_��2����*�JXktF>��unO	��RSd���s���y�`�|l�u ��xf��Zhkp�<�j�����������1�d���oh�F3��)�I�=�|&�-�7+Xl3��Z5Ȭ;��H&��TJ�DY��q�}	�-�b�Nx��i�{��!��`C��)'lb��N#�$���葍�(-�Ԏ���a�q�|��|����HF/$�*'����1HF�\�X'��<z�SX j O�؍cn7�9ٙ=���t�Ƣ񺅱_�{~�Cx����q�}�>\��p��y�۹W
sF?�ܒ�Ax.0{yVڅ��hX/��^p!�xb�h(E���%�;	c�|�˒n3͚ݬq�~�C�6�%瘸�d�/,Z_�Ð�f��n���[��7��[\~�<v{AH���Z|���S
27I���f���B7��:{�r��_/�.Y��DuM��֔�@8�hwn;%�f(K
8�d��*նI��dQ�����+)�4��>��q��q4; Z4f�Y�¼�G�V.E�1��4���s���(&�R4&��1�|�=��i���>�PB�<��\��0����E�N��S"� ��t�u�b+8�-�V���Dhܞ��:��P<^G �|� Ō>�5p<F�s (��L���gyv7h���G��e�}�b˾�Ăm��U^�m�#���T_�6嵞z�5�sr�f;;�����GX���x���{\:s����5�j	�KP6��9H���t��X3gǽM�� �r�CQ
�)�)�۠�b�N1y�P���I��W�bd{���|a�Jo�rL0��vU�c�����x�ӟÂ4�7���y�;,pNWB"��W���f�wD�����*�����|���#WZ1�C@v�� RD�?$ĂHM:xå��
�J��)&��y?�r�j�St#�N��B9��pKa�f��$8�c"������~�M����<n�A|��O�§��
��E�V��Ŗ\)
����XE6���MQ������d�8�t�3	���*.,hxo��Z��`F�2�0QZ�9)��j4;ӄ���$}�%CZ&� Hކ�A� ���!Jizۣ�:����Ȑ��Q���6��B@�� As	������r<��i��KM*�'�SJ��[a1��ix�p������w����A?[�U�5���Y|��>z�
���'�^���bi4ñH��(�x/
~C�E !�y548/�2�Z��W
�\�E�g�j����t������s��$,C��(]?����`NNp�'�F�l���%��8h�$#]�'q_�;:N�w��{}�5Wz�v�%��Xes_2Y!gT�	�G�
�Z�А;f�@Y�(�nxGP5���ӀU��F{͙�����3��Ba���a�PPD0�s�[o��~/�܋G��8�-.|����Z`A��2�8f�A?�ⶥW�V��䭤���R�:��-���m"�r	��B~@
�I	R���A�$��{���~�
����7���z	�E�6ћ(�&a��c��v�5.�AjL��l̥�qȲ ���%�|��A�t��t�bL����U�&b���DwZK���D�$�p<���O�����@�D�����"�>�����\��Ghp}w����x�/�w�w܅���1��,>���
�o}�wv����v�)�I�OG��V��OB��=u��d��d�
�<�@8��9��� %�kZ���H��o"�e� 1W�������^ux��z�`m�,�`ae�5*FFt�A�0\�¹��	�+�����a�*�B�aL\�e<r9��(;LH�����/����>��ir �k5Mp 0`/���w�	�9�#��,B�{��gB��[���Y�����g�
:}�W=�N�_�����|�[88<�9é�l.�I�X�W�f[AI���sg�/�Զu�O�R��z?$q�G4a��e�&s?>�-cD.��<����u����Ξqm��A�1�d���1�c;X�am�7�Q��S3�h���K��d�)>��1�\�;/M�Zo����6rYgY��!Ө�:�Sj�)/z͗��OY佱~�f{�N�к��2n�yǻ��_��X�y?�� _�'~�_��W�-�D�x�-��fiM������5ň����BC.o9Y/���L�A�_|����`��ݗu��u�6	��l�gL��_����0�� �-A��k�0h݃�K���@��{C���c��N8�!��ד��q6��g1��J��ȈS%��X	�xKxB�r��*����)F4�@�R����aZc��>J�ٝร9���÷����k��h^�V���_q�5:��
]%�,�ZُT�$��f�R()�k�hoYwI�ܜ]ws5��Y(���Pj1:�9��T�PI�+�?<x���5-֪��t��iA��D^"����1891�;���a>W�ʢgw�-��OT����%A7��9�l�5�~r���r�zmѭ���6-�&L8��<K�@i��ź�Я�";̀1Bӎ�X\���XO�R��	��r+ར����K�иk�$<��q2(��@x���3���`;�s����#��vpp����ϡ98��y���_G��C0'G���7�����>�[��3���t3CC@�\�m[�w��.<�3i�h#<��f���Ι���ZE)����P���"�?���A�*��WZCA�c'P�RVak��טC4;@���0V��$����p  �I��r�ʨm��e�`n>֯q�R(r�<��U�F�+��3�-�n��)��D�S�cv����;5��LZ�0�H�����ZT����u1yջߒq�ր�[�`�1{�W^�ē<�au�Z�{���F��_f��˺�
���+�s���|��3�Z��]�G"r�	�B��Yx�ť����p��g�Ʃ{����>�3����/���e,���ͱC��h����~{z����"�᲼o�z��59�3�A�r    IDAT��1�)�=g��M���+ra���hƼ������-@�Xh��0Ъ�1��sJA������B�;	���T��a5��b,�BC ���*�LYX�����Ų't��&Ƣi�if��ܸ*"�ͥ�w:>�q�O��_� ְh�s����e�('�Rʻ���C	=!�f���,�N�S����>�Q#�{[&Ɓ�Q�T�l���D��R[�@ŹHܗ�Y�Ve)�p�_1��&�� �>��fѢ��Y�m4���!�g^����{>�O��{7n\~�����߿��w����5�����;>`�O�h��։^{M�;��4�7R�J����R�����#-|ɐ ;�q�<S��)�O>&��wK��ɲT{w
&.�fc��M2b�-�����ƙ��IP�)�ZM�-�[M�k��m���u�,-[�g����럻.#7�t��-���b�Lg�s���6���,�Nc_+���Oc�X�m��bvϽ���Ga�~/��|�s8��j`O:43X���I��'��H<�aw2�4��������^q΢I������	�L����������`BaiUE�~��p��iJ�)L��$�TJ����У��R8��ġ�p��ic`awL{CT���CA����yv�X��$F�I��+�rA�D\ٽ�@��}��I�%�&"�q��Xf ,z��4ԭ6�_� 6xq5ǹ�~o�����5X�\��×���������Yc�������hܶI�4�m�K���Y�j�+఑xŊ,�8I)�x L����G�hg��~*���@ (�s�x�9���T�P�u�ТPcc�Ʈm*9|�S�w�Q���l��9��G����h����=7�Y$�%�/c(�����R�륵��!�.r�D<����L�t@y6�VGdjD��#�����-�V���_��u�^�s�
�����O����r	�羃s{�P�����Y�6ñ_�# �K��sT
5᭦��1����՝���������$�y;+F�?��c�џ*�3"_��J� aD�v[9̪P�K�C��p��M�5<�`(�K�G)��*�%�)�e�Ц#2����R:�H؃K�Oj�)�郉TeM� 5ѐ�vB�P� �{\bw�����e��9$<�׮]��h�&oM���8x�q��C��so|#��w�
��;���?�Iܵ�Bwxi`YCi��l;+�ƻ�{��銵f��/0`*r\�+=����`v[3
�����x�ʱ�ʸ� 2	TF�Gj�o�dS��fJ��dN���X�����Q���%\ghE������Ȣ_}?Fߪh��LoL��ܱ�46!�B�$��X��`A�g�6����y����N;��"}�"�$i�&���y�$�,�,֝�-������O};�n���xv����8�2��G��K/|��Bi�~עYi�b����<�6�}PjJ~Q�)&?%t����|��H2ڭ`���.����^�q[������������5O^ q�!Y�򆔨R%�ޔ��0)��3h]��A�_)X���,%( 0zx)+j���l}V,By�+� �u�kT,�WR6zY�a.}Q��FD��D�M�~u����kK��d\����?�ν���q�:�\z��Ͽ��?����݅�4�NV�����e�P��hvv����z��r�D���V��bZz�'�/��gf��y��FU�E�٠�P������B����o`�9�����͖�e�e�I�l��+�*0�R�uU4!c,BZ�ic�]g`Þ�+(�-,*e�}�'jRx�Xr�؇E���i�˲�0�s�ܛJ��r���J��p,j���z��1Uﻪ6�?�ON@��	����z	�W�S�[`�.��,�=������{'f��)/�������sx����k �w�"�˃�bh���_��9-��5��á� {����|��T�g̹i���S�S3C"�&A����N:2[�t�Je}+�,M�ؒ��`HD:�հ��`]ٔY�1jx�;8z�c4R�pgb]��%�o��1��B�x)�&�6%�q�b
ן�D��o��7�(lӠ7X���h��<���~���c����KxU����'�?�(^5��t��Ŋ���g�������b���=1�<:v> �B���47��>��R��n������3�	<Ԗ�0��$��iC�R�4�9�|�I���c~S��R��j�g�p\\�P&|��l�2g�6j�i���7����b�:'#�ް��7ۗ(���Rc����%���IܖIm���m�q^zE{E��t��\�WR�BNPY����n�6|�5Xl�Jws9�k��@s���j`��߮`���o��o�H�����,ϜƝ��ih|���=�\��}&��Fn����E*g�7�'�\��!�/�֞���X���u3h�~��pwE�����%���-5
��9�"�E!ͥ�P������h���b$�"��� Q�/<�u88���˒vB V �P�����coMBF�7��\��hP~�1�m�`��0G^x&�Q��ȳ�yc���>8�H�G
�
��;��ټ�U68>���=��'ރN7��V��y�?�9�1 ��l� �����N;�V��v=V�lo�����G���~1�<V�dr콮A��"r��Գ4^+�O�!���:�r<���'8�nPB�xI�%��CP
���MR�Ĺ�sc��=�Qkϖst�� c ��3��F�JQd�cu%�W�*xR���%jIB��p��&��}�W/���J4Ɗ�%�{��Pߔ�}��>6��~���u�L����0����ʢ��~
 0kf`,�vk�VP�q۩Sx��3��G�f�:�~�ؿ�ո��?�K�_ą��3�{��\F0�0�����X��f��z,'̜)zSs\>+����i�3���NZ�d��r�Z�3$����,�yJ�TC����A7'���5^�L��B�.K\��H���ا@r ��$��^���	��P>ۏR*�pO�k\ �q�{ֆ�<�{��Z�3�Z�fd'��e�yX���b8�ѰFc�9i4M�þG�,~���Sg�/;��/�/��n�t=���]��
����8Y^�{�D��u��'�8��+/c�\���<ľ��35�"w^M'G�T��Q�ZGz)�q�+��L�c@A�Xv8!�����d��<ue(��06B	sx��'cL('FC�,��DH!<�r��Gd۶EӸ��}�c�^W	DI,�%?y@
U���~��.Ǆ"I�)SLh|�%A�~ׄ�a��}"�~�8%
2 [���'����0�n��f0W��e@��K�q�=gp����[��۸��pt����A���~{?�V��Y+s�>�籲�zHu��	Yʵ_{�ޮ�����0��:<-d�����U�$��Z�I���7[��U-z�@0Њ@��ѹ(�AH9������z�v�5
3�艁�w�b���	�(7`��EP�q��#.1q6p�(R�4�K��2ٱ���0 j|Z@�Mΐb-�r�!턐<66�;W��(�DP��T�)�}w��R/�/\�k�:�u�?�C�\��|�ֶ��W�z���z�����%�������1��q�?ƭ˗�������?��vk��
'�{��a��24Z� ��;��/0M����}GCp�I��X�fǫc�~�]8u�-8���8z����r�[_H�1	���]x��u&��i���P�W�ϰ��SK"���Lk�t繙��f'�+r֤0�2Ƹ�FB�2Z�>���@���0�J��p��OBR��pqM���S0mz'M�y�Ѣg�я�l�u�RCa����p�^��(�?�괞"#��;����&\��R(�a{' �ib��`�A9K��.�`��ƍ������&,�*Ͳb�ȿ	wA-Oy� ��Ě��źcX�0[h\��a���^��g����[�'o�Q,�]x��������˟����x�鱠=�=&����9����勩؏�΄�]!f��1jH�hB�n��L#�ٶm�,�7�X*�a������Pz�N�����&��`��)�5�x�}]:09G�����&ǃvǢ����W<e���)(��0N�s�F58���4l=P�ײn�aG��Yvg�ܞ��։|~Cդ��$�R
ݲs�aO�3�wD��!^/��%0_P��H����29g�,Y1id��R� 7I�cŽg<�.΅#'f��]�V�+w��Z�e��~�c��őjq�sx��:n{���5���!�������gt�V�p�w`k���`:ٿ���3s?��"�)��#�ҔDD��`���q�X���˃l�ְx�Jj3�����Y(-JCmO�ίf(�&�N��(�T'�d��XZ�OJnN�.�W	��&���ɍ�c���r��V���Ҹo��59��o���Oy�|.ocϕ�8�q����qa��4G~S��$@|���w0�,�}��9FO������������K_�]��9�z�<��_�g�?�+�~�v
��f�zt���0�͡צ�k�-�|8D~�K2�R��xa�5<��by�CP�Bʹ�$�M��	���x9z��$�!mp8o�J�X�P���czF�������0��VT]�a,T�܌]��@1�鞓hy`�w=�� ��݋ȑ���m��U	C�^m��ݫ~ԇ�E�h��W1��B!r��EH��
��Azg{x�C��[��a����=�g��c�ݸ�n�<YC��lt֒�_�����,!�E;� �PP�a�N�c���%/^�Z��{JZ0�8�f�`�t&��|���iЩ�|��8|R{5��v��Bw%-M�5ӭ�.�<ӫ=?%H���=?�fN����d�Sm�ڝj
�1Xkc_FE,I����`��x�HN�a�C[N��`@:R��H�7�鿄G���1E�Xw"F|3��J������?�����cy�x�d��7ԙ9ԩ��^j���S�Z�U
l��Y��Zc�U�Z8��L�_�8�+��J�����2�[ۂ֍�?,=�Xs�@���̇����38K��� �RhT��1z�06(Ƙ�R�ȁj4mn(F�r�$;'�VN ��tyhmp�o;��q�ҧ����m�
{uT�X��\>s.aa wsrѓ.P���ø�����Žm����������5��� ��X�������)N��n�x&������F"D�劙������{���<��0t� ��1����v9F��B��d&/�Űn�^��C��f����vI�б>W�ls�>C����E�"��N#��Dzw��^��������M��6eL��b�Su���n������}�mLBc+c.�0ȶXy�(��V��2����L��U=x�c��p��y���'��=8���x�]�]Y�pt��羅28�cu�}Z`�U֫r-�i���b^�9�)��|����)H�����vN�d�����Z:�ϴn�֟�A�Պ ۃY�@Ù�ÑXe�����"�z�"��?/��C5���&������g
��A�ɛl����v� �9��~���'���#8�c�����b�7		,�f/��������Ie8�G*@7X�����x��������)���ʧ�_��A-/c�j-�3��Y��V�]�ݝ�.ߧ%�7�X>FaR;k��Zh��6M�5�6A�����c�G����D�����4eP%�ȧp�ד�����!b?���|��B��0�L6Nl�B��6[��>����P24	�+)c�x!ڶlSϘP!}&d}c�T�ٗ�J��@J�p���u�h�1�����7��k'�B�.ɵ�p��:n|�S88s����oĽ?�_���?Y�.}u u��*P���m[�Ot??����)9��Ƴ�6g��z�wh�f�w�&����@����Ι��.��-93Ѯ�B��ab].6X�(�tn�1`,��
�bؾx���� ��렔F�= �/�4��~bi/�]}�v�Y�7.�r(k�:�=L���e7h�C�> �� ��1h��0������gJ�٤I���)c�~��=0���<�����>�۰�z�/�7|���K���v��VƢ��N�>9�\5�=�Lð�+Z�V躵[�V�����K��Mg�GY�APM�3	��ys�P��ZCNTKb掱x"�i ���k�l��m��̇�NwMJߵ�H+�w�a_�^�c	��כ��x��)�Ķ֨1�5V��Z��d�m���T��m_J�l�k���)��M8�f�Md.i��������k��?_獙��ڢ�9LG�ewZ�O�'��N����ƙ��}�|/��t	Gy{����3��j�p��:��1��ʴi|(�1_'RY�4okk��L���'���7p��鏁gs�T�%�s���Ki/��vސ���ѝ%�,î-l�;�E�6� ��_�}�	%��ݓ�Cg�G���0�&9RJ)k �D4pE�K
$��j��f����0�#g��5�ZM0�R��`��t����3w���[���y�k�o��_�`}��|��
��m3��;h����Q���ĺS��n�FO���'���`0���w4)X0���ǀ�,t?m��E>W/�`&���]w��~B𪐩xâ�'4ґ��
'���R�'�1��yY�ڽ�wƴ����R#f5x���P8�_3�V�CP**cǄõ��m�W�qDq|9=7�NwƽiAj���Q+�Ϸ�e�^/�׌;j	�����?ǋ��8p�2���x���ނ�4�jm�f�(�1�+q'��W��e=ec��r|���uCZ������ɩ�cs��&�]�ORX�'��Ƕ�����M�Sk�i��naTM��K	�'}) ���}��+�c`��x��Z��� ai�����d���#9$D��#7E:b�M��_�`�d�Q��j������n���?MNP
���1|0V0��'އ��gq�'/����it��A�-q�va�\J�f@��O�y��ط��Z��V�(��8��vǤ9�@�'x[p���%�1lљ�r��ehk��K�3���%0۴���k�K�Hph2V. i�'0���;��{&h���1�C�)/��(��~�шPL��o%�R��f�l�)��cB��~e�v�y�/��Zd�z_��xv�к6ha�°�c0���zA!�����b�a	����V�0��s�v\���O���S������{�O��y�<��1�&�`��+A�ϧ�07V��\�M�M�k�>ӻ:�N4 ��k	�s�dfg!QJ��іTb=�a0�L綛����7b�`,��Bh�E)�9�T��Jh���ʠ�"OH k; .`��{� �B�V�C�c���a���9�� >��qi�-A5 ��{Z{X��Cg-fq���KAZ�|��4�	lg���:��l�MGN�"�9q	LEN�����	n�FG�|q�})fX(�a�n�Bs�����vo�S�
��1��/�C\�};��ɟ�.��_�l�,��r޻``�.8�3�Ƭ�9�- �zfz�./r�� БM�g��<�.�X���z��V���U�+#`��Ojd��%�ÃY,]c��C����۸U�`N!��TF� 7��g�H�}�"2"�b?�]gT�w�$��"�zc�h��Z�Њ�9�8�R8�Ҍh�Y?F�n��S��te�$���J9��T��-=kE@�\	�Mփp�d�q\B�2pL*�$;�7�u��͎$s�x��^3'�\
�%��N�*Fi���}��>fR�i�'�}l�$�!�fF`�hH�;���Y����x�;��s����~�-?��8x�<���'=�����N�1S,M�v��w'�����Z E$ L�%^jV���*��V����q20f"�U+(n<�8+'�;��9Y�Ƣ�=t���X�Z�`v�����A��K3 �0,zW\��    IDAT�[g�܁�E�4 �`���sS��1�F�ڭE �x�� G�ƍ���@�0��^&�&�;L��5S�dJ��Eo�����gR��'���${���D�+��5l�B^����D��Fw�����/�0��7�m?�a�}�Ҍ�o|O���qr�
v�8<>���i�v����E��Mh���p�m���J�%���c@0�1ͥ�ixٯ����~S[���T�@Ș9~o�&�����¬���k�R<�ƫ�������+i�VjmM㭵q3+x��a%���7�Fv��_��U��R۾����쥋x�K�é38u۫�<�8.��Q<��Wq�0L+���ڂ{�mT��jև)�k��ֹ�������r��>"r���7�z��%=�4�o����R�PW�G"���d � ɿ�3�B��1�8u�DN��˅���>X�n�h����ג��2��{S��]I4�c��ޝ*d,����k���<a�����w�ܣ��hn@��w��8��_�@��Z�mv�T�����v+x�"����g��M�\����i2�ݱ���)S��kLp	�k��{a��8�5TAۦ��`/��1!�^\P�3v��j�Sp�脬w�V�J��6��X��_ɐ�-����9������S���������o'�c��y?����7a���5��9aI=fMef˕)�������]q^+ckrl���%��~k_x������loHR�]�n�n{�{����e7$L �@+e��Hhl��w��P����`���a�\��M�ĸܵ�Hn�
�l���u�ޟjs��`������0=���g (@׿��8�؛q��P�	���?��O|g�1;3�=c�Z�~U�k�}y-,$Y�T?�D����؄�rj�$�e$:Y�������Z}c�Li�D�����5�M�a�8�nU��& �1�4�!t�8��~����*�����٘00U&d������M��#<e��uo����k8�֢�{t'�8� ���*��{����?:8�ț����G8~��8bB�f=ÚJ��,�7��d�c���S�M�$���yR��p�b,���es����n�ɂ
��?�˺Sq2�a@�M%��m�PG�d���,{9���ar��_]�R��
���}�݄Y�&\�Fc}t�3gn��f���~��ʯb���0�5��<���ٟ�������\Ǭ�Ew��B�4�S����MN��[7e�nv~���T~/�>O�Z���p8^��0n��U$�w���)�SJ��}r�aFo��|6�R
��˘;��Ş Z?J����-���������V#��z�h����H�6J<L;s��
H���)��-��+)S����n��q�� /�s8�v��s'��]�걷�峸x�#�w��3j�k�E�N���{��4xL��<fJ�+�E+�9q2�@�*�%� D���P���~�-.�\9���#s������U�� �HSJ��?�8V5α�3�����#d�8dx�tq� <[3�OI��6�O)e�i�e���{�p��Ǖ�5辇���k8���qj��\�����.��|�b���e۝͡�P��+,��m`���cxO���C�v3��;y�l�����njet,�9�|Q��,�	y�����ف��x�E���Tm�`����\N=Dl�$��������#�S�v��m��6���/uA��br����<�}6��C�A$f���;4��m����x�#��S����v~#��]��X43����V5Y��p�8|�Χ�[��z����2=v{��k�\��Xه��I��"�[� �"�,��ƺG�U��$�vb��2�Rɖ�^�	$�B�[¾��ކ���'vy{�iЬ���.^����so�QtKB��g��?�m���'qj���5:��?���E�Ֆ��$%�<:���'�>��=���lZ�c̽��67kc5ֶ����p�)S�uS����cQ����G�u>@Q�C
�?c`R@l��i<�u[��l.Stff_�O���1�6�N=���|-m�\�mK9�7��������
���|�����~��c�O��������bt~�����<�$T��m���:P{N��ل) �����!�G�M4h��Y8���^_�����N�1)1|�}1Ơ�{�}��V���rK�@�&����R~�֧�w�N���Y{n6����Wq�����'ޅKk���ů~_����`�VK���h�q��Utm3�wS�S�o�P�I���V�*?rQ��3��v�m�ڭ�P�m�٩v�a2S8/��2~��j�k׮��:h�Ѷ-�]�EkW�/����=�~ҽ�f>V��W����8��v��Yc��E&@gPSs�Fg�ʘ�[hww˗�a�q�Ya�4p��y|��?��O}{8����;p��߆�[��+��GX=>>�f|��1E�6=;,'Џ��ks��Kc�:6�6�)�k�R�#�+k��պ_�W��Z&�'��&�h>�G0ȝ��L>z0.�<t�;d��֎)nazv��@5`6ѝ�u����[o�S��Հ�a�
Vu�d����cc{���1h0��3�� �O0�l�oM)S[9 �51�\�.�<�5 �֪��,̦�8��P��c]~�圁F���Ņ`��[p������;ѨX=�i|�w���2��]��5��0S
Kk�&�V7�w��L�]��s��j�'Z���V.N5��H� ����K�=���GC���.�����f��(�4Lۣ_ �0�K�@�@V�j8�����(U�pj��$'�{ƢA�6�U)?o�s��x�\��)w^>|�Y2�&���c$�]l�F��D��0W5k��b��a��g�̜�
�C�ó>��)���KN��u��M� +ԧ��#҈)�`(¦Om첌g���m��;avGR.Ui�T%Nj�Od����y�.sa�X���vк��i��X�`�M �IP�G��z3��&<��M%
 ��� n�5J�5L������������\{ǟ���և��z���pߛ߁���˭�����Vi@
��ԍB�<�W )zM��:�a�5|�q���*���ӎ�Y������aݬ;���8���^1"���^�|�?a� �{��[��{0�Ӟ�4���۸P�g�d��x�Y� hjAp4+ui��[ZD5�#?+�#=�Ky}�Zzx&j,�MKMS�׶eL+=5�G>}o�3ہaƊ�Sg����ᶷ<�G��X���O}�S8|�%���=4�Ma#Vj�H�p�p��0w@��DlQ���"�=F�Xh�A�`5k`n�����vv�X�ccp�8HBd��a�� ǢF�Â��6'��Ɣ�>G9�Ssdb5VJm%;�3����Q�E��j}�pL�m��LYQJ�7��|��8��P�v-��8R+�4���,f��ƬW�zc]^h�D��8?�Z+cV+fF߯��g�M3�L5Pk�}cq��gq��t�����x�ïÎjв��?�s	��=6����r��ޛZ��fF
c,��()
��<
4�h�&��ё��.�WI��z�0��r	�;װ�tҋ@!J5�:Ǒ�kt���{�̑g[������O���2E��fJ��`MVCA��y���pr�4�A8��/��_}��4��E�
L��|�HG�'���K�4�ߑ��sgJ�k��Et�,�WX�3v���.�]�N���Z�naw�a��Y�S^>_��S�tl����q���v�p>�����϶��pB}c�&�pVޯ�1�[t�|(��c{�c���
��qcKW�ʆs܄����sWð�%f�ŬcPg�֦��u�sf��9������-���;Sc�hp��QX�V պ��n�3�<�]<��o��?�����ӛq��Ǳb���{��O���P�G̰�tKY'mu�ܖ0��H�[s&/�Y
��o�ɣ�p�a��e��7D�֤ڜ�p2� �~Mx)}���bR��D��=C�c�х0�p�a1՞���&D�b):5�iS�"`��n���*죍��ZG�w���hp���s���a���quy�ٍ����!���8�hp��.�_ɈʾJg��3#(��y7�3M[��3X�?c�+�����i �`���V��y�A�ػм��xf��j}���N\ٗпm	]9���Y�m%w	������N�-�$e�5M������?F$��-ǱF���M�}F�nml}'M�u؇s1`��eY�k�U�V8k��0;Ѱk ��i� 2t�=�on��q�z�����^��X��I)�3zN�����B��X?�e\����g.`�{;��8辇pa钳80F���ΰou�;Տڼ+۬�1:�[Ei=�I���G��JZ�m�ڟ��G'I9!;"��F��q����c� �*"r�,#y'k���I*�Ob��i��Y���&�����Ci\[�����G~w��p|t��Z������W��Y�r9�O���Ҕ]�p�of�����9-�c�}��2@�C�p��ZX�̱X,p��8�����'���?�?�����B���]�ʌ1�қ}lQ�{�I�ilk�����:CYW��P16���"vSQ��`���g��>��\��,���؄�A �cP_�8�mm����	T���R0�Z��R�,��p�M�1GTG��m���<Å�^��\?} �*�L`7�<W+���T�`�3j`WՂ��+t0��[��,��͗0�g_�f��������Ƶ�Y9I)��@Wc��}�:6���mل�M��X�JY⬸.�Zd�5>[�}Y#7s�H�%���R�c���Ҁ�A�M�|m>=�IK*���f���6Მ�qJ*�� �K��=+\�-f=��}��hϜ���'�Y<���>��Fk�?K�vd}v�|*$S*̗%�&��1��v���Pɹ���г9X���\�z��������]<����a���q��bi-�߀1]��FdƎN�Y`j��o��|�V���&�������T�4�1x��%l����Z��m��1�l��1X��G&_2�C:��C��:�I���g�����]��"�����߀�1֍[O*9q&��9�m��<U�Vx3rCm� ���>E��sl�e߃Icݯ��^��/���z
�f���	<���n�V��z[k�'n�pȡ��!��ܷYOSnYwM`u`(�	�@�h��G�^	�ر����!qVc���z���mN{[��9-^H��<s+Q0�i9t������@2���0��9��L�4�m��8'F.�ݘ&R{ǲ�j�v�9�w{�]x�{�N��(��c��.����}�i̵��34���K�6�S�3p��Y	���M�[�I" ��}cv�`�O3s4�1�Due� K�L1X[k�(FC�'G�݊�o|3^�����x�2������q����nâ#p7N�$�o��IB0F��b$[P��|��l�6�ߢ��h$�荽+�0Ō���&i�n��l3ܯ	��Q֙����P�>q���ȶ%��;X}�^Hw�P ��>��4蒗|���N߆��^���{�?��g��w?�Q�U�kV;U/Z���ao�D:*�i)���1��� ��Ō ��gemqf��������bv������5���`k������ֺ4�j���6	�@�ZZ@7ͽr]QF��30�и�M��D�cD�đه�^ �2�B��bd}�kZQY,��\R���cZO�;g�����o(���_:\%8�zL�ۆXL�m����&$��n�=���,;ƩW��}�O��Q�n<�����7��S�awwL��B�~t,���F8v��@�7�"ʜ����}�0�
�������}th0��~<���ٽ����_ǅ?�]\���p����s��Uu�����,%�j{˵:�:�f9o��i��Z��h䲔��n��D����c8�%a�_Ã�]������1���ڙ������7���~yTUw�c޼�0��   $!�H�HJ��%W\*�{m���7��������ՊK!J")J�D< ���p���xW��􇬪Ϊ��~ �Q�^ב�?3�W���v|}#mч�s��秐9v�����O��я4Ǧ�|@��[ec��=W����%��sB+�<��9�Z�HPSK&S\9��?�K��&�_e40[[㞏<��'�0��&�k��eq�cs۳����ۣ
�pH;7A��p]�8�f��0gDV��غ�9���3g�����<��R�`Zi�R�cp^b��#/s����Ei�� �C)I�i"8�pk�F@�suk-�BR%A���> ?�C9�q��Rz���GP&	�V��n|T�@*IQ�8�1��b���ul�ր����w��u�*��p6dL*���;�in������ck3��k����?�n8��c��O��"�\DS
���0x�ϳ�a�@�>�N΂F✿j�DԪ��;��bl�/�h6cS��H-��H�� !YS�q�l��r._#��������$7�a/�k�.q�/������ ��ز�Θ������L�2���i��h�%�R|��J��<V�s>�����
��\�}~�J�i9��62q��{��%D|~���E��jU�g���0�w��Y��Tkl^`�Gb�R�����Ӿ H>�@� M8N4kY ���CӺ��4"����6`�b�{dݽ7����{~��o�
�P������7�:~-��ߊ<����3�ua��o����cb(�b�l`fSdR"��c�u]=�I������x.�M�]�|�.�VH,����*G�;fɀck�$;��Js���nmc����ˌ/���lB6ؤ��DLQ�@��:9��cq���^kU��eW{������R#���f�J��%%Z�Ֆ~9g�ƒi/�O˒InP(FiB�
�rH�VV�VT3"0NR:0�׺�D�I�Π���Pʏ]*��%�T���U�7� \� ���y�\N���d��qeYѣ���8��w76p[�h��6 ����\i�
�{&3�lG�ֻE]�8�e�K�;�ɲEu�~&d�&I79?3\���q�}w{���}���W�\�iY`�֔� w9*]ܨ]�Uf1�Ug���)�m�������c��2P妤0%NX�����G��ƅ����:��}�3d�mQLv8q�"?��/��?=Fb,i��Sgdݚ��������J�]�����<t�j���l�Eªۋ1%}�1���ol!1��eg�ݠ9������)��1SPG���8�/�5sUe>�B>5��#�����R�"���_��Ў�~]���Ӌ�b2�rb}�������"W�~s��}���g���ڥ1[����!����ּ������g�b���a�.�]�� ��E	ŌK�>�/�fw�N��'�c7ތf[2=�0)3+�:�$��}TDw�q-��CX����{�֚$IPJ5���ºb��hZ+��ss-�q���n���:�P(Ŋ�Xt�N��ڇ܌%�>�w��Q��
1'�aD�X�"��"�p�ɡC�]�z�����p4����^s�{�e���l�����'cp��z�Q�K|Cas葆¶�j�kR��NJ�����#§.�:0�Q�p�D�����)eiq�d7�ŝ��,�]g�1c=?��_~�7��wȷ�"s�<�)]�u%�έ��5��n�g�`�%�ٻ��#2}��p鮿UH���eL�2frU9��bLl����w�+�D���8y���ǐ��p�e��m��Q���5��!�q����:�%�J'u�&Qi�	��e�MgH��'�!���_�s_=�.7��Yn��Os�=��ۻ�@e�lc��dC)�K�����Xqε��%PLl^�0��������5��~��$��nč7��Jr3f�R`�Y�ro���2��L(���~�k��I}6c0]�\eDm�Vi%j��ۧ��K��^v�L׏~7fI�trn,LNщ%�f��J�9�&�M�l�/.$������A��,�ޏ��>�!&���>�#��.kJ���Y��
WA��i�E7(Q    IDAT��E��`��|�=*������~u1e�s�����`E����,˰F1>����G���%/-�f����^��_��{�k�C0���a�S����2/ˤ�.�֝ﾲ
�tϦcA8~��ZW����Ga�����X�1N}Pw�K�����������F>TiyƤ��=���x�޵��a���j3b_K�"~�SK�1�tg�F'&�����x����ܷ���ŗ0b��]��O�噳LP(aH�%���j�I�V��n���o/�a��|��\��k�e!w1Pl�=�S���?�r����?�Q��f&��
�e�Ÿ�����!>֣0�}c��#�Z���k��-��p���B�}���[�v��/�kA���}xSv9�����<�����fU��.�kc0�:Þǆ�"���Ήza�p@��ǒ��&-�2�r�w�b��s8��7�ؼ�n�hD~�m^��7�{�)!94���`���>
�Vʤ�j=���X�K����QK¸S����EʾX�~���m����KO<�+�eŘL��`�u�4[Õ�	ISo=���hL-�kW�Jٱ���'��[~5"�_g�p��v�ӹ���c����K)I�"�
J�d���}L�s0h׏��u�^Ex�r�C����6�1e�#�51��^d�c	��4�%�O(�q�H��l�7���\��/�~�����{胜��O��~�RhL>EP@���
��#��]W���Z|w]���a��ST�b��g~�䙟1�q�����#�G~l����S0Pf������>b_�0�]�_|tW*�ה��p]�i�����{o�v�~7�/Cc������Yi�!!*_��;��c�� �@� @�/��\��w��L�������މ>s���<��G��N2�6�����mg9ؽ���ۼ�أ��z-�BH�NQ�R���ح\ڶs��u��M����~б=0k�HWZ�r~�n� ��\�Y��!����
{�iJ9���ɿ��$o�#$g��ԉO�Q�u�&�t1�d�:\��w�QF�9�2�]����
I�x���G��z����� O��{u���_sl$�y��j�Z�v���\؅6�	|��	J|�,�E��l���9,g9I�aeB�
6ӌ��e^��_��_��F:q�#��=��#��mv���Pޠ�v��$86h�;�n��g����©]�&�i�%���䰴Gq�M~��_a�ҫ�ƻ�4[�>�4S��a��V̎n�	_}�%T��������1u�5Ax�K���Q�Z���Q�Ƙ޹�eY����gw:�t��?B"���(-�@8k��Yth���%�QYB�nPM�PΪ� Һׇ���י��K��6A�q�]��&�ݷ:t���#��]��[et�:�����?%��+�rLj�1Z�%u��eFA�4���6�y�.����u>�����:,�Ɓ�8)p:ũu6�{?���g)��Q���5��w�U0�g
I�h}��̦h	�������^�Rz�e�˸u�q-)����E/��o���(�������>��Wwآ���O�]�lKꥹLr��.#ў��b�Pi�����H5�~tC�.�m~�"�{�9X��S6�C���SJ�ԂV������]^���	Nmmq��əG>�΅�\|�뼲{����{�87~#9o��������������[�B<c)Q��m�UܺD�}�����F���P��g��{���'ٽ|�a6�L^HȂFu��]s1A�~&"gw]A;�_cc�߷���"{A�v���6.hI�`��]�K���G���Q��}o����P�G>QB�d�ĢŽ����9����Y���C>1o��?��EW�����Ω�(Na��X���\����|y�)�:��t�2?��י�}��c#�d�+f�c�C�4(mA;HT�������1�]˂��|Y��7wH��)�R�шL3ҍM������a4�$������|�Y6��� ����p`�TXRm�䇨�n�h�T�%���'6w}@�X�`R�e~�ݲLJ�G��.R�Cr�~��%O��<�����T
�(���&c��u��UG�������k"��.��B�};�[?c��f(6WE	��l$�P��d��1����~��/�淿�*��i����q�ݿ�=��۫�d��"݈��0�}cj���A`l�"Q�T�tʰL�n�aY���Ɨy��믱�;n��~n~���q�t��tns��#ײ�׽_��]o���=Pӕ�خ�o��B4)���ڥ��=�P�����Nw�V�u�g��x���q��4A8��^R���4~�~d @)�u%EYVzuϵk>��3��WgC�:��,q��6��h�b(�_��|p��|�3�D
�D)��c����wmR3�9����5u��#�#�G�C�K��Sw΁sHY�9�:����kK�p5E���^'��H�Ag��N���M����7J�V���.~�k�H�L�K	��-6JS�r	���[�)��4c�����yP���[j?o���b_z.S �rƦZC̼�'I3�88~#�������~���3�}����?p�;�`�)JkF�8�p��K	R�S(�|�p��>�n6��4?�
�B����/g���輚��7���;"���UˊG����沂�oO)��U�n�ж�;�.B��R��a�"�n����a b�k�y����f��:-��>�U0�FU3M��k�\��B�:��ffi���R(����E?3Ε(�TuՌ���՞w�,����}��� �}�����!���-�
���˜�$V֠t
B�� ?���s�sz�8�c���3���7�z�+W_�MP2�5]�.,F�
���h�]�_)�ǈL�^'��z~O��HQY�;�0!��D��y~	7p�=�o��G�{�g؝���\ A��	R�"J�����c%o��z��>V@�@V��1#9�</�J�h����]%*�D�ERX���$��T:TR9�3��)� ��AiE����PR⬣^��b�K�qe�tl8��s�}����3�yf���Dcj�.�b�J�GQw*�]��,��ew�J�7���x²Lrx�w��	����ƚ7X����";u=�=�QFǶXw��W^����I^RLf�~��ҧ����zgq��j�>�׊W�e��R+�xק>������������K˫�~��L3&����������m�o�}�j-�m�Xݱu~����UgU�L��b�����$��{}Y�����7�y�UK[���Gc�\O��>c��e��X���-S�H4NIr,S[2�%3g�E�	M�ŕ[�TQ��̷�N��y��r���y��|�������d(�!K(J�$����N^��okB��iA�{�q����"�'n:˻��Ӕ�$Zz"���Qt���qSC��O�����}�5�Ƥ����-O��.��R�᷍�T�X�iX�HW�ѕHb�
U��D�����G0��Qu�Y6���%6a���b�h��kC����"�`=r�K6o7��?��h2��Op��/0b�D��o/�����j\�P��Xh�4�(�P��?z�t9��g���'��qQ'l���ͯr��_c���p���,�J;���ֵmHm%(|�'D��i��-a��k�hua[C�B����SX/CN�>�%v4�G���>&��/�{}�M}�o��/�v��V�����G;�K���ѵ��,�5���h�Ȁ��O�Y�3-s
g!�dk#��!.Q���<}�S0Њ4MX��g~�Ͼ�e�d�])8v�{���O2=vWfcReq��"I2�$k�v���(%��b��P�g��\�\��12}�u^|��ߺ@>�b�އpۧ��R�|�8-qJ�|����D ����F+�m�{���4Q��~u.�>w������� ��XHS�׉�F]`?�c+^_[�K���߬����e�/��_6����l�s�:��_BiZ�c,w܍=uƕ��q���eK0!5���h���Iv��|0��<Ӈ���(�`���hj�W'�N�ɯ}쳤�[)�/��׾Fv�
gNlS3�Y�v
��o�P�J��o����s�N��.���=T�w�X{G)˘�p\1D^}�a�=J��b����ۿ������}�s^-�	J@T��b����� ;�h�hߐ��N���^�e�iJ�e���s��IN]w-��۬��W�Xj�a�=RR�֞�f�"'�d͍����O���8�7>���f_I������I��YtN`�+��b����i���~<���ZQ��
�ٔu7e��S����۬�v/�~�#�WR�VB��
��,KR�E�[V�k�Z���(3��]a �^�:H�c������Uk��C�E�矶l��/�P���.��Z�I��5xc�:����JZ�z��ZW-�ظ�ԭ+K4ɚFZ:d�xkz���[8~�]�)�����e���8�%��Ô�([h�W-��rf�.VЊJ����`,ؽ�6��o�G�ﺓd6ac�<�����ҵ�3%��� �X��iB"����q��(g��s�#j}L`~-D�b��8���n��e�iU�.V�C/2b�����w��[����{��������h,k����6/1���p�xw���._e��զ��P�RR���"�A6Ɨy�O���K��lIy�iN}�a�[�`�2L�4# Ԣd��{1��2c��(!�RڍNX1gu	�:�(������*��1�Wv�k[������'���a,(��0�%��UWw�s��%BO�ӎ��)��5�-���b��c떣����Њ��݌+[�cb�#t]@uTx��|Ѳ�:j,#'y4$�W�qC�>���(g�gS��1[�M��\�2���'����0� Ǘy�'?`��0eN�$;����,��5��kW��Veՙ�U\����+/3�a6d��i�~�X���9�@M���7��ۏ���Ô\Y�EI�S�Y�y)�_����ţ�>�rTF%V_���>�a�G9C�c4����w���O��؞<j���UD~Y�Gm�'��m���H�a�g�T!� ���/���K���%���}�/JK1�p��Gy8%q�v��к*���$IH�`�ed��W~��_�ϘW��̧l�s77}�w1�o�ⴄT�LI6�a�ø.�m��I�k,R��<ᓴ8�p�@� �JZd�����W~�*w�SgX��יe	c[P����U�������.����=˄��
5Ρ6��nn�)��Q��C�o��9@���,b�*�e�,ƹw%����hw���� 	����"���4`��Q9dߠn����ۘ����+?�����LSN�'HC�XqX���q3����뫳�7P��n
W������?�N�b��O~ȋ�e��)��!�B1t�I1�p����f���w���/Mw��+��6v�}W��z��-[[u�bAy�{}.}�������Ǹ�b����UOHJ�4��vl�e�o�l���%��GMJ�.+B�J�؛�2J��YB,&+1�0>�!m�.%�9d��O}�+��;�7^cm�7~�c���OR�>î�1�3��בh���>�C�ƺeq���q��V!D`�V�P� F1+r��e��P����1Ǯ����]�u'�j�Q�+�t%FXd�)\�r�W1�}�:�a���m;F'c4q^G�b���K�k���S�8\3���0�!b�(�9J���󩥫vv���.����"q� �e�#V�""X�1�6�3������v�F�d����ʏ~��X�l6#/K2����'��[�-�ɯ��{�������i>��g}m��"��s?�[_�÷vH�d�Oj,n� �9�ZJ�rR=�H*\��q���g ����1H}�����pGa ���{o�CRݾ��lN��_�,�;�>��E��!jW�91�_�5m5A���Ǿ�,���1����,yYbq�/˒b:[o����4��l�&C��;��Nx�k_�ҏ~�����u�������h���cT�Nְ��"�o]֍ߣd�dV�(3^~������02ct��=I�hH5z�bl�<%�i��*��c�s�kq�ދgm]�\��o�7�=�j=�%4oK�̝A�;���J�LR�&"��?y�����
�X�u��Yb��o>AUhSW"�Z�dK�\+�m�9��:^q�a]��3��8�����φ�$8]�kZ@�M����^��/��xNUJ�
��J��L2�6�c������S���O��}#E��O����8J85"#�%S5��s�
>�L�0T��'B���~��ih۪���X�y�P+���)�vks����g�?un��Ǚ����e���r��_Ƽ�c��5f6�(Hȇ#
%PӒ�K02�
�D���R����
�>a~�znJ�(�ø&�_;���"/)��hmp!�i}ݢJ-�81"Α�»�:��R �5�����ZE���:�zra4��-q�� ���ۅM;��i��ZW]���k"�<sE��(hjKv�֖#�\�3e�V$
%����ÖB� �y�ẟB�&D4֡�D	�
�����Jb̐��:/w�"~RP&����1��xm�8%)
�R�}�0(�I� ���]^�����(�j�;u3����8y�)r��,�Zc��P�b�43R�pI��!�T�/Q{7�qt��I����u9Uw�Jp%W��(P*����)��~B~��t�N�x��?�>v������шLM��{(��Wmx�PX'�&�*^i+e��8�ο�D���$�~=9c��c����
��M�^X���T4)MS�N++{D1�3+�Za� ��q����-�:�1��)��g�
\uD�u��CRc�&+;B�H��@H�LpȆ�V�g5���}�~�/�23D^!Ҍ-��T���wҏ.A�qY�ι�𪑊���]?ƻx�ts����+<��G���`]I^�X����I`W#��ˬ�'|֧f���9q-�o|�-0yHT�!]AjK
�y��������k� �� ��w���͡"W;+aݍSw��ϲ�lnc��t���2�7և���>Lt�^��>_6�>ɬ�yw�����߆0���Q�U�m�!<C��kbg{5zWZg;*��ﺟ�~��t]�)��s��[Z�����~�}?Z�[T'+j<��⋜{��%;s�k�� Ɉ��l��QN�h���4R%U�UIc��я��<-+��=�h�p�����Oq��և�l�|�n��%��a�K�67PI�Gl�X�5�%��v/��S�]�c��{�F� ��-Bo��6�+���m�Ѵ_yw4}��{ˁ k4�r��|�Ӊ8�X� b��P:�\��GD��2?ː�nX��"���ބ�̻��cg�}�5W0{�u�=�J��
�A&zAz\F��������Z|�!�b�p��z|��@��)f����l�� ��1��,���?����W��r��t��)��|�B�F��6va>�TV�~ƬV�"4�������2F��}k���]�b��n���e�\V_wE�ASg�l��ph���>:��;��:�$u� �/!��3o[�*M\2W'���x��p�X�?����K�دj���h=���[�,�\A��K�7�G�p�[��a���A����,E㼶C$��bj�g��iY=�~��N\3T�2��j�JXO���o?�c�I�x�N�u?l�c�2В�8
�N���ZSq���e��9�x����j�����j��y��>氻�����.dtk[�����m�AF1⣪P�M��uK��"d�A�	~TFo좵n]ˁ��k��q�!c!D�}Ͽ�/��
s809�)'�}���n��9b�m^��o3�g��ګ�T���qG�.�˯���u�`���o��NgH�o���o�>�{od_�Y7{�������c+�&��q�B�F�Ssʦ�H��O�}H�(sK��q.z���K%����v<�W-�Jҭ��Wߺ=ʺ�ǵ��c��YGU����+k�(#aE;��dRk�����_g|��.Bj���p|}�Bx�Bߌ���&,����O���
�Q�:��\Qr����){    IDAT{��O��[����>:�Y!����:E�e$I7r^�h�o^[0ZFLd��/$�Ɓ-J��#$��b�p���~���[��s�Ïp���0��$d���n����>�+��G?�D�1�1v�~}�����儂o��B05��	W�N^� �׳]���o� nގl}��ѬS��d�ٺD�s-U��ۇD��¿���71IK�pF�U!�����҆�?����x�@(�3puoLv�����=��\y�����b]*DQ2�'͂�t�����^lA7�;`����X����`���}�r���p��m]������3O��5�OI���k9�s����q�p޺a�[�>b�m�<Bi)y*V�s�{	�Wؗ:�DW���X��@|/Ş����c��-L�����J���#��R���\6q�=R��vT�FU_�1�������8���cs���W�z=8�Ota�Gb�L�����:���T$l�}?���g\c'у!Z{��ٴ�̋H��ġO�m�E��f�b/X'��$6/9�
���'���w��u��w���x'c ��`����*5o�u��1t�����'�@%�$IP�F%�ٷ���Q������I����?�:j�Ҋ�y~��j��>[�0�]��b�[5ϟC-�F�Ჾ��s��׫-�z!��)��a��Ai�㡇��� �f��r��3��dJV	]<�po����18���ژ(v�����z�Z&>Fw>f4Xcw�0�o����<k�O�ؔ�[Wy��
��O��X{@�Ǡ�ޥ�x	���>�H_8پ4�}p��c��K��c.5�ڭ�u�<�1��I	ZK���*.�/c� (@׿b�����}��^���(���&J�Gׅ�;'�Z��������Z��ma��\���얭���+�x��^�3�����;)G]�B�f�Ϊ�S7m�s���x�k_%y���\��������%#qY�N�,HӔ�t�� ��FG-�p签G�s"Ek� 'Ha9x�%~��oQ��2�����\j�R]�	Ga�$J�=�W���H�.���.�އg�m�*���&��Llm��G0�~r��R������̮�6\�xc��(�}����0�A���g�iY�:c�V�A�e�lU	��1�Q�7*�c��M�(�b��k�0+8���y���F�J��!u�B!�C9|jZ׿��~�NB&��[0��]_--Ed�&r�K%VY�KJ5"{�]��8˄)�._ᵯ��|�K.%�K֫��;� ֐�粛j�w>z�[��\9K�{�t�񻘼���[�>�ƨM��!��932D�~,Cl�;1�9l�
��E;�|�fW*	$���@eY׿Jҩ�XK�����5%|�t�:��j���[����үVB�%��m���p�e��7�������9ԴĦ[l��>��7�oJ�+�	���yG��;��*F�s���}$e!��8rla1dL�cc�W����*6n��cﺟ"I�N�NN���d���^��-���w���t�d6��yN���>�7�7�i���e}|�����:c�g.�����p�Ǌl����Nc�s�&�Z_�1G��vaNBB�7uQ�"�@Y޷�5���� ���Di=�r~B�C:\�&�ǚT��쳌/������`V���}��Dy��nT���;݃ZR{E��p������#-õaל9��{��0M����O~��e;��S�-4ÙF�3�,Y��A�Q��q���QhL��[s�\�6����i�b��49y1m�sm[V�����/�s�ϰ�i���\�c���FU_�~oJn5�`�	�3�n��QJ�(�2�/+��mǐ}�r��(�.E��q>��u'P�x�;�BN�l��[o���j��Y�����1��t��g���>�5���_e�-�t�!�����Ll�e��^x�\:�Y2$��6O�����:]ۅ�cvC�PK���fa1A��`O����n�����.�ע�_����Hp�!Rz��_h���5��Y���,�x�� M\i�JW�y�&�������:� Q>#]"e�����ʨG��
'S�P$�D��I}�7�Rz�d��YI�[�SHBX�H4����8Z�j�[5L�!C �%0+n�#��Pb���O}�;��/~�X�2����K!���Y-�HKQ�؊�QJ5y�-ՙ�h����s��?�w�X��0��#%%��h���`M%I�� �d&n`@����in��r�G~��xFy�e����}�*��l�1��k�����IL"��2,%�̘�uGǹ���]�s67���['F@`��|�+���-�\��ȇ@���ZI2��Ɓ,)UN�*I�`�g)ؗn�2:�)5ߚB�P $��
�"����� �[>���&v1�c�zU��P_�J�����v���T���_����~�xfT���{�2Od��Ü��=)�A�� D�'8t���U�m�Ъ�܄ ����#5�e�Z�x Zq8���i���UF�5��D�H�P��7��ؼ�F���9OJ��cY��>;{o#F뜾��R��ϾHve%'h�c�U&8Q6���FV�H �~�i+<.T͜{,�6.ʲl�H=߿ �M+��D
� �($8�/\Aek��vN�r���+\y�E6�����pS�3�
�ʗ�v���\�N��x�s>r�Td�(�ȴO)���MBxC��	
k1���
g+&����j]y�Y`-��.a6��@���
��TX'�U��AYz��Tg�i��G_�l^��2XJJ��w��_��_�$�H�3�he,�U�<���Y/��߾�m#�Ru�k�����8ι&p¯Z��A�>HS�0�HuJ���?�������I�򐗞x���|?J�~(��6}�`�cR�a*������R� ��!zu�`0�=)�=�:\g��;)8���s��{��t�K�z�7�~=�1���p�C�Vm֒��l^ �d����������y���.m���d0����9�5��О�^}�@:�� �sf��(AST���&w�Ʊ9)�bʚ�O�(����x�H<�#����r�j�׾�O�+F�0\V�~(�����[g���o��gm�ߤ�//����/{��%/wq��l�q��Sg)�c�ю.9��1	,��kWb�>����|+=�*T�lZ0�)�x�������N^˽���\>v�K�h�I$�,!����]+���R�Y�;Kg���d3�����k6��/?�-Ƥ�6ظ�y�q�`�fqW�欶1��c�����I)��Ř3#Z��� §.�zo(#_��Z���x�M$��G������sM<��B1Dۇ|k�S�Ď���%�ֻ]׆n���[�U/��e����"(ϵi�m�3K�+ԝ��q�m�l����=�{�
*QP�diU�k��h/:���0A�AQ�
�ߨ�eG [-:��7ƠF[�\{߃��7s�N��>�Sfo\d�X�1%2�H�18�Ш4C8�(}�3kK��f�a��㜼�Z\�B��
�Ӂ����9�I�1X�ΒI&}4?�-�2gZ��Q#��Ր�g���`@�#�$�T�n!"�!�&0N����B8�fm�H�-f9B(�
���y�3�����:��%[��yD;7�T�[^�݈
S����m���!
�1� \������U8�rq���x�5�ay's�m'��:�l	02��0����������(�7ݍ��v`@�[�8G�q#�ݨ���[��G�v�m�:j��&�/��!��e����°u�v���>�0Ô�D؊xҩU%W����u!��^�ٳZ{�5ֵ����1¾j-Ş�̖��Fbm]�>hXH(:���I�]$�E��M��(�Ќu��pP�>!Z��H�V��*�Tir�+q�:~�s�N^ì8 ��:���&��Dc�k�8`1�Á.n��nY (�6��:�� �t����O��ri�y7�a�N����=�c��)Z����,�� ���ɤa�2�8���a�����/����Ғe��j
c�N���!k��J�	��	�1�)2��h��՜�c=�9s;o���1�0t]G��6~��p������7�}AlO�1���_|w~�v͙q���܂([[,������a�I!�<`Om����^����Q#�YK7I�	֕��C����e�*Dj[��Ʋv�inb��.��_
A1˱�J(
C&Ǚ�������`}�4w���q͍8[ɀ$��Q:j��/���}.��v1LP�*���ť���'��Oؾ�Nnx�['+����hvA��"��K���B��6���F��վXO�.؏z�c�F��R���d��;�6���XuY����:�p�F6�L������lG���}/6�>��(%6Q~�k�E�p���F���r涻�"av�^��oa/��@	��ҕ/�����N��tԈͷ�m�U��6A@̳ӅC:XO�xKIn�ݏq��0�˨�_���s�b1P�LL����)���k�JC*Zz{����,�u�ƕ��?��x�'�����S�M$i�V���s�t��^=-)*D`�E��5��1�D�5.�y�]�������[?�G��n@��4�-��~/���"��8�6tL*oI.ϕ��v�/��[���5�/:?C�L{;�ƜHt�*���^��oR�)�fG���u=�o���1�ʰ6,[MkX���ɣ�X��
2���:�<�0�6�^|�G��O0�<���}����:�(�8!	��hL+|��#��]6G��P:o,<�a._������d��'��� �F���&�R�&��QK���[w�C��o��E���~��a�?a=^>���3|V�����Mb���$��u�{$���S��O:��3=�Ѷ��~�0�w�}��~� ׊���*�dB){�fo� ��^~�7��8�����Jʬ�s-f�=NɾA(nޏ:f���\� F�"���z��J�k@|ԥ�SCv�Y�[n�(^}���럒��I
���'y(�a�T#L���py��
7Lɇ�r���ڒ�Z�`0`��&��$IН���$ܷțw\�HVkJ�	"�0��Ӓ��g�����?ñnc��Q#Դ�,��1 F}g��{1B�l��U�X�Qd�Lb�RH)�^���v�W;�z#t�����l��B=�8�Dx�>�����n�C�������M��Ǹ<J��� h-�p^F�cc�>�.�cߖ�!KR�p�2�DHP�P��,����o3�<��� ���2�qŴ�4EÉ��k��&r����0�t!��8#k��@�u��p�=���M&�M_��k�'�65�_U�i͖�C���B��s�����L�,�V�,����E�%z+�j�p�IىZ�<w�2��}&�0�q,PI�[rC��Pme����k�3�i#����)q�w����0�a��9}��$kC�@#��L�k)�\^��p�6�9�	�6��\�h� ��I:P9����[�	�! R�q�����?���&�����_断m�e�]b�(�t$��R
�4�L#�CY�2%�Ʉ��Qf�r��6�(L�)J��C�xJf���:#��UsT_�xk�B�VdIʬ4\r%�k����!�>�!��M��&��/��ޢ�'d�-ݺ�Zf߽[�}�@���W�~,�>�ʼϕ:�U���l����j^���a̍���v�Q�Z�eG�j�k�O��i�3�8v�Z��y7[�<�����������D��(�j���*��V���y ��49J�<J)��
�F�Ή���w��q�����G���OP&���Y�F�\�1uε�U���#��X�zd�(.H�V0q�M-ї��G_�o��*ɱ-N�ykk��l�a8	8J��>�4ܣ1�4���l�Le�^��ص�.Zm,�}}0�[Kι�V#�>�M����plmKʣ�{�aX�N�~�}yۥ�۟#��H�9/i��Q���e��ׁ�����N�9��~�ַ׹Z�q�ܫ��0�%��C�u��5��ķrD�)j"_]�}7G��E��}`ij�8�tM��\��?���1�~q����]ʽ=�����)�$G^U�aV�(qX-qΒXHg=-IJ��7�͸R�ɕc}}��a)�T�([cj��=����P�cR����i�c�ָ�������<r����e�?�(/��"�t��O�sy���&��n���M�}XVտl_t�z�{b�t�R����{n4�F�a��Dk ;}�D���VB�:{�66ή��������շa�"��u��<�Yn��@$ل?��,�V�Y\�a�+����R"��ڐ�tڤB.&6���U
�.q���^�H9�n���?���k��Kǣ��cЉN���օ�gmsU�?��
��1�4�����Ϣm�ю�kOq�����mE���"������a�{
b@����L}LqۀU�'V�o�������3�Ԕ�^��pT��Jzeτ5�����,@Z�V�4Ѥ���g]��(�\J�R!�$Q�4�h%�?��o,�@�3�Ki���y�T�|�Rp,^Vw>�L�FS�P��9��Q�z�����rM��I	�Ddar�L��2e���8��g��?�G^����QLC�18<��*�k�Xg�*Glip�A=��� W��~&���|G�>�~�5��mU��J2kPVb� �!��m�������k�7\�� #�<�7��%R�����C+��^x)ӯ?g�$NH���4��$R�TIo�"�J����ۂ_o����7��Q�7���GV�L�#����C��8�&��0����rm���>������#��1J�9�9$K�W��y����]a�x�u
��jMV7�����}��.��+p�JW%*�^E�'ՑH�&s�}S�����a\M���N:��|�^�Q����y�<����F�O�h�%3��rU?]�����bh{��.a�LB��8�}���N�]Cy�5�N���s��7ٻp��DpX�KHtJa�v$y%�����C
8����sp���l��6G+M�c�8D*1Xd"�U����>~ɉ�Ҕ�ŷ8����d8.�hfJ��$q��t�G_ð�7k��	�%�5 ��V2{�Ϻ��O�h�m[!��	�l9�3g��Lr�q�␗�{	5�c8����La�,Qr�u�C49<��Т}�$��rRT�����|筭p�B��k�1`��:oI�*�����<�sBa̰Ls����$J�)H���@��ǱBb�$ϽP�脡6�dW�H@`EmF&��W8~��8���H�
Y/�:V|}&�À�]j��BW��'2\<�����ͤ�uYK�ͺ�P�P߯�5t��
�kC��Ln+���ӘB0��k��s�2�J�F8�(�3�m�G$�`5"��޽�u�*�RM!(�p8�ɔ��c6o����{/Ce�;��Ȋ)kـ�����F�����{>Mr��~�:�̛6c� X,�0 ̔� 1I�W�,�ږ,W��*���U�k\e_�%�JWW�E�9�$$&���X �����8�3�=���ꚙ���sΓ���,!��|V����xX�17ZC�f$h�]����y���h�E�&\���ÿ���.qh0)����;^��8}����p��ni�z}ĥ���~=�Ei�g�T;?�h�$j�EMw����x���}�5��$^r4�y�������E��$3ǽ>�����G�ť"cs���o�p$3�ҘV��ks��؆�A�o��yۥAo~g�Q�p��s��������0����qD�6B�`�n��p�4�ծw�������.�@>�qy�61��|��Ͻ�3�c��
��C�W���i|�`؅_�㬌P˻�-��*w�`+ ��-��.]kՕ^o]t����rDV����e=)�p���\����uD]?��s�] -5�T���cz;��u�a7���K}�7b�t�z�q�����G��͇�g��L��������f()^��T��Nz�$�N+�2N}��~U?��6�!��RQh0>CyO.b���{sx�Ȍ��o��w�� Q��sh�NU�ڭKa��}Ȳ�Y���5n)��rG�L    IDAT��k����#��|��gd������?���;�2�&�i��:B�}}V�.��ƻ��]Wi ��Yiqt��Y�I��?�+]����y�ꈹ"���U�}d6]��43֜�Dq�g�㕿����*f�}��ğ���ػS0�:ĝ���ڢ�v�xm��&�]��#:����C�EG��N�Eu���+/p��+�������|�;�3��-R�9�<�(|w��.F�=��s5��o�w�c����`���1�LIU���76�z���(�џ�E/�������}8���S��ӷS���	�3}���=�}�+��q���N7�l�-:7�.�����B,�*��z��Uȴ�і/�@u"���ۮ��Ϯ��H�(�B*�)�?�1�>�$~���";��b-��N0��P"��w16]�w��.�T�t��S1e=��̊"�v��Z2����3�|�in{�� ��?�\��fc
�R1��z7i_�]D�!�ղ��.�4�Bc�M�cɭ�;8�=�������Y�pw�������92���$��D�M�n��_���&��񮜣Vݫ����A*�$�:�܅<���5~K������Zo�}jê����}N��X�o<�u�����)�N�$�������䥿���Pn��ξ�������ܙ��#v��x$��O��څԻ�߭�^Z��ʰF�'���͗x�;�b��3�����F9�Nn�K�Pޕ��.�	Ⴙ�����ص��qU�8�*J'���FJrDC:���2������~}��"�0Sdxo�:B��\'}�l{=-i_D���T��t���i������Z[QӘ���ƷMc�EY��{ėO��'a.I��^;Z�tmξ���=�N�M*K��~��j[�w�c�ҵ ��/�����J�'O1A �/}�kܼ�*��$�8�QJ��w\uF�}�#�sdQ��BN�Y\�ǥ^ �f�kN=�>�>�0�.]��+����A b|��q�+���Aγ����V��W|i�������S���5����������8���Q�1)S��-.~��g{�tƥl�d}�a:`:���f8���J;n�o�K��*n~U�]����\Roe<Ww���Z�ܥv�н\,���%����\�����u9W�!�G�>1��`�M��ï��W����X���o��<��y�X�9K���n�uW���`�oU��{�<FF��L�у�X:��6��l�J%��ĳ���3��zH��.+PN��P�+�#��}ޯ��QD���t��?�>�/��։S����9A�4q����9�&����{]�s���y��:�՞�/1�=BO=�TH� JxWa�����B��β��j�A,��T���~���X;�[;�K[J�k�7�8��R��Ou����A�q�/�{1��)��!��	�X���9��"�x�VP�t�s��>�E��/�*�Q��}�ԯ�E�x8������k��C�%kv�K�����G�N�|��8�lc�x�����WI4���N	/���Ň��3���?�Y>�V����y���=��U6"M�,F+�P��DG8�\']�B��mb~U��k�=�.X����	swۖ�}��~LE�_��A`�jn�B�+m���l�h�K*i��.�A�:Y��3��[2)H�60�pl�=.|��y�k_d�w��>�q���?`W���#ȝ������c7\Vk�c�?�|�BƹŸ�Y1cc���K\y��$Y�>� ��z�u���|.���=��^�Ҵ��o�}k��=�Q�#�*$j��\���~���;2ƭ���i�B�V]'�]����W=�&�� �}�R_�s�;��1�=��F3kC�*撆Fl�@s�R}�vS�/���GX�L��)�C/��mB0�.��A[�m��P�{P���$��"�B��+�t�G>�I��{�5$�wP�֣�[���=EQ� ;R�$bmx�2R��zoI�Th(	Q�:NV��l;ǉ'�&9~��t���mn��Qx�(l�p���s�A�*�>g>:�AW��U���!�s�+3������C�Û�;o!��9����H��9�Z�3�M�r4���,�� ui�*<sՇv���w囯�S_��3�>����/����]k� �G]�/�M5%��~5K঒x���O��q[Қ>��k���y�r�h=���Qٔ��S�H㔣^r�K�;o}�ˬog䳘���y���g�s&�M�n%������X�1Z�}�u�4��T�o
M�ϐ�`0�ܼ���<Gv�mf<p���QD1F�Jcr�^���Uvk���������������0�4ki�o3~�u�w��9��#�t�ۻ{�\)��J�� �}��E�&!=R��	��b.���&�u�שg)'KW�����N�8��k�Bi�b��b]��M���T�V�r�w�`[a�\G����:�9�(��4����v��^�2<@1���ܒ;���~7�CG�	o����n��C��8CԎ?�6��/�>[�6C�W��h-��~!,��!5S��C��ȻZ�w�WL/_B[�d:EG ��H��&�6�*�G�ۈ�B�sX� ��|7�~���~ ifܾ�?���q�����h�I"���pk�@�llbo6	�W��ޏ�3��j���>]k�`����B��>տ���;A|�޾�����_ ���u�3�X���t�؞�>��*�2��qx=bS�]��dNa3��>��/����}�u�tp�3��)�o��]�p�d���_Ő�����Ƴ��F+�$j@�w����#���x�u�\�ч���O"FC��H�@X��s���,v�0�1�<h�[�v�1�1�8
뉕$q9��ב�)�C'x艧9|�	�(���k-Y�u҅.����>�l���4�v>�4�z�>�}��ų`Wk���u�5�q�+���c���J��yxU)q���Jy�0H�ё�ySJ�TP�|���-��3]�JR*��Ò�WX#:,�<sx'����,�2�$�,U�:�s�Hk<
�R�K"C���y��(�����l;8���X+֑�m�YC���ۼ�Wϱ~�#3.
T�6C��B#�4���f�$g�<Ғ*���vx�'[�d�$��#0�W��U��@ZO�I�d=̹Q���G�M
n�^�?�0�p{l9��%���� '�0�p�������=M"��7?�lD�s�� �9�
�cl��i�U�
6�:v6fmk�̆,c���qyg��>�;�|ϯq��;w��ů��s����Ø� ����8�8rL݄b��@i��6�Q��aL��c��'2�s�V	9�j�*Cj�p5�NR�B8s���S���1 lM�����sU�^���Aj@*v~y�
�x'�����(�0GB�P��SՑ��]%f�n��1!���ㆺ:��.��L�aWZ
�$$Zᐠҥ�yջ�3le�݉�;����W�y��`M�����c�I�}��gx�3���\���1���
��Ѕ$E��EЖf�� )u�uZ�_�o��'x�/Q�/�$Կ����g]l2%�!ټ3��?�#���2���#d[���txaq�a2�L����\T]M�*
%D0.��-8�T�R��%�0�j_, �@�;r�y�ȥX�ȱQ�_�ʕ/��G���p��1�CED�+��UX��Ϗ �G���`�Jz��Ę���Ԩ(F�/Tm��(�Z�h��Z_��ˆ�Z�*/=s�L�W����4����\P��Wx!dLn����һ��4
'6/prQd�P&a}�ڮ	��FV����s�M�gئOu:/�!R����3��Θ�'�I����g����i�Ǳ�T��>!�e���� �(fn��ko��.r���RY��U����-`S�M���ns��M�R���a6���o�6��F�+�߼I"Q��ޡu@X!����څ�R8u���ީ`���� EG�D����q$�hĥ��H��)����z����b����&��_������:f6��XX���Pe�k�U�	��[�o�C�"E�+�|�SɆ?�+����%��k�9��i�{�qN[ဦ��AJ�
��?!q< B3�	JHf�c-qc�"�<�d�����qq�����o���{�
f�s���|���^?��	b�Ix��'�&����Վ�؇G�Ҏy��ti��m*�=�sO�t|���o3���Ɯ8}�G>�Q�Gh�Ɉ�硎���l\ީ�zW��9��y�t��a��c)&�\�p�;�E1w�}��:��	^(�wh���_�#�׌n��|w}ֿ���*������}<D��z�]���-�/�S��K���O5�<��9�FDX.:��� W��@�IM�V4b8\��%�L�P���'�g�}�o��ǣm��w�O~�$G��3
?f�y|�	@�sYJ�=V��K�z�U�>+�^'�sX�'��*k�	�[Q,X�Cr3������~������~�;�n�$��$sy����;����{\+���1(�E:GQL�l*͚���
d��M2�E��� {�i���?$~�֏�_��W�.��ȕ�e�D���^��c% <�/Κ��(�(��'J=��3J
8펠8%��o�էz<�Y���ڰ��_��"��gҸoH����F�u��rCB�6�HH�d��-�l� ���9����'��9I����_���:������G�i%��DD�Sx�U�$Ju��}c���jF�o���W�"'
�#���E����L�����=���12#�J�ľ�Xu�r�}��E/�2oAE�˧�[��q�A(]2�Ǡ~�õ_���+o�76y����D
E4�Ȣ�n��u8����e/������.m���ޞ��-����E�j�� h��M��\vqp�I�`]>�]�W���"�ϭV�Xn2��DQL!7�)�lN���̚V�r��>n��e8�g9��Q�{�Y�0Eۜ��u�l_����Q[oOvK����֥ͫ�K���(<c2��l�v�YƣSYp��˼��/�E���z�qvn�eGv���k��{%��8�7HJ��($N
���7�kM,5:"������k�?��
���\���9��`�5���
N�����PSȹE����,��d9�M�-�sC���N���gV�߷�b�7b̋�-��b�b�?Ț�gv��}}��8��ɼǥ��[��|�]���6r��m�"!��M��^�֗�\���N���g~�ܰ+$I�1:N�S��_��^Я�	]Lq�و7b����c4��c.�����u��?�0��xB[kzqS#g��k	�9�s���
s[�w�Ϗ-ǣ8�4�͘���^�9�sO�F��
AX���¯��9���Э]���]_�^�(��ei��\W�{�{�pE/�@�쪤ޱ6�Z�/pM)���R���̥tK5U{y�*o�[���ar���q��8�P��enL��M2�<�����{k�d�����|�W��u�"�D�w'~P����/�`�VQ��Lb�n�38y�G�}c���_�s�A��E�-��aE)ͫEң���i_���o#�P��KA�cf�ಅ�v��&��0��x��\��:ͣ��)l]������׾�-օ�Xc��YE$�Ndۄ����39
�C2L��6���w=�1����Vf�5�c0�v��O��g�������ĥ��*m��n5߶��s����{��&�_hۺ�V���-NinIū�)�2C����y,��%���S{���"S���=6Ә����?����f̉g?ƃ��<���!Ɋ��X�3�����K]��۰h�����/$�L h�Y��W_x�������3ϐmn���XK-:�2�n-ý�wԒ�����H(��
M8�F8"ܹ�����2v�,�E�I��$	kæ�}��Y�uN���"wC�wJ�����㫹�� g��e���%��PXrw�0�v���en����s��;	�� t-�: ��&��x�r�cq�ޓ =�:nn��E�<��>\Xb�o,��p��𱐺#\�Ջ���o[p�3�J�9�z��Et�V��'k�	�42�o�y�iT�Ɉq!X{�'�x�X8��L_;O*Z*��b�@����2[X:�'07����s���<#G��>N|�c��CL�A�-4I��L��;t��~�7)┑5�7^ᕯ~uk�42��IӔ|�#:�=�}�}�?c���(��ܼ�����ǿ������'��'��,6׌����>���an�i���q�}ﵟuU�'�J<x��v}��o�j�GQ &�(���������#\6�>�����W��>��S�!���a�)������������%�\̽����c'�t�.]3��;a�n�ݯ&�˼�U�}3��Ɣ9�Lf9J�"�+��{Ư���`��G���{co�G͊|���������f�r5���r]m,��)�!�	�8�!.�&����(���#gY��n
,��m���.��♮��_K�ڂjV�c�c&��N�l����Q��!Ƴ���g�m�w���i�"nr.�3Y�Sz'����\a�eh%�d�_�������&X�JR����N���măH>��	�L��f��0���"�q��`P{V-�D�s+ll�T;3���(�{?w�~G��LY���x�����a�v�K?~�k?�jf1��
��۠�����'�TW[e�"-1Z�B�s�g?��_�/�8v7^iFC�l��=1�E#���O��o}�)9���~��7�q(I�
��"�0LB\h��+u�Be��@����Ơ��q�G�<�;_`�G9v�~N���͵M�;��ƥ�~KZ��5Z�}D���*�Z=��=�=���`����{�z��}}{�~׸������~����=��?�/��O�;�Ǟ�j�Z��t�U�=uF�����,u�+&��w�K6g׹��/1���Y�$�IO�f؛�xD:�Ө�ƻ��8 mx��D���s�@G���HD8�q쑷�d�ꫨ��#ws��f�y�"wN`}0���n.�a�8zX�
�,�#�п���K��q���A�� "Ɣ�$
�\x��/�C8ͩ�c����$���κ�J���B�ު��z��N�f=��B/�B;�<�T��&K��
�΄g���9�ސ�z$�. �W*�[�g��f� ��L�0�����#n첑�����_{g���w"M����~�w����F#��6�x�cɀYV��B���7���%K�T���e �&�u�Z)�<?�|�r�	��Ƭog����9�0���1W�ֱٌ^ u�����|��p_iKKu�מ���b:�P����(���"ﾛI�023a���U	�μ��?�in+�$ϸ���y�g���H!��I�2�
S�Q���Km�L� /�Hh�����i����7��U��.p��K�ٻNzl}_F� ��d�;��J��p���ˏ����w"ɷ��tOv?��"
�3�y�i�{�)F�?�n�����Ob��,J�y<�:ު#ƶ �'��T�w'���H'.�ɹ/}��7oa2ǻ?�����CƓY1�`9�I��#��� �[���
3E�O��gh	2nWE1c`g\y��o�`;���>��E�\�t�/��0�!�MGxgA��� �-r�K/�!vA).��2��"ٴ`x�	�ÛDQD�#�a�o�}��c����I9��W�ȴf��뤇�(������u���c(��� ��d�o��b�6%�)�yys6����*�QΡuL��x��NA��� �&Qk�(�+��-J$J	
�8\پ)7����+:'�/?����ջ�c" &X��Gy��G���c;���~�����X7E\Ѽ��A���8�8��2����ʸ�t`EI	�t:*	}�"!)��4��%Eȣ-�)A��6'������ed������	�'iH�h,��<�����],���t���C�qU�h��!�cƌD�5~�譗Ho�`8���9W���%޺�x2aC����������cQ��B�Q�V����Y�`�l�{���Z����Г��"�]�̹�"��������ȭÌ�.�>�5.���'��M�>F��
��b9    IDAT��r�u��6`�j��w%��缽�+�J"Q���0��XkI���c~��*)��
)t�;-q0j�n��a;�O����Zr���tO����,�A���{'���P\������W8�}����|���͟q�ԃ����h��`]���&�~θ8|�+�
pʣ���8�]��4�KQ�������f�œ����3Os'�+������h��X�[�X>n��΄��͡V�����n�.��#	��@��j�����y��l&k�^\|�IdY�,�R(p��t�-�W�.�����P^!�~�B�|��د���ף���1~��!c���"͚7l�klE3v�ã���b��lD!��/�^�8��m�W׊���/c����|�9�5JƵ{ʠ[��%�]7�J��˱�A�XٰT�b��Eh�1ֈ�ZUl�2ć�.'�S���'�Igۥ"�R"d�-,I���� �ԇwLh�J3ێ�5O���c�C�-qv���m��
�@��f�slmmA���2�~�K��"�1��5#����(�\�ܥUis{ss;�P����>��M��� D
_���?q�ͷ�.[Uɩ����X�<��y���r�s�&o-��]�x�_�W_|W��1{i�C�(����$�˹���r헿 �S�(i���D$��G��6���/(��em����r������~���f������[���"�Q���;�-�����މ���|��F$y��
��%�G�m�TW�3�XHg�T�.���b�W�,,�e��E�4�?r\�ڒ�Z�ؓ�hM�������ϙ����O?�	>�{�%��] @�ܚ��/���%i��Hf޿�v��  f\+_|�9��׉�'O����G1j��"�ǋ��,ݥ�X�����U���l�B��kʺ���#��[�;;�
Gz�~&i�l�!%�0��![�p�]*_�F��1��c
�-¾V��s���6�[�I�=���<�A ��J.����M��:ݪӟ>��z?��ă�E{渻&�	���xt��=ҹ�ۣ�s4]/�+�\]��K�/�����@���@����o���nOmp�Qa�8��{O�VLR�y�)r��^�cRp��?������Fx��n��낋�3�W�
�*�V�gl�"˅��$c뙊!bc��b� υ�{�C�4��~ѷzư��K�;��3rd�����s���d;L䄽�	�G#���'�:u?.����~�[�}����D2	@�l��Y���5��)�R�x��k2����ܐ[����'PI�ھɥ���s�rH
J��km��o#�.Fz�v�~�Q���^=cJ%I�41eC:�d暱̻�mU�ge��OQ�6"�VLCAp��Q�/	 =L�)�J��Flܾʍo�=��0��8��Gx�g~s�^r�0ٱr��J9������y����Az��@ٜ�;���y�/����m2'8��q衧ٵ[�T�~�_����F����І��э{�+I!�M9��or��W���̧>���w�"�T"̧�H< �
T�W��QL{t��&q�K ���~�"o��e���|��g%����&��R��
�M��4���ź�vx��%[[K�T�m`��%��3��Y�;���������
Q��v��y���A��b�7غ��)j���9�����5.�!;Jn�X����"��`�iiXr����njK������`�Tb�T]��*��B�EhE\RTe0�%�s�˄{�� ��1L$Q��_'.;ͦ5��a���9m��UeռV�HPJ�&��6�au�n�|k>�,3�-�}��d/�ȱa�-�pxl3�6+n�=����rE^̈�;yƝ�C��Oq�c���\�o~�7�����4��N�PJ1HW����*�v�f^����w)%�'�`j2o���,��n��Wo���_Z�{� f˥ힷ������;Ӗ8�m��7���?|���?ev�&������9��O��n2�-i$���"]I�wAs'*�����Z���N�����������|��>�)��C�Ⱦbڃp�Xo}��Kbl�� D��a����a��ŭk!���0��)�8��"쾁��Rh_��*6C�X�u6iH�E쇩����r�e��)D����� '
�|�q ���c��7�S�p���nyoT�a%U�3��)+��&����N��U�S)j�ٮ�(B�9��=�l��;�DPn���	K%�ϧ�����U��f�`.[��N2�%]�
a*9�6��zȁ�9��{��JHF�3���,G�tI��n����o��eĳ�����JU�����-�cGH�`��9������X���Q�>������,�(4�J���({�#Fg1b�n��O�=��3�7�d��Y� s��x���@���r�t,�Z�u& �	��m�r�o}���ɿC[g�'����9��sķo�#�q3���&S�_�h�[/C�ņ_�L�aU��R=���(b�-�T��n�և(��L����5���_=��W��6�[U��4n�l0ĺ�6/�����翄����?�iFO���B3�C��ܚ9��&��}8[��\�"��w��F�QD֟~G{�q^*le]^]T�ҫ�}�y9H_.h�m.c
��b0���m�$��'xwx�̚�]Sٙ��x�-���m�Ӆo��_���r�)�ݹ��u��y1����G�1vY��W��[v]mT�����{�i��@�k8�����$����֐����>�wᏥ�7o��T b������]��
��%׊c�C ]�� )D�F\�<� �3!o<R ��s`A�<��y��>���T�����J����6y�8�6|]��&�mb｝K'�yP�õJ�!=q9P�������s�(Ҡ4Z�,p|��#ڌȿ�x���J��B9�F`�)J��s�!x�D1$�M^��W�7�1Z0�n�2�"�^e��}R� ?Ԥ�M��8���C���g�m"vn����������&�$&SQ<`m8�(�6��k��{}R[WUi��#T�=�d�3G�9ĉ{O�qx�٤�~tⱼ������ҮR�L�	��c�KL]{�>G�WR��!�G$D�%��7~������|���=��'y�s���O���w&h5���I�R�(��~�4RuX���Ȱ���x��������}���F�)B*_��`>M�tਫ਼�����ͣ�%\����]���f�fs�.�{�IN߇!^�u��u��>\�(Mj��k_���|��� n��#��;���y߃l�w��7��������|mB�5]Bk5�K¢�}� ���l��{��+��I�}tD�;��� ��������ǡ�١��D��:Q'�P�>uOHa.ک�&���`K�BE4�ً���Ǟx�e�
������+(�gtڄ���U�^�ʅs�koݜ	q��@��JQ n�������sث׸��_��c���,�M�Q4-~+K[I����0��~�)�س9&/Pӂj�f9L�69��Omn����%����ƣ�D�,ށ�!{^�8"d�j�ޅ(�+<��q�|��﹟��u�/~�[��G�.��F\��9yflD)"Z �>"�J���(՟�����p�����ܺx��[wB�"ݹG��a����j��E����5��X��*B6���*�x�M�6�1�s��-�t�7��/�/�L~s̱'��=���m0q��Q��~�^)�v-��.�"KF����a�L>Ef7x�+���6����Sl��8-�J��J�[j/+"�qo�s�,�}g�ΙSlڂ?�	���_�N��ɩ�A'X/06̩���BT��_��p�x�+�\�<C ����I�²1��^���7��>u���O��鄘3�����������uF_�H>�R�Ei�s!Y�m��=���~�ZB��b%�ύVj���w��*5��o��bl[�W�T�몗�ή�|}����]���8�_��4*IpiB�������c��%67L�c��������R�:�N������i�{�H�``��<��A���T
��7q7o2���|d��6���w}S�k�/2�@��1	 �P������,VE��67^���=��#�YA����R��YH�4��.Q��Z�}�~�ͳ�Q�Mf���op���O<���7��#���d��L�s�6^��u�.�ܫ�O��]R��#Ak�f2dd%����I Tj�|�u�����5K�#��Q�B��}WG�]Ｊ�ߙ��J��!� �ӽ1�T���������9a�+�}�r���fbU�?�w�����b>�N���h v���6��ˈ�ap�nN�c�#�VeJ�p��J�����Jk�U�D�z?�@a9���=vo^G`,5ɑ�Ἒ�^��o�U�Tg��;uƱ[��fd=u��1Γj��Kor���wI�F��x�pem¥�5iF�aZ���x�o��gEpo���]���)��#�2�<XH���HF��t�"�4M�{^ |P~k��HC(�PA%#Ps�ĶhLC�!cQ��:$-\�
�A�i��x�!C�R�!,�<]D!c�\��&��^� @���'@"��eDC�s��E����ч�_�����G���HH�SQ`��XA�$���<�q�S���\�	��q�uFi�F'�x�*\�� ��X�Q&�H�є�%�I���������1���J�s%��(!1!�Y���̿��CZ���k�k�>�g��m-�b��hw��s=��8!W3.&�����c"��s�/}��J#&�0ÒF����2^�"s��_6�$9x�pGZ�T�C$�鐋w��}g��O�;��/��K?�!Z;�l�aD�@>�P�6��X H��!Ŧ�xi����L����(�f&3`�� ����E���W� 4|�=`C��=3�F�"�(�p�Σ�Q��A��!�9l��V�-��I�#,FX	K��T��q��^��(��@%�u��Q��V�|�*r4�L��x���ZQ�R^&Q��<'x��~���
Bx�O���&��1&�D��L	2� \�pq�sW�$wx�W(#�t%zPB�n�ǎ!���˯�9;��3N�9|��O�ͭ�%4�\c��=��#��}�R�*�\�3�6T��^�4F1����I����rm������v
w�I6�9����:�$���|�W1�(k�B-��"l^*b���i҃���ք(5���W��+/��#���&�^��df���il�AVL!�a2x�ؽQx\r�W�J���ґ�+	Zέ��,iA���h�%�B�
��I��� �>����!ǀ�$)Q��f�<��[�t�9��"h�|e��J�W�!��"�q�����>(�����_V�sdTI��E�ǕvI����/��ԈB݂�Ug�w-�zu�ȶ���_߇S)�pH/�:�(�X�D��1+J)t#TDQ�1�#���5�u��M��T�B�F*�����ǚ�2t�0:�ة3<��Sl�P��0�p��
���a�F�����6�{��UE�õ"s9&�!,�rꁇ�؝l�s��K�^����H��Q���3�^"�g-a�'R��:{�#}�A>��_���S�1���_�k�l�u=X�4���ۛqaS+�92�)��0�1��ʉb�y�~Pɿ!)Vhk~�i��\o�V�%��`!~[AQI��Uuj�W_���#e� �Ϭ{C�G�0�`K�4�j��rm��k���[�S�KWx�_E��G����{���1�ͣ%2E����"���՚A �BP+�f6!�y���+�)���Ü�Я��:�n1��)�T�x�l<Ca��l��Jr���a��{����kI�\~���^�8y������(�y��^H~.�����u�U�����(F	�@�DN0��Ę�ȗ��tJ"#�Lc�5D�H���������RJ���i�Ь7���6���㝎9���j�4p�X�_}ʃ�z�7T��]mP���w�T]P��ڄ�>�U���	2����5�wdɀ�=���	
�0&�0���2W{�O�c��#��U<NϢ�JbT�h� ��,r�8j��	W��~����G��U1�h�[[��6�;��~0^U��D�'�$���܀c=Α�ũ=�c��96�c2
�v��^c�%�ed�c�C��M�w�l�ru����r�ϒk�.p`��`6&���f�1��X���"����H�0yA6��*&Mc�0HY ʀ6}Ġ�}A��SbS�D�?�zV�N�WK_[8-\��T�6����(�e��)Z*ֆ�DQBf-f��_����^���oD���\��W����`���D��e�D�Q�@	��x��.D�,����9���l���O���շ�i���8�}g�)�0h<��ܡE�;���eW9�꼂�;Z�h�yƕs/r�G?d|�����C�sK�<*�qX�a]�	}n��S�L�X�}�6�gd��������"��~���yw0�t'd���^�D9�v&��c�Lp73�K����/�3�+������aT��UD~A���.h²��v?7 ������R}��@�|���d�:�e�ߢ�^���6TW�i�C�X�"�1�d�Q�<���"��@I�t�to� �"�����2�Y����,��Z��U�9��&R��7�!B>�83�8cv�"����h�B�|����ݑ�l�o�v[�x�w-��)(lN��l��N2��Hin��2���10�|b�3��,Y��9ܪ�X(
鉣��y��IG�sɡ��r��>��,�O���/�ĥo�#Q��g��+а�M炭�d�I�X뙭�߈�:
�ٙ�[O��ɠ���:�����O� Ј���O�k���m�_����7WI�#)S��Q�p!��L�%Y�D	�Q���gB:2?���_X�5mx�ā��]��|��������8���2�8�N.'3S�R���+�}�EB�,�$�f��~�~��=uu�F�D��c�8BF��zw0�f4���'�w��UOaBIt��l�hz��8BDd�5��&cJ!��8R4c���6�_%അ�:c��88O���cI~��~�sf;{�����~�5�TX������r���~4�x�.{�u�Sj�Uˠ������[�.=-SM��,���!�r�P����k��U��\��W�^��3�:��,��{1��4�`��}0.2R	~ga2��D*�9Gn�F��2�/ݿj�<�V���V��j�ԸC-�Ŭ��cZ�S�?�$X�!f{����,��g3��T7�oU��|a���~��Ǩ5�	�oe�0���wq����S�}�W��-��YO��J�3�r���\�6d�a.�@�<ϑf�Ipm���Ȅ��$�<����u.~�;�M'��%I��iI�-�H8_���O`l�R���+��β�Sn%��m���U�����ZյHC���p�!��CHSF� r�AH3��Q������0��(��ˋʐ+��ȧFD�x�m��#L�������8�:]��ud�˖?K&�9�����R��-^�ǿ�\��^[��G>�ُ~�b�0�VH�GQ�G5l�U"d���`C"A\��������z�$��;?骎���t�L�1�0 � A��YJ�6$qcC|R�bc�u���Pl(Vk�Ii)�A��0��oo�ǔI�YU�N�:�6HnvT�����������:����<�U6N�%�#%J�����ݥ�}{�gm}�a�w�=.��c4c-��|����9.>�<N�x�H�-V�g�9딪�y���m�|��s��JL"p{׹��O�wva��0��AI"�ԍ .|@u<�널�y����W���{DZ�^�bA��ߚ{#����u�N�X�a���o������ꇄ�4�NjM�b���Q�]��r�iJ_C��%��d�[�3��|X���D��FXa�Dg{�~��fx�(�!tģ�!,����#��k�;��v�>�XĆVhbx���Ïq����3�7����\��8�    IDAT+-F&c��ͷ�|�-I��"�roA3&�IM�P�>0�x��ș'g,�۟1��mt�㼊��E$�R�R�V5�@�%H(�x﹝����\x��p���?f��[�>�w
����;�y����h�&
�	C&Ӏ��<������9��/�'�ԝu�K�V�<Tվ:H`��6s��O�S�j��D���B�1o7}1KV�'mA@J�֚a���W�w�~�_c���\m��[v�t!��<��Y�K��19`��,���R|�&~r��Θ���k�ؕ��T�����{Hs���Q��%Gb'����x���SO����Oq�9t�HS�D������~�}�{�AV	c�{�����>x����%&{S�>��z�K�jݠm{03?�q.~�����u�Fxk�bi��B��;er�Sd	�;-)� /le���-JBي/��m����m�Ro����U�׌�B�Jd��f�}|�^�;��^�L���v��J4ldbre�Ir!�����`�ô��s��к�t%���ޡ������ii�B���&�~�O^�)�����Be�Ҝ��TĦ�K��m���%���8�2(
A���g�"7�̲;ȫ7���L���e4�yق�]G�ݶҷ{d����GZȝ'����S�B���u>��������r/!�x;ŕs�b���J�R!�N�0;�f@���s�Γgw��e����2��7�E�"B��8kK��Ih�KJ,^D*�CBq�~N|��x�����ɯr���q�2j��k}�ty���d+�C��X!��a����k�z�2XK�v�ߵ��)UUf���i�����o�/�+/����ӿ��L��bόc4zK3�[7]Y��v��MH�
M�5��%7^�	[2�=Kr�s�kC�y���Z�a2�a� R�xQ���[�~�&�sm�z�Y�#Ǚ�bU8!��9�g���8-�c��& ����^1����5n~�>))��M���R����W,������=ڭ�ƅ�w���Ԉ2@��b:'����A0��1NH���B����r�p�U�M������A7���n�B#8��[��d�y!��(�("���{9��-cE$�v�SJ-����51�BS$�v�ﾴ>�LW�i��s�5B@Y�ڰ1� ����׹��$SS��JJk+-h!l4����[<��pl����C��J�Ԋ2V�nn�8����ĵ�>�}Q:�,� �a/Co�n�gH�_X���y@)�
�%&`vv�<���]�;�x��ELw$)s+@jD���b8�Z
����@jf�_EY����;w������9��6�_̙�BaI�]w�l=õ�x���� �Ђ����7����/IN�b>�P�Z����w}�{�#��h��&�@0_�x�������r���W�U��1�_��"�ʆV&���V$�b����bb��x���[�;Ͼ���m��ak&ҮV�Q��˷R
!1�R)Lȹ���L_��r�>��Ϟ!M�(!���D=��N�4��3ʬ@(E�Ǩ��Md9�X3K��UN?�89%E>C�V����1��q�>b��w��TK�pR�0����mL�(
/H�!�yּ��$+��Y�i��RsH���-�3Kb:�L7�MN�>��c�р�%^	�
�T���E��<a]����8]�]���ݬ�6��A�N��׽�n��kZ��d����ϵ�C���DX�>��M�k������`��P(��h�AH��4%�#�T�a�-��&� �z�q�T��|@i��ǼQg�[��є���:���#s���;�rN��1��	�)�!��-��-F�!E���d��RvDdX:�d,��|@�z�� � 	D�HP�"R�\B�"�=HO4�W�y�47W�#V0����,�6����O_A_���Jq��!�܀T(�Ϛȁ�E�x� ĺ��h QB��zΩ�SB4��`�@di(���v�y�[�I�a��I殰�MI�cv˂a��}$c�O�~�)����~0E�U3G1��dꎲ��י����O���wAc��˒��C��bci�I)A-� ��"����m)81<��t��/�����a��f�ὗ��wC�=E.b b��Q�`�{�hT�L�1(�Ρ�Ya��u���%b}�%�r�U��O�@>���� ���)�I��y��� 6� ؼ� +RVu�Z��Pa��K��ȧ����Gĵw��	��M�g��?��Zñ�a3sX	�p�0�tٸ�$X��� 8�A�}�(�[�[�Nl�G\}���m������q�/rEiv�g0�QCf��`� Ʌ%��'n�lE�$����;�s�e1)rx��8�0#MA�,܇m��fu0�se�P���AJO��ݶ��d�
�Rbf��(�Kfh����f��0e��3_d���k�x3&Iv(�	�*ȫ>DG�oec�>/���@L��Z��D@ƺ"A��[N�q.��T)��!G��=d|"'�7�#�:�0��%��R�֠�)��@�y�t�b$��+��-���q�D)��	ZF�
U�<����@J�(J)"Р��8�P�P*+!���sD��	�h]	�>�=�P�:"+�`E�ģm�KJR�J���5ٳPm��V���D�Nk���0�յv���ܧ���B�ƚ��g-��ɀ,˘�S��H-�;��S�����*�(�k���zq,�i̻5z�X>*���D�Ek���{iW(��&�JD: ���֢M��6�x�;���:B�g�i��!v�`L�#eD�2*eg�$=�4��tF���yN(m���eڮ�Nb�P�����'y����ęS�^����1�rY(�0J`�m"w�$��5�5���x��*04C)ߞ1lq��O�>p���M^���c��Wi��V�T%#i���(P��\]���R�˶i�~7+.={���o��;�q�\Z�봶�bS��������S�N��ڲ}�_����=v�OO6T�Cb���b>�X�dB �l [CY����^������1eN���O����9�Ԕ�}\�a;�|�9"��sU����%��o�������;3��ǜ>�|��[N�B�ʃ���aֻ�����U��$IH�F��>i�z�6A�?u����C)I"4���~Fz-m�Y�:t���q�Uø�,dd=P7�p�ǯv���m�s��h��d6���QHuX�Y�5�]��ig��S��!�Bm]����As�ݛ�9�*|�z��ܤ���k�S6y�s��k�{w"���3/-u��y}�f�C�;ˋ�۷���Xځ��#M�Q���jT� w�8��c���˦���c��ݬI�H�c��-�p��#z,� ��[}oD5s�3g��(I*5s��G�8I��8�ݽ��z�.Zr�-�Y���LD]"����;k�QT���<oN���^��`�I>�1��}������C�����a�6�QQY���s����9�ŋ`<��~��/��E� �Yt*dDm\1�u���l� �h3d���g�����G�1-���\��?'��91�H�~�{Tr�V��MQ�Hc�!$�S
� �X���6��]���f�r�_\�o`M!,�b��U��d��5Ԥv���G|��������J����o~��G����Ҕ�,�S�6�!Y6�m� PV)ODk�􎑑��.W~�C�K��P�}��G�ǩ���`�,о�'�|�H)�P�I �����з��bș/~��'!���]�~�����������{2΍���9ʛ��{�&�Ol����|Dz�)�H?��)mf�.��=�>o(s_0K���p�������3J,�dHY���2��F����f��`���?��J)� �C��E�2���ǧ���*�j���}�n��;4e�z�5é����Y�#�=Ob< "���Y�C���>�sP����E쁁�e֑9�O>I�Z��%�I�J���Md���ih1B�9cQ�n3m/���7��+{�O'"?8O@PŃ_z����0�\1A���W%5�Xd��+ʘ=�y7������w����/$��Q�!���I��%av��ｇ��RB��_豴F�@��Qc6�?�C��v��c��d��1L�%���r����XK Oa3����;�6|�p�W~��AN������+�n�`,S��$�����`�?��n�R!��tw��A�m�[�����C-l��������H_�uh������nv�k��d/����.J�����y���3ӛ8�H�)s����ĭ]W��������&�M�ѷ�����-Jf�c�<��d��iLmꉦU���6�K�c%(��?A�!G.~�?B�������1|�~Z�
��7�5R�{7���Op�� ��i��0h�Rd�����_�pb�?�� }������n�"���i+ <���iK?*^��R���:,_�ފ�����S[�,��ݹ���m5w���mP����~��t�=j�t�Knb!�4��Π�ڝ�vk��D�mί�i��!�,rc���Xk
G��.Ǘ�a̋�>�y.�ƔB���R�T�Z=�y��&_��{A��iw�v3�RؒR��.�C�7�!��7�S���t��J��L�d%enu~C��2"�:��^_n黅��9Ǥ�IN���_���1:����bJ"*�6�qu��)B��v������׾F�|�^"�3�3� -#�
!V�+]3���E�|:����ǜ|��x�[�̝���q���Wy�������-�I(,��[k�q��N,�T�RJ��Yg��(���U��A�F�^�:�P��F�:�}�.ϸ��"6��.��o������ٔ������G�}��b��F2��"�rp�]�Mi���<BJJ瘗��$��Ə�=�G&���|�����zQ��`8��t�}̨���ZG%�,&���g|��+��Qd��-�$��k�1��� Z*�C�J,��5�e�#��b�8�y�w���c��|�n�����5��=��C?@����t@���>��*vD�]��`E �!�C+�r��V�J�(�{�|fitǻ��ْ0Q׺��dr����ܓ5�$$i���R���.a�����S�v��(˺��'��e$Ū��m
-��:�B@%E���1�ӈd�3,I�1�u����V��H��}�a�`�8�x�﯊^�U�_���]J=�S �S�"j^j4�H� IAq�2�(P�&��߷�̋X,�)�Ojm���X
�qcwa�\�B��n�FtF�M� غx�����ѐ��en��C݊_���X&}k�M<=%�N�b5��|�٤��O~Ļ�}��X,�$Z
����k�
���gcs�������<�c��u�.�g�J�_��������li�������a�5#�ZSzGVx��䮤�!h����jT]V��nV�2������`���l�O�'���CMy���q�����o�-���}������sub�A�#5#�V���YM& '<�� �&T ����v�}�ro�p�8�|��̷��iE�M�{�.!��\��%Zj��y����\��a��m �>Er�~r/p~~���?��ۿ�(��"�v�%ER��&�;W@Hv�~�SO�@n�Z���F�g�[���흃���;Z�h4��hu�<��s}?����ٴ�zI��ൾ{���N�[��A����^����t��m���ճ��|��&��
�!���Ж�]_�A�c�}i:X�,��e??��&i��^��b�$.��g%�(L:�C	�=ʽ;�R�h4���j���zBҷ�Ѕ'�Li�գ��ʂ���h��!^k����ϥW~L��"`FY"\�sK-PR��ti��Ϻ���vm�Qk�AD�TP�%�i�
�;X=��ϸ��|��0���@$*β�C6~��}�&��Ǟx��>.g�w����b;6����^x��R~�,A���;�};ESf�g�ǜ|�Kl>�(�+��2y�\}���?��|��)Rl4�+j5V,!�F��Fh�u&E��	O���[�;��wJ|��T���Ž��=�}�#�'.C͆�B���On���+\��f��w��?�y.~����9ؤK�8���ʸ����h
mi��.}�'/}�d�Ji�.N�e?j�<�]IB���/YybE1b��:vRI�y�٥�щ���p���ǢX._���?�:_7�J���V�N�
��܍�|���b��l��0��b`��E���x]����a}���3W��p8J���
��a2!
�?���9&"��;P� ,��u�T����6�U߹��P�(|}�o�ƌ��kd�OP����m2v0���f��A�~ͩ����� �~��VM*���[��^Z���/�*�1H)1j@�9r��h�Fb����\��#lsns[��y��B�op���^�W`V}�u�~X5�����y����NI�`r�&��+hb �oR��A�27�v�B��w������J꒝JQV�B�G�Q8����]����#�2��� Ix�0yn��<��W8����"�ꛯs��W��)a�
�pi=�t�h4�X��Ԍ{d�+���{���|���/������ǆ�Ǆ0���F1�4�i4�E�B �$I���mQ�"�|�I�"��z�ᶠ���u�{��H��)�m���=�L'B�ؑBLJB�Ē�psr�r0�����?��d�L�<���x�_�0C���\�^�})0J���!,x�w�Rr�w�\��,��N������6�|e��9�Zb���j���j� ŉ��0�|��~�2���:��yҔ��*@�c��h�J*18��U�R�0�e~���2�w����y�\�P!�I��=���4��~��x��_�P0�s�r�bF������pw���"����ג�,>��HŊ寫��j�-��:���k}��t�o�����6O���M�F�Te8#4�GJ��Y�
�*?Y�=��B�@ ��*2&U�Q������"�ȅ���"�R*������$��Q�D"t�:�3 �BJ����"H��>���(�D����q�˚.�߽�-��Wp�s�&�A��쥟���ƒB
FN�m<6d�S��b���
��"�B���j�4�\M��.4y�h�r�g)���+��`�^=��w�e�<r[��ȡd�_c�2��M$�
pH�(mV��h�(��m�l�Rl��s��ޮ�`2RE,ZIR�b�N=�􃏱u�n�9�ܣ�{��QJ�L�S�rW��2�R���M�Z����^"(xJD�)���d�h�4���$��$��'�����.��f�5"H�W�4a��,gCD�@X�2�U
�4>@i�v�A�m2u�_d�s�����|��~�?!߾E�,�p�JRr�:C�(��YRmH���%���=����Y6��>oQnJ�K�Q8Pz�P�ҫ�uH
�V1��v��@M�q�T"]��+�Q"6�,���A{Ű����ܗ�D�he�W��e�zI	�;�����=e�H�*<[�����v�Ý���i�c�e�+g$Y�N�\dO@V�"��8� 4����a��ܳ"9��q��O�'��)��8�M`w|��dW8�Ԅ �֑(I�%��+�B�F���R��#�!��&���$-�dh6�1ߧ��\V�DF<f�T��; F]��VX��-��1����dR
��,L)�"�RϦ���	����8p�l��<���ZA)��AYх$��E��d��.��V�}n)Z����H`|ms���?���-� �{��ws�x�D:�הJ�"��꺷?;B�g4��Tq��#�!("\zPiB#��Uf�GV|."Jh���U�7��&�b>��q}T8)13�R|k�{e��B��@+��=b`0B#\���d�E�Uɼ�s/Gw���.��s�徇����h�d��?K)�b4��&MS�N D� !,���;ѫ���bR��K=w�z�������7Ʌ"'�˂a�Ѕ���~���gi瘪N�j��ޔ�t�0/rL�R��t�p��y�,��I�    IDAT=�(�z��l�x �߸�P:���l�?�N�̢X�̤"٢���rF�#���<g�5(FJ�e�ظx��>���QŔ��������ɋ��U�{4�sXׁ��֒�9d)3�r[���)"����E�V;o�1�k����m{���.b��u`>���A�P	�
�����E[K�/���_�?�?���.�4�ع�9��s��-
UR�%޺��;0��p������7~����X'�>Ϲ'�g"v�QS��9GĸP+4�۔�tBZX�|FP�m3x�4�e�k1;�ʹ�]�>�}�Nˬ߹Ԋ��cnOf��%��1�����:����{��Ż�J��cq!��|�%j`H7��Db�HZ��kW}���_7o�������.F��u]�������:˰se� �葉�9A�7�67l��՟�G{��^�a���#ۻ�5�t��.Cꛜ���'�A �&M�hm✕��RV~��0׍�o�����6���xa%�^�V	���t���I��e Y�-1z-��0��1]#�����:#�4L�k�؛O�~�*y�a��ٹ��"/g�?����fXi�}�4��\h�G�DA���3�=ǩ�!�����>�ĶR1Eh���k�=��i���a�H�\��W9���$�"n_�x���	B�
/!jl�E�\$��쪟�E�N���JnKd^ ��D�Րm�2�00 G�w���]WA+� \,;���y���G���Ec�l�s�����mrB�8�����|���-��y��_�E��#�U�z�Ui;u�N��C��wSF2���b�:����\���ak��LU��!�� K�fkk�P�sF��{�ٕ���1�p���z�L %@ڿ������\��ꮹ�q��}J�}f���%OQd�)�zA���+W�R�.�����R�dG�術��+�h����҅�*2z�txb`��S:[��cu���~�meQ4�hRʕT��o�� O�=���-}�}W���A�v����Y(/Rj��|�mf��t������Lb�����m\�E.�2Aj��>�L@��t?ǀ�LP!��	g��d1}��Z.!���t��W��ۚT)�;�y'�2w��6�}��!M'S\V,��;�Yw>z~��`;uk�ag�5��I�S*��!G�?�3�=��O<Ά1�̑nn3�������1�z#$Ey�����s}�=O!Gy�ϳq�(��y�/���ǟ�
��6ź5���/>�����j/<�sG�}�SO>�L@>���������q���HM"�+�/P4� J/�%J)Bq��4�:��r��x7Ż���bxػ�j{}m�+���$��-��X�`�N̔i"U̾'�y�(_0�{�7���_�DF����l<�(S%�F'����c�� ?��\Ok3��{�D����"�(Ԉ�3�	�`Ii�i���ޖ���s����)�;�>������.f�'�2��Pj�kau�������ٗ�T*�x����9~�!N~�I��9�0!5�1}�d�������ںiQ�B/+W2Tk��Y��>���EU��y	O�A��Z�r���w����FL�^��'�)!��1Ƨ�察e�]2I��t_�)�g�[�/~�3�$�&ǺÈ���1�F ��5�,%yWFM:�4�5&�N?�����PT���[��h�m��l�t
�}��=�̕XW���I�hL��|��	�{�w��߻��Q�,�eI �|��D ����x��>�h4b��.�._��'S��1H�,�֊�� �9J�ذ!�'��s��L��Zt���GOP��]���*�f$���e����ɽg���;��'>�%��y��wnp��1)'X/[P�� �\�_� !%Jk6�	��j�ޑ\���RjȂf�'k1��v/��9������>��A%\�pK���H��h��Ϫ�j	L"[���|5�R[��v��&w��}��/~���f��^�Wd�N+���KD=�{A�{�~�׈�h)� ����@i>P�r���Q��0� "��`@�w�[ｍ����p�$�V�R+�saFj8����{��n��߭/�����>�ͫ�����s��3c�\�[����M?Z��1�uL��� 	A�bL^��� �
�F����h�/ �ˣ�3���>{�_m{_�Z�-����[i�3����K�޾��7x�w�" ˼��6y�S}��?�%�]���Hl��>��_�.��Z���kYp�U%	V���w���(�����=�{߀��p/s�(���V-� B�%4V�`HQl$9�'�V��ܦ-��|�G�|b�kM����>�$᳏>�W^��w���ի���ź�t�0H�$c����໨T�G�k�Z� |��Gℤ�'4s��Ot>%ѱ���M|X�t5�o��>�޻GRZϑ��7	��0��ob�n!�	$�W�ߢN�Ԃ.���hV�����w��O������?����S��S�Ze��t��>m�nG�[�Y�n!8���s�W��GNrm. ��P��5h�H��j��f�V����6C�����v'@���}�	0�.���R�0Q��"�.v�n6(\�����1��Gh_ �[��Nkr�_[��)�r�R�E'�� ��9[ڀ���U p�����4����ۺ��������]���#D6Ë�y=���F�;�η�����X �h��J�TY;u�,�#<1��� w.BWkRc{��{��Ϫ�*�n�u��}�D�%kj�-�"
˫�����=�� @D�5J9�'��@I%��,	)!L�.�?��t6ԃ\.pP�.�����w��7!�?PV�_�c�N�QW�DU�Mp�f,�_�!��D��D,�")P��Ɩ���Pf�_�D�O�|�M�����};HKl׮���oIJ����	W������lʄc��l�҄�9Fmn!�����q���Q�+}j��+�A�*78u�4ag�~6A���e̊��h��ځmB�X��X�Sngt�~n�	��������ݿ�q�ܛ�@�z׵�E��}~m<z�N���_����.���ȗ�����昫���x��۝��ˮ� V߫ġ�!��W~���Ϳ����l��>��:ƥF�l�Pi�]Сv_%�D%��&x.�����C�)vv���/�6�x+�*��+!][�Z�vŌT�l���K?�!���l��?�pg�·��7~캚�����b@�+-Ӽ@�Ău�rp�-��+�Y]]�k���_}f�uB[����g2�p��w�9J&6����D+�h8<T������,B@�'�ʪ�*���%��L]�����m
)�u}_�_�[}���m�r����@����9-X]!��������כ��=W�+K��{;�����^�횉�Ei3ضo��ݏ�.�}~���_�ׅ�)��ٶJNV���,
ݱ�C���T�@��{s�#|`s{�$I%)��_����h�}7���8����u�Yp-F���#���.c�Iܢ����]��;��@�,�!R�$��Q�k�,,s�'��E��׿��sg	Zr��gX�#L����dw�	2@�$P8rk=`SMy�fﾅ+�H
K^V\^t߷�ݰ����F�_�џ�<� H�&�{w����>�(Ѻ�꾫���^'��"���X�안�S<�����+�߷��<� P]7J�r?�x�$#����8��{�Q���vN�г/�q�(f<�W@U�tZ��l�&h���9�l��e����������O��.>����ft+�a���u��B[;�͸ލ�{K�gxe�9w���?���n<�a{� ��ǐڭo?�i�RJ�	~2�Oge�f��[.������Gi���+�.k"��qe�-�|�8~��ΟE�R��X뱅ède�梫��U��������v�ƿՂo�3V�ӟ��}�}�	2����FR�{��� �`ʮ
rX�6P:�:�@=�
�"���"qx%:"���#58��3�!��G�*��BE	[�X�^�oI�n�%�dE�㘜��;/|^5�G}�'x�u�dC��=��� ���v�C�U�w�
�,sUI	"�C��dD�
���k��9�Kuz�\���ʞwoA�Ҡ5吉(�>q{|�K&��W^�	�� �T��n	X�5���������uO��R-��BA��v���Pr[r�0v��K��~�~�l;E�2w��1'1n����� ���2�!0BRj�P9�� �D��4��S��^�����.#a ��e�`�9�i���d,8S��p�b��g�Y�'_�_�wt�}�����z�cN�e�` ���U	��5L�B!��(�<�Ch�0�&d�g�H��9��
'��cs���Wx�����ΊM�Y�JRP����K��"Ȁ�����"-6�
?Cct
R₈�C(���XMH��������}�(6�}��~�_p��ܵ��$C�H���<#����`��vU[����ۜL���W��|�-�,C�?���#���9j�8�'��h\у�"�ZJL��Sl'�b���>�tJ�~ã6Ƙ|�(�칀)�S8��k���ItP(/	l.�Dl�:��[�l���gƈ�K�I��nJ�����Aļi���̈
����
�[6n�g7F�a�a	3#��D��]HGr�;�-�p�w�M5ʗ�Ļ�akQ�)��F!���T�z���:�o�s7��	ň�X�W�M�	lL����_A_����Cl>�"�/�	�V3���M�|�2i�#��j\%�ǌ��\�;�8,�+"������"ӶnJl)�V<
�" dB���5�
�u�Ʋ�8\ۅ�o�E�.z����=B�:G�%e��T�0
4>&� �cI[B@K����-�蘦�����;�E&Qko=)���v�#I!��~�u�.=�-5U0�"��/nm)��uM@J�X	b�w�s�}�ο
�0A��Ã��O��EE0�k��6��f�{��u� KL��,�Uߏ7woE�	sSwm��{��6GN�A�	�@>ۥ�ܥte�x��8�{�ΛW��x�V� %��l١t׮]������ah�ͮך�1�!I��Z�p��\|�)6��+W���7���,"pF��nYi9v�8�K�����[�c�ϒmJ6����~���['��Y��e��v�h��r����+<J� �HH�Y\�Ʌgc�����k�g��s�����s.~��월R�l��
d]I�X�t׎�c����|��%ds4�,w�'��r�x��+f�)�9L�����KOń�s�
��b EV�t�0�bA�|�ay>��g�JJ�('�&\����]�2��$*#�c�"Z����F%+�r��v��Zf�~o�k�ⶵn(��1����e�L��D�U�om>P&}sҧ��}iO|V�(.��(�)�o^c>�!D$I)%eYRι��ܧՅn_�ͱ#➴[�|�5V!JjK�j[;�׭���v��a�;�4�5�9m�w��i�|N��'iB}��)��<�܅ ��^���CG �;�Q�}׶�#�!C堗!�9\1�����꠼:�(�:~�A�<tJw.��T&�#Z5��Z�D(	�w��@x?f���S�����:%�-0�����y�x�/r�G�[�̕��#�NQj�2�y�MQ2P�XX&��@�z��M���W(�B�H���M�h��%����Ŝ��*��
�X�+�_�0E�����I�0ۛq��w��'/�-$&�(#�#r����f4H��N���l~�󈡧��u�|����lF��!;����ʁ_%�-��:һq�G�-�ڃE-j�p�^�36��!��������_v���n���_�gy�r�#�&�J!1=�~_�H�6�/,1=�t$�d�����\�ǜ|�E��-%y�B�ʹFh�c2��6j�>�|�t9r6A��>v�앞YQ��A��ф�k�k�

%0R1�˸����.r���a���d�;G"UcMjӁØv��A֋5�Lw�Hr�=�v�������IY�7�G�ۊ%����󽶾k��G�Q�l���M�H�0HG�6
�T1���0��}v�Na��ܚGAQ���+\{l�XXz���
^�^!�&�V��s?�]���e�N�}�r]�ߝ�����b�]�S�y1�������|M��L�ҳD���Q���.�l�ͮ�P�ڬ�J��Dm��l}Ԁ7}�G8a� ũ�z�X���h���d R!���3�-#���-$�.�n��nVC����:�ar�����W�|Fb��y���݇U
�l���N�r�71�	CSU�
r�ɷ[#TV�ƻ�bZ����H-��a�G	�@��)�]��BQ�'V�BȄ)�0:B!c
��}{�#	�z��Į���7�2��l�@���Γ���<�4[�;�k�y�������`dȊ�b2C�fK̽o�t-,��ki�B�җ���!H��	�t�lZ�a�;Wy���+/��i�Ȏ����_⮅4M���FI�X�,�
�E�HT��Dy;��;o�w�
&p��'8��x��&�
fW�KOq��.�9D����K\�ǭ��#�~�A����9�`�l�7?!Dk���=;M�XD�V�2��]�$�J�(E QI�K������D��\��s�:����]�' �gZXPW��
Ǳsr��g`�0�sYe��i�Rj�v�!�S�{�}�rQ�iq�ų*-W�r(+�_�Rϫk�8皌�z��5�1����_�I�@̨P��9bx
�����s�=+�JK�Y�?�&�?��>���D��������Cn_[_���V�[����:6����׾���W����*�#�u(-���!Kc󫮄�D�0� ���b�5�o3��wJ���	"�u��*���*Ӥh��	��$0T9� ��`3U	���ɷ�>��t�`{��ZP�ItQ�����'q����v�=s��Q�T$J2�}��^y�?!���T������a���\N�D�}_�b���fs�,�,]5�Ք���/c,@���!�(��`��̰��;J�"���������)(�%�dN⏜�_�5����9ӗ^b�G��@Iz|��
a�u�F;��W���J U UB@�}�1�(@�C@%G�*-�Q���'|�_��y�\�<��]�a8E Wzd�K�p$�X�)z��\{�u.��6�9��w�?���W�$������̪��m�z��{zzf�!gH��H��!S�˂ ��?�?�˰%@HK��$�
�Y؜����o���23"�8�YYYY���� �[Kf�z��=k� ��S*�9��VW;/%Z^�ޅfs[��������?����=����ǫo�Mr�P4�C�:������H����RR�P9���w�{!�`X�j� m9��^F����V.����˃�kG�q��r���
���6�&�?=��2��Q�z�2Z���}�� <��pv��֫�S�x�lO9ҧ2��kޅ��E�=7��d��*����r)ݡ6,��0 4���3F��	SzN�;���fN:=���)1�7(�s�sv���3� p�"0in�����}&��w�3�m��L��9������Ԗ�)�ÐUV8��IDEѪb(�K.HN��|S=X7�%ȋ$�!g�r����J�*υ�����S����R�;�ϸ��#֓�m���9�*�U��B���ʊ9�]�7ׂo��4L�~i^20dE�2�������-^��o��-��	��h�@t�+������|nsT\��h�����.����x�7y������O>%Da�t��D��k��[��i�$�7�(��C9La�4tWV!�[��Rb��q���­��Η�����H<~S!bۑ�<hR����g�-�s&J�	��)��?�v�
�~���9�s��	��"�{�!jm�[���A�UTU��+W�|��g��Zq������*��*XA+E=T컙�����Ͼm4�#\�y��k�b���q���/jK�u�O�*< ut���O�ٱW!�*\�-(�#�ix�Ppe������0sS��Us�q��&��~[�����1�?qZ��y)�    IDAT#�Wc:X/f�9���7�`���0�;�ܻ�p*�����I��<�oN�q&�蜆6�Ԇڌ}��P�Ԗ��#B� q9�8e����)<�t�G͹��.
x[��ܓ��� ��u�'�v�<����KD��ܗch|:���9V��N xrI`}�G=��O��9�s��?��]U���w"$q��Z�x�}d�o���Q���Ჲ�j�d���b�X��o5��#R��R�	�%H@��[�*M�F�'�'	��`_� bN)��]y흯����N%䧏�>fUhb���۫��`h밢��8�p���&���l�\�Җ��}v�~Ȧj����mF�.��S���M�D�PCc(��,�LF,<�D�'�t�٬jv�S��A�m[�}�	������g)��_G��e�*��uE^��|�#�
�8!;O]6��ὢ���}:h5�:%���"&�f���,H��P	T}G�9��BG��X���v����pIٸꀳ�%�k�����o��U$����꠸�F-	K{妿��s�xʼ^_��W�y��b���*V2AN��_=X��k�2V���H�RSD��pq�
،YT�*�j�)�����Cf��t�4�<F������QL�|�s��艹<��VT�c��%&30�s�� �-��X9�nل1�r&�(� 9.J�G��H��T8��?3yF��<%�4QFӸ�!�gn*�̙<�D��Φ�V>�j�C�Tg�'<F�0K� !�	"����׋�|O�'献�k�l��W$�\5�~�V��NU��]�ԡ�a/�9Y�)yq�+{H�#�$�j�C�ێ�����И�H��('{b:�a+HƇ�j�B�q��}v��9��)O>���ϟ����n�*T��a>/����F��zV�����w�������_r���w-�:T*�ړsd�=�$�-@K����m�PE�t�X��Q�Q��7dQ�U���Td�[ڔy��O`Ms���/�Ʒ~���D�4�Y��A(��=�>qUMĪ�iۑv;��+�1��[_���͚�E �T�Q��Z��H���M��{�͊>e"�쵒�]��UA[:�}��t���	t�!}��� 5]]�o~�XO�����ĺ2osz��^�a-�Q;Ue�����?�.��T5����;�@���`����u�C��s�y�6<7�����z�����mǒ��M��:�ғo�q�X1������q����*�C[�z9Rڒ����ʗ���#x�/9ʒ��
b\H�ң�G\񓩁A�k�[W�d�)RK��@�^��|�(��'|�h�pI]�$Z��e��'K&�ՙFV"�s�g�m.���b�I���%����~�!�[�F���+��$*�T)[�s�I%�''�5��d��`y�S���>;!;�LE�v�sf"N���i�����E,J[�Ej*�>7�\h����}o��}�?�3x_W̛�7��`N_cy���Ɓ����.
9�Pjo��)%b��=��6�HU�\�#�Z���s4$��<���R��(������Iє��M^.&���^���5]�
�k_�Ƴv{�ǟ�T��=��Zc5��}&�E,ȱQ�o<99���g��p������?�7��>e�ʫ��p��Ż������5�cR'8�4wH}�N��7��⻬����Ǉ��_p�լ��ꖪw�Ržj��Q�!iO�D���zӱ"��OQ�|�6|����n�'{ǵ4��[�a�׬BM"I;�c���kRm�Ȋ��"�c�z�=ҿ��?����;�ҷ�.{�Cj���T�qU0�����"�֬��;\<�@UG��ş��>E���/�*�o�&�v=w�@���4
0úMϸ��3�:P��J��סr8��g}��o!5�Mo��mD+˾�bqLq�Uu븵
\9Ƕ�y��{z^<��A+O��[�ʑ��5���
�boy���p�T���^J�A]��Ue#W�p�	�G����:��n�hv�RT8��d;��M�y�( � �Z0�c�+�s���}�=�{�e���Ԓ�kX�	r�]�"(Hn��ȭ?�-�^�K�K��V���d��KT*��o#��E��Ka�@��=��`]p��hBŦj̚�"`z�3Eh�hq�zb�S�G����M)"���cD����E�6�P�DW�D���5�)V�,JՊ���x�|���-gt��*:K�;�y�A{��~�����R���\�J`�<<�����P~7ۑ��G]�k�1?���4�!���u��n�j�$�pI[�����,�W�,��ꔔ2�v��{����Q3E,:�O��0z�L����E��\��
��+cn��Il�t�;{������Ǽ'F��RB4����8i���CV�^�M����ny��C�������8B�~cR��.�1j���O�Ѱf���op_�����d��>c����ɗsǦ�h�G���ԁ�3UH.(�yR��;�����ÿ睿�-�ߺGZop���@�&|��plr4s,��{a�S��=��G���ko!UźnJ����,���~�@s���HY���m�d��z,r�B��T�7�T�Q#Nr�h[�?f��;�D+��+�9�����6?��ٝ�B8�e�۔��u��������n0�J��T������W�x��'�V�F�C��/)�z%������BV$"c _.e�-���BJ�Xf&P�:�T�ȴ��+嚧s�E��Sd��}8�J��`1�D�.ʪ�i��8c�1���)S���1�Q��2�˔��K��j��?�%,L�p������f8�c���Q��)}/jc��L�y۰����!�:��"�WLLs������s����7�|�ӧ����E��}�L�!,�./�c�/f��@���P����[o��+�M#��Į7�b17ǈ�04��7���[~��kK��	��J_c���pn�C]���\UU��u�����r2tVp�q����P����* ��5o}�/����������7�驶W\��|�����/I}J�'־��C�Ф�\Ν�.�4�A����O��mՐo�e����B��(���˩)٫.s�Tb�P׏��'?�տ�4UEUU��O
q�|�N��3�)���w��j�����_�������c�w���Gy���1���	\_=���?㋿��V�e����dN�&��L]� 5�%�K ��t�9�Բ�d�R�e\���x��ǩb7�c���s�AsE	��wH�$��}�Mn�����2���
�I���\����q-��F,6JI81.�3��͑S&c
���\��)��'<)%s�r��	�3����(�"f��)�֚;��'��@���"�[ �jI� Q���ORD�R��хS��t1�4�2�#��	c4ӑM�)f��~���<S�~g��L7�%�,B�qΉ���r<��\�ho0�V'�&$e�]���{с[�t~�5���ʄ.�kzm����ɞ�Y��倞f-���E���r��e����ze���0YNk*u��k�ӖP��σPŻ�ogd^�&w��`c��:T�i�΂��$�`)~hM�{OUR�r��d|U��Vd���}�_�'�=���^��/���=O?��������O�G����G{�.ۮcS�5!��S���g�*ɔP.�$�����cf�ƛ|���MX_��Ɠ
��6�Q���4�L����VL��7	�4(7ǿ�a�Ӑ&��X&����׿�5V��ޠ��~���ﶰ�^����������o�Zo:�Sr؃��2|��_�*&mY��Y� ������qO1��?W�y�~>gK㾱ߪ�"K������W��wi�bY%vM�s�塏粌O���qPz�T��R�̧c^���qɤ*��8)��c�w�����������#��ߧ���s!\�9^��6����N5�pa���$�� U�s���=���"���P E�ܔG)א�������kK�~�^�"0ms�10�,XE/&�gƤ��|N��M����hg�˃=�v�@F�ia�i�IXЄN�Dp@��a�;G�j��$m%+U�4G��+i��������;�9�P�z
�47��ϵ]ߡ����l�V��L���%P�o`1�8o1F�h���
W��R��J���6���_%���|��u���j`����s��K��;�˛���,g�rx�t�^i����� Ql;Ү%�L��k|���{��.��#�2���.����b���	z��`�)s��4-i�v���D&����눩g{ݡ�5�x�.�����t�����Q|ױ}�9���8�%z;�����_6��us;g��;4�s��'�e�g��8�zz>�1���3�K���t.K�s�^���Va}AT;"�"9��njiQ��]?sSL�-O�L��ilȒ�sr�ϯ�A&�1��7O�CSq��M7i��r$�99������
U�v�j7Ӑ�;oSIs���`9ƙ�t���wKL�軣�L�C�	��X����8��s�!"G��t���L�\��X��&��x#M�a����i��e���ک�f�g�A8#z����2jpSЈ���%�!�:��޴��3^W���G���I��tL���4��l����W�Z���7��RV���z$$q����3�?�\�AHj��3��!�����o���ﲕ��yK[u��%�4q���_|����o��]�M�1���A���TU�ŝ�5$P�b�	m
M ��^��)�O�a��©��*8P̬����{L-��:��s�#��l\_?����x��=���[���z~��uLM�-���e�������	�����yYfz2v9���W�X�H��ʗ���T��qK���7/�l-1���ea ���M��(a� �B0Εh���4	�}��׬2	�������������w	��h/8?�؏�,ӕ��sm��gX���&v#�%�l��p.3t�E����K�SS�M�P���a=��$�E�s���p@��D��A�{?ʥS_p��5=`s&�2���BK��q��<���&���m��s�~� 0hf:"�rHm/�c��M�NUQ�ٷݑ�4��I��%��Hb�z,�--"�z��hC�+Z���6օl�Ź,}���n�'��SDS$�ۃ+)F4�s�,Ox�4Y�I�f��/�����ﲿ�#V�Ry�}��M���ez���_�����'{r�ǲgʾB�!�{�]$x���;rL�ۖ���%`��DM�R�XSo�̔A}X�%�Ź�g���|T2+C�kw�*�MmX㕣��?���ѕ��~���T,��9"_���#^N��ϵ�sz�T�'h���ίPU��7��ۇ#@gh�[`�/�_/CӖ��0Is�	�Dh�Mhj��&�iB2͚�����i1۟�s�7��4��o���>��Tܘ�=��R�8R4�>��P����%�HbpŬ85S��Lß���Hc:j#ibF�3�%�������r﹤<^����1�����~�9��6��H��6����,3���9����c��K�Y�~���{`��A�Τ]r�gL�\�!�e�W_78��S�����9���6Zy4���(�na��x8+�3^$���������j��jK)J���,#������������\Ea������������wp��졉��K����R�]J\���mw���sb,�8	�u���JV�v���.��r�}]�aA�2b�H���#d�KB��)O�_�ҤTKJ�$��S�Ū�2�{A;�!/�'�@D�K��5�e����H5ĝpr&���3Z��ɐ�S^��/��3O!��=5�ve¼���9f?���\�l?�ӯ9��P�Ճ�R�ʬZ�}�0��f�#��&�I8�����,���ǽ�����T��p���r����U��d݃z��>���g�y"�[JKԎ.����ՙ��ڴx,�b4"�����GJ��Py�l�-��{oV��*���81�+x@~s��C0CprFc1=&�Z* �66LjF�S�������㶿�j���|X�g��=8W��A�T.���{�Bg�b$������#��c^&<ZH?���TE��8	��)9	�]����zz����tґ����X�-rF4�|��$��JT����{��.�������{�*�$By�Uph�ӵ[R��Պ��1��E-����	<Y�˦«����n˭����a��mW펋�.�78���(����(>wt8*��^S]�qA�}nd�3�G�q��s*'���{�U$'������BNJ�9)u��.r�Wl��׎M��펰Z�Վ�&R]s�vH�qig���Q�kQ�Xi��	*h?}�'��B�fNϷj��hG��&ʎ�|�EϞ}�E����.+����!�S�>8��1��:u��S5[�ꖍV��6.�c﮸��Ⱦ�B�تgU�F=ɷ�%����ӅH����"����Hlwh� ��eZJ�Ԍ?%��+<[��x�}Ɠ���U69*��R𦏤&���kb��#�,7:��h�
�y����oY�۶#Q��gY�	������H%�`Z{�U��'��I����N^��t.<ng�X�d/Q�<b�Z.�[�w 骥WeJpWV��.�$���-+�I�=�z��8o��8'���)�	j���V�(�]�{Ż����nK����1Z�l����*��B38B�HI�. !��S��:[�3���( ��@!�處��`��
��9�"q���hs���:����`Dq�pfr��j���e˨��B���␴���<�or@��	3��5uO�ǋ��T���C%��-X0��!V@���n����/���v��c��/yN����f��cű�\,��y]��O�+_;�dO�]��>E��,���c>|��˧O��ʊ}�,?tx)%h���f��K��y�����	~4b4���M�uM/��IV%+�ǩǫ�/~�<rpoZ)���@" �k����|B��􏪒5��FM}�yYK��j���|EJ��#�i�u��z�R��
V2�Z@��'g�uC
J�$�ӽ�@?^�@P\��FH1ӥhQ�c��cR��bs�mY�j>y��[wo�}�{|�'�{vŝ�-4)1[�;)�C"�85�ISy��������Q5k������K�� �FLsW� �J���Vu��e�E����{lћ��C*�:-¢�5���j��v8�����uU�Ê��-[r�`�!Mo.@w�֘��ZvƸ��ċ,}Sz6�s����y���Y�xZ�:R�A6ԡ��f��@K�4������S~1�i�6̓�r�'ɂ��aO x<Y���f�⋒�H��z<��3�dh��7Z�}~ŝ�6�=����6>8�G�2�(�XϳƱ�`<����a�J|��[.*�+���j5�	��{�'�l~��7����D�(���h2Z��ȩ�9�s&��̵���U�Q�9�pL�:H��&��q@2;h	� ����l`2�����9<��Pc�yV��{nݹO������q��r�r�����|����$��
:��,-���R_U��q��'G�A�/��0�{c���*��(z�"�Nx���<y��^X�C�7��Ϲh8K>�cfd��٪�ŔQ��"&�ȫ5b�BJ��	ΏVDGK�ά(�G\�|�:O��WH��M��g��AUU�W��Rd���=W���?�c��ϐ��<�:�W﬉�~�����	����H�
�x�zE�C�D#t�*!	h�}��e!:e�d�?�]w�hy��67����Wa)^��u \�|���@� p��~�9��#���bG��do�nH�*�.)�xr��(D@$�N��!�(��0
����!K�^Rh���6<���$<y�}? ��!�ba=҅캉�`9D���K4~�v,���%�ąa`�3���R�K������kv�}�yw4����W������ѧ��;�]\2���o8'�ee�j*���ܮ��Ym����5U����)?b��f)H��U����AFJ(�U
�4�Ą�M�Ҹ@�c0���/�D��������vt�:<M    IDAT��0ѨA�R�J3�	-΍��C[�h1&̃�q�oIV�xv�^��ϟ�����Mɦ��]ד/�������6ͽW�D`�\���
K�7�!�}���ĲACh���ȮD[��}f��r��AUm����, *�2�� �,,�l��YW5�>����#*�33��J��1��S�"�(���:��NP1���~M� ��Vo���g )������b�(Q�`�=J��i>k�w	6��Is�>݃'T^��3��
RF��D���$Y��ə��!?�_�g������_c�ګ�������1���ͳ?����^�����0j(��ݖ�
D�))��>s�\�ڌ�64��q���>�я�O��
�8��k@h���!I"I�����PQՍ	�<Z�oLi+�pm�-��$�3����6e�@��~��8�xGw}�:8�XΝ	�������tH��h�W��x��s������;UqR�jë�����U�1�j�Ӷ;C\G��(�V:N)�<l@U��U\�C˓��WCP<�E�,l��|r��!����X�T��Wk..o���_�^H[��-1����DK�����1�1{P����	.g�F��E$W�>��������ּ�^���vk?ƣ)Ƴpr���|{����^��`,��L�� M�DҚJt-sx�M��8���9Xr�6��5Hi9���|�i�ĐQ`Ea���/S�<0>t�a�gU2ٲ��#�j�;���,ȗ5�/]7��#�rl���l���s���.�qօن���/��_�>^p�x��T�i�5�xuE��6�^�ZѦ=�3#I�|�̧� ��V�(j~.��`����d��qD���9���1�aG� -@ҿ:��T�W$G��s��!�1Q_��կ}����A�+|�x���!j���Q���|Ԧ��#��ׄ}�V�7��O���=�3��TUE������ffw�0�T#��_����C6�\��X5�������ן�ʭ;��{�]$;O��T
}�ȕT�}M@�z�7+>x��W��
�_�������{���1��.�	t��p8xAK݂%=���,�c�=��	Xb��K� �5ѧ�TUI�@{� O��-.�ޣ�ܢM����$ M@�!�iZ��Y%�5�L�����a��6;�=sE�&�~�M�9�*��q�|4�+\\d��L��[A���ӱO��qN�=5�3Ӏ���&���y�E,���DJ��!���W57A.��CC�q��s�����g��g����6kT� �R�*�w�Fq}XC��+2#�U�����[�^�Zw�	���ϟ���E��	�0�С|{v�u\EO���1@pF2��j�%J&����S���A�M7��f| u�r��LPǦ���5B�,EC�C�~7? ��|��&�A�9g���R�Y:��K��>=����h����Ao��u҄
4��w�3��;|����'�7��G'}I�4XRh^P[C�n����F/R@fp���U#����9��
}�.�/�I�/�~��U�Tb�{����\I9Pd�I��'��xp�B�	�y�D��� %����0�̃ˠ� �c�G��9�����kw��}��<�}���>e$%�U ������UhU�^��'}���R��_z���/s�wiDhV+4yR$����d����<T��יn���3r墳�t\��\\��]���Z|pd�Fꪁ��^�W;�w���gx"���t>p<ן~@��hL��Q�yn*�.E�XƳd���d��:��*��$�Q�-3����9#|�O��4��}�����2Y蔎~�ȟ��������b��"/e#��^�
j��K4�e�lßK���=F��T�?�i�.�!�b���Qt�k��g��S }=?��<
Z3���X���,-4mw�P���b9K�}ܲ�wH��lV���$��xWXY������Į�,W�m�651G��s��zRn�b�Za��Q��!��ދ`��S��8���td�zB����/L~z͒V���n2S/],������e}��ִl-�
��O���a��d9k�d��9B��62��:���g�g������j�፯}�6�.�<z����^�|�fz-�˖
e��m��8�}���CD�W~�k���׉��%�	V�������'䂌���O�G�Р���<�*�T�'d�Z���da�����k>���>@|����P�LG���5��yU��2��q��������9UThV��o�֗D�H"�P
��/� &�X1�I�O��k֫�\'���6���gU;���츾�Y0��O=��:@���Z�+��p��l�Q�����UR�D	�q�{�P���
~��c����T�2sgR%b�[��b��oے�bܚ��k7�B��YuV�X-ۮ'�[���!��G�tI��7ͭ�Kgd�|@k;(@:2
!q��+tv^���~<7��kD�*�Mx&�;�>)5�-�b(*5o��<�<�?�K4�E��8�x֡*�$o��(�Ij��cN��ں��CE��^U�u �$�/���kѱ�z��U�\S�*�uv��ytM�d�Ư��/��t~\�t
 g���R|t]in�yMs<5�G�NM�c��4��C���Rg�5Gܛ>c��,�������M��#��ك]�9���ڋƼx�p���WOS�8x��Ѫ�O		���$8-�y���q���O�e�����Q�������o����7�ФT8����o�uR�;�ŏ)4� �/��gR�r�]Lt)�EX�)a���	q3 ?v����ȳ�>!^=1wAU�>X|UQW)EL=rG/#�%��=����C��G�E��Ľ/��嫯���z�eߵ��̫����'��~e��D{�N�]���œrO��S��~��Kͭ�%V��Kf�^[Id�H��o��������|�w�C�Zq��<�����^�Nh���e�)�IbA��A�Z��8a��9�����\𖡠�T>�Рs�o�%�Dլ�u���#>������s�H����Y���+b�ߍ������.�)m<�z��$�,�9�@��i~M.{�Ua,#cg��7T�^*�������ئ�/��<k�L���x�r��u���g�Zz�E��Ex0��v� ^΂��t�If@�5�O5�l��Z�WHv�{;��&�?�NL�.Ym�ܠpM�>~�>r�%�b�=� ���!�$)��oQ+څ3�9��>+*_C_o
Ꜩ�V�J��
�OhT#�j��":���P���L�BB6�ɸ�w=�l�}P|vT��r�Z�L�۔XgG�+�ޡ�W���-����~	�����%Bu$D	\����o���,R AR��5�҇庒�~}Q�=�?���X�RG�J��&@�l�5&3��CD����� �L���5Z�i�P���Zko�K}�T�Y���;\G���?�:%��oj�EX��&�ڎ�w�Α���\%$�C�����#Ǟ��^3MӰ�n����D�.y�W�&��5�k�I�H�=�+D* �z�fֻ�*��.�\Wt�w�u�xR��=�y&���U�'{vx�������2�����,�>����W��<��U#��9�����_�����a�.�����
�ЧD�B�#]�*=�Hū�ˆk���i�h{��hE�ޣ��Np�.� ��<EG-��H�g�6�$�#��m❯�����7���x�?�3����ZwAV���O-=~A�@ސ�=�ۓCǣnŽ����_�u>�s�����C����c�6�����=��
�I��O�J���;v�ҭ6�*s�:�O��~�C�;-W��ʯQ��iG̲x�hh����%�(}��Q~��1�o#���'�Zc��q���p=Ƣ,�9s�B#�/�l��1�܋�*�
%%�X�Zisg�"��r�adFK��ar$=XJs]P�N6=�'��9��m��Мs�%�Hto���z@�qNY�}E﷤�� ����'\����d{0�`�!�UL�ԳA�q�8��R��"�YLHN��
��<	�Lƕ��s|�u�ۖ�4�D�z��t�؁�I��7����-�����|gC����3?��>@�ؓ�	��6��1�7�tc�wF�6ka�m���Z���aS���o~�M�z,�5�R~9�X����,<�Gv)�KV�q�z�}KK�p�n�����M�/Y$�������|��MS�R"��*��'�6MU4�i�|M�,�������P���<f����g�o���֪�س�z��9MmY�ǌ�Ү4�*x�������*_~�m�Wy��Yf����"8�זZ*2��[�ܾK��k<M=�S¦Ƌ�����l�9<��泋iON{������'��?�Cx��~U��o���x<���i����\	�g�cs��l��Y�D_;��q}Es�z�_�o}��zܓ��|L}M�Dl;\+����d+X�DE������/����=��O~J��)uj�ԡ��Ǽ��9<�����d1u]�$�.Eb�E^%�Bz��N�I�+4�K���TT��d,�d�`�i���w8h����M��6��9��YKG��p2��&H�mF_��G��CߦBҔ�h�=q1��r��U �L�w��I7���Ƴ��c?�&�r��g=9���� ��ob��/��)����<��]���~)O���4�ab�~�'�KI�p�QJԧL��L[�������e�T�(j�<@��ggi����py������ ����|�K~��"���y��T���U>����3�UM�+nݺͼ ����c���L`>��χ�M�Z�����|��g�\NTάZ _�q��hm��p熠�L �>��~�q�o�U��X��v�����Ԥ8��%8����d���1�?y��xǭ׾���o��;��h��}˥ `u��h�#kO�\�;\����q�B�ʭw��W���K|���ʪa��+1SB:7]��["������#���w�����_�y�u|~̣�����Zi*T��`��-���*W[a�U�r���Dý/��S'TW����Az���B��J;�� �s���Ugs������WH��YY���� �d� H�y��J�LL!k�6ׄ;��\�Gh�)�q�Q;���r����2�y����v�wA|���M�-�lu�䚥{Y?��]����������	�$A�۸�4}On�%�Cȉ��'��9���93Ec
�;�i\Kg�t�
Sw 2���������H�A@ 7��qB�&�֦Lf�q�Es�8q)��Db4�����fS�@F�RJ8�R
o����ʱ�9N��M-
�z�!0G�ZZ��{�q7�*R���"����^���B�b�{N}���{����t펐O|�Ï?4�puC�Z j~�A�6���7��5�˹�>'���	Iw�b�ۢ�*�ۗr��G�.3N�������i�'��sڇO�l.���6�2;��w�!�Г���׃����|�'�g|�6+���_���:*�
�hƹpt?u��H���������Ct�������?��g[�X��o�._���.\���6�.�X�N�L�p>t��@t�ٱ{����@�p�wy�o�����&��>�������!!+�Ԃ&jY�}��>�յ}G�H�kv��.qs�_7���\6"��ǚs>c18�����	��R̈a|Ľ�C<�����}k
�,�i�b)��V\���o� ����{�ݎ��9���m��ڋ �8�ʆ��x��(�S�4
r"d�L�2��~/�ї�O�Xrڪ����3�r]�x�D���!��%\��Ǐ���b�Ss��5��9=2�����l?Lg�鈎�4�C;0�c~�~���_�}�tN-�~ДG�����sL؇N���;�'�5Gւ	c�;P�j� ��A����P�"9nK�4c�=�W�"��@%&I�y�˼�λt�@y�L�����ub6<~�9z������{_[)ݾ��D�k��tY�F~~oU%�LNʀŞ���,�>߀`+���aÏB!�9��HrЊ�[o��%1g<B�E�^C�9,dӖ3�"�*G ��?��_|�������9� �؏ź�k�4O&{4f�>�*G�Z���Gtۇ��%����5���T\i>�W��jV�5�jE]5�}�Ʊ�o���K����7�����C��;��Ϣ��y����'G"�'1�{�����Z
�[w�?��~�;���k^��[����O�>�U��#�<�7Y} �:��`��~�V6�y��֌Ӗt�����7j�jn3F���,�Xa2 t	�jE������ݖ[�`q����P[�/����eO�%���ݯ|���|��پ��Wb�!&\���x��QI�=g����~.���jY(�P��|Z��f�㆛�O!����~�6�O���p���5��司��3�i�F?��0̳ϚTs�A�d�΍��S%p��vt�F>�k�(�t��HǱU�U�!g`������b�g�|�	:"\��rn4����5��ξ��% �O���u�j�2�=�?�z����68�p
"1gt}lqU Q�ݎz�fǱz�>�� g!-ޣ/��6��M17	/����>�﫦���.W���2�s�9���Yn2�O��&��jnȨO$pa���������<�6o}��������zb~��C��V���mA��9QE��I��N�G]��>�r��(�G��~���mۢ^�\�\t�U���S��m^��/�6���;�8�Pr^g9M�Ѯ3��n�������Bp���<���v���;��?������)�:���y�KZ��Ͼ �m_+���c���7~�/�������㚧������{�1��v�Ka�����͵�.�(=��}/��o�����y���'�}�z�s�k[�(�����v�n$�ȯ�=>A���Ɨ�ү�M���h��WO�R? ���V���\�^��.�\e��W���o��k>�����Xoj+BT�!�	���D��t��rdݜ�с]��TS��Q���d .��ꛄ��>/��-���!ܰ������{���O��?�駟�i@ԡ�,��s��ߓ�EJ�[q�O����ð��#�	�PAϠ4�4�s���X{�fI����w�̬���4 ��6Vn �EC���LI�-�'B�_���3̄�Bc�c"<�4�(�(�$n"���h��ܾ[U�r�8�YYYY����ڲ2O��ٟ���s��\�i!em�n�6�%k&�	<�R�rPT�<�H�J�|_��������Q�����_�~���;���cu�s���,�Wl�(%(�)�P�����Z���[H����q7	�?��[\��y��g�N�ɋ�
A��+���a����nֈn����!F�:�Åȼ�����E��������S癆�W��W>:�A�zTL5�A�J8�`9�bFF�g?���r�A+�N��s k_m$2A�����AU����vnc���~q�,����e��g�M���4JǸ� ���o�V�ݟ���?an|BY�L�z�/��M��}���]5�֒�"��;}�omW��q�i^�����}
��c.��ſ����&c)�F!�(M�!�5��h�ٻ�W��(H�!�}��l<�f�0��}.���H�LTR3ɚ�w�լvg1VR:Cr�Y�<�z�QŌ�+�����	�Aym�VG�-Arɉ�Ԡܜ�ﾆ��%It�
����c�B9���u�uL�+����Z)�$|eqe����Z��~�^�h�R ��g}j�7)|1$ַ�H/ڤ#	EAug_� D��5>�ƽ��F(�������c�FX��j�}����K#�/��Pk�p]**�u�=��MU����dF�J�ެ�j�.�6J�Z�(�ֿ+���J)<��*�E����Z�{�?�b2�B/Mp��j�5}�:��9�I��bz���;��J�$JG)�uJ���M��Y���&vq�Z�`Õ�    IDAT@2�LZ�a�g�}�y�ls������kw�����I�>�k�;j-5�)��yy�2���7�:er���9]���8�}S�{-����
�-؂�?`��mB�����:�����i|�r���Q��=�JIt�1�8����^���%'�~����iF�BT���8_PUs�L��m��%�c����w���?y�� f�����SO��|p=�<Cs�nn��ٔ3����� �dLu�}~���Ov~���L+�2����lJ�%,�)�ir��Qy��:F�������|�m�YŶ�jD9OaBX�z�{�d�P�@������,���Mv�]��s�R�֪��Z���X�_S�>���Fd)NBb�p�T��*1J��!2�Z����������<$���j��T�r�$�*�Q˕��ߋv� ~=s�WEH�~�c�}Ai
o�ޓOV�9��u��7}�q��J�R���u�a5�X�nU8��b�:�G���F�RJ�JP��-Q��e}ԋ���;_Ea2��bU��"@�ã2M)J�j�LE��	FEk+,R�-�oI�D�ZEbe��}��m��uu���t��m�<ʃt�+bQ'YD�'�)2Pلl$1�!�F��u.����M�ed6IU����&�9�1�#X�w��#XK�Əc���D�K=)M d��)���H�	�n�Zε0cE��c�g�(F�&$�"qX�p�0�<�����.������`�z "eB,s*��EK���F���p�kq�$�F�n*�5�흊0���� N;f̑#A��o�g0*E�ĉF@�,N��č�)b����@��vR<7�I�l�1���0�u�<q?�}�-+�*����@$����mM�Ԅ<�#���B	(5��ܘ�\����Gd���^�:�'�Z��i����8U�]�,q��R'*ly����4��!������{I9Ҥ�\��ϻ�������k���䗮P�Y�D�"�B��r5"a���pY��*b�{J	��!�.�{�f��=w��?0��+X���4�s��I�鄢�Pׂh������g���g%����rx�,g��,�l���0�rl:Co*��)F@ad�|�v��I,�%�Ra�B�1�,�$da�4p�_2��˨���U��U�U�2̣�,ηM��9���l	�b��0uY2b�T{�T�&G ��S�1Z��-�L�� j��uLU����*3�Ay�I#`7�saۧ���s��)Ey���D%�2�]� u�ͺ�J�\ˤ����)D���>�w/BE�D��S8��pZ3�6H�&y�蠑>�!��R)��xvu�5 k� !��� ��!�AFDH���*�'��@�E dߒ�ڽ"H���(�̨�2�0B��$�� T����E,D]�k@��x�s�q���S�f�FS��	h���6��d]_��	�X�Kf��J��������oYYdbVҿ�` G��e��Q��N_�m�G��`:�!����e^��	���Q�lE�k_t����Ǯ�0tָb���`�̴2�����=O���O�p�DiL")3C�(D��,p�р]Y!T2x������v����he�_�A�JP�<�7w�Z�T%�s�%����	��}�}��6��WZf������'W��

/9���4:8��[��2��Q����jF�V%R�i.����������S_���#߻���f9FT����{���$!D��t8B ͣ��	]����gs&�3Έ���)A|�5�n���66E�����7����/�"�����:�g���1����5C�xDP5�YmMp6��[��ן�o}��܍O���/�Zrn����121��m¼�z�͎���'��
��A���tc��=�@}���ɄYp^Q�=ގ�唲�Q�C˶� [���E�4��՘�<ʉ��a��]��=�!e�5ro���\��ۼ�z��:�~i�E����:��:ȭI�t��ꃥ������wRJ\��@ �k!JEs�V?��h���������D��V
�d�����%k����"kh�2��9�? Cl.=d�ۢ��n��⺂�-�Y��JK�j��Z��yԍ��k&�����LK���Z�c��-�>zk����
_%�c��Dw�����kS
�� Z�s4כ͇�h������*JTYpp�r��9٦���Zm]�X�T��G��Qf��D�jl����#�T�Q�*�lʠ�'����|���g�E�a�#�]&���ИmewgQTTA�y���E�D��1�	p�.�/]|dJJ)���Bx�������՟�)jr?'^�:a�׋9c��B�Ob���
ӫ+ߝ��ϥ��"�$۾��|������Ԩ�u�ch/u�rfl��T���>��w�v�%V���C�i�:�QTH,BƠ��*G���=Ʊ�����U���7������:�A��<��r%���>����Bh6�>͹/}�
�μ���Co��{���x�ŮQ%cF�fb�l�%Bt���ªן��ա�|�6t�\��O<�����wns�ױ����S�����.�o�;4�G�k�X�mB�$�Z����ֶ�����(%�ֵ�4V�~�kI�y��%V�n~���>��q]�"������5�(Գ��ʄC4@v3�h�,���z7�.ш�4���EbJ�#�Ng��A�bw�@�k��\g���'�ߧ���"�#QF�|��%I��檘�f���Xh��
���¥��8�]��hj_�����P��%| !�*�_y�>��w6Z#�1>D�T���<޹�t�W�eh����mCX37��ֵ�P/w��.��SlqȜ�ѹ�8��yG	�Dw�uNjo\�)w�u.�0���Gos���x���<�ŗ(��2��I���>G#-�L�昮(?x�)3ax��������mL1݌�|>�V� �JǬ*	ac!���ڒ���B�Q�2��F�^r���I_��5s��U�RUX�g�\9�]�D#�ܲ���u)c�\/9H�(1̽���/rߋ��4�M7���ט^���B�W��0�	1`�>$!"!ʔ�O|�cϜG��n�n݊.��ؒ@X��w���2�����29u�9���޺��CM����G����Qܺc�A����ݼ������i
��SЧw���ں�����:�7~"H�o�$�)�.�T��&�v�9vt�P��!�ꀸ �@�Ȥ���}~! q]��ǁ�+!���}[�O_���ˮ����f����ҹ!k�N5~��_��x�#���iJ�y����y�"Sݖ5��g@R�N|嫘�m25�Ō4x��T�cn*��%�F_��>�n�"=)�Epc+}�G����}��јE�C@'
�w>����!I4�+�S�u���%;���֭�#��!�͘7��{-�ad"��a����ipxeH����1�|��4����owLʋ`�-�3������ޯI�'5Ǐ��DG���l�N��1?=Ib-��mnq����0'�5������䈇��M�#O2�:��N��1�&#0
'$��0�F�ٞ+F9l�	��(�
�(+�XO��klHp�� ����ȲB:Ɇ<Ɩ>��e-���Z�W�G��-@u�4B�ʔ[6�{��O<�Xyn�����ۧOGK@X\��X�d-\+��ף Q�Bu���{7���s��7���l�u̦?F��z{¼(9LF|������=N~�2�}���;��:־rV���1���?����V=��jUU��$Z!L��{��:&߯���.�ِ �d)��v|��JE��j�Q�|���f���o�9���C�":j<�L9~�ľ��$I�Ib`hON_���QLe�C�21]��!��k(iV��M ԝ��ؽs	��h��h4��ߝ��>��u7��j=Si��a���ٳ�<w�Ys鱱��QSn�|DL���e4��_����@k��KV.�|H���x�'T�`ZQ9��M�Y)�	A��CsޞS'nIa[�O{4�55cb��F�ׯp��/�v�Id�d|��R�X�}X];�y.�a9��{�x� ��k�1Ĺ����ؗu��n�\���yQ M��&u��sk�B*���	7~�3&�.�[6{�s_�=���`d�$MЩ$d*Vg�-�����NJ�D�dAc�����§����6�u߲���,D`(mb���KU"��к�L���Gj�L��p�Ԅ�� y�	
;c��K?�;�+�Ʌ���>�H�ø�H\�_U��*��!�x��g�2S��7_��P����AS�A��R�M��ǣ�ۏ>�i����?D9X;c�-8Y�pM8r�U�ٺ�ۖ�o��� �6��GD�~=y�Z�h�CM�:0�֛��h6*
�!���(.�Z�=9�CB�����������-Ʊy� �o�w�9��4M#���5vͰ��e���i��vd�D��K�	}������C��P�ʡl@�U�\K�E�4�C}Z�ai|����Z�R��V�F)���{!8������?�MRD�����ۜ�r�Կ�u�`����j���.*џ��7��:H��C�@U�TJm���'�i�}:�cլ���c10~w[C����������.x�pl�S�k7��2��!�P����0?`�-�ܣk���xf�2�,�������Y���'8�T['�u0N�ye�k��XFU�	&KJ��@q�d�`l���1�_�>���
�~�l��[���l���9�,w�c�Z�Ts��L3O���U��(Cld8�r5?�%�Mc��Qw���T'щ�4��$�L��^�a���΅�Hm>�l|%$ӓ��ķ�[x�sd圛��1�o��S�b8.g���Ѫ��m��*=��/~���}���Q\��h���?'H�r#z�q�J
�#�1�a:�oڴ߾��mC���?M�����C e,�H�����3�~���C4xM�^{��u���uiQ3���W���x�&������!�g���t���s���bY�S�|���
�����}���E=�{i}�a1 ��hC�>�&!B�*���$HRc��n��,[�1v	��d3�؇��Oj�fB`:�����;;��ὧ���[�)rlmm��F���3��ώ���X�kZ���1�7X��t�ݢ�4���#e�J�����T�et�꽬�.�<0`�Z�F:7�;�!��wP�	ac��?ǹ�z�b-:��1�r�Ս��� ��mQ^���/���g���SOs�N�i��*Te�$�� ��r��*�:I�b�!�ۛ�勼�w���k0/�N?�3��&�gqZ������I�1Sɶ�TCT��i CbrGR	DU�ʂ����>bں�����UxB9é9!-�XL	�Rk�V{�Z���K�� b����g<���a��W����������Q����8��e�*���s���0�68��9�q�����]�@�u�����J�DEYM��%,����Pz�1G	۟���#F`�
����1���{0^�/Cty]?���K�T��O2�D�=5m���Z*[��r�1�n��w+Zz� �Q8b����:N,c��e�t��V�mqf��Wߥ�}�n�j�"u�}�du���`��m�h��}8�k�Z��#CL7S5��d�!�)N	lph���^ͱ\PhB�CG-埋5�j���:��{O��`y�&`�	{���R��E؜���+����������|��WX���<���O�S�%H�� (:���7�!@P�ܻ�I! �%�!e�)���l����Þz�2/�2�TT�t�*�idI�`h�N��D�k�T���:�)XWC���K�B�uUk]l����D����]�vq������l����ܿ�JS��L|� )�`]I)�x�
)TG��A,,����S?%57��6F(R�=�4�3Rlh�(c4� �$��<%3%�9.ߧ:�%�hW��gqe���I�4�lm�P�_����o���T�8�����d�s�l��W��p&��,G�RD��(-�8p%�5/p�C�[�&�z��Ǘ��F���jP���)8]�A�>q�RX�
X��A�*�p�P-�s�h��2� c����}o0^�a=2��.K����/�>b�`����9�ׯ2+��2�y,VTy�T�c�ؙ��Q��
4c��XH�-=|�o8��s��|��ox4������h/A�t;�A�0�B�zM��H�`��g��ǎ������աŸa�1Ŋ��jه<$����ܫ6��k� x�(����P�8���&�x���&�$Gp�P8y�y�q���f²u5�U�v>�����{���m�`%d�O� h-�dX@i�'	�L�L@�=�<�L>�؜P1C���b��R4>�D"}�w_���-F�ŴZ�[��%RTH��b��"�J_ã��+\z�J�Dh�4qO�Z��%��H��FF�WB,�eE��9o!�APZ�ts|b���� c����5m�	��[��i��v�B��U�W�����nnQ���^��G?�{���ѦqO�$�ٖ"@>/�ۻC��̕��$F�\D�`�WQ��cڗ���C�ꫦ�e��O�2�v$����ػy����N�G�R|L���AjEс�m��O��GW�鷾�b�����߸͛?�)��)�C;��cfJ�pH �Ht�:Ru|�+������Ûש._���>�(O��e�*Ì��ST@��j�*��j��E?��(i��dQ@0��Z�t�������}{�2��&�}�T>�ua��M��1V��DL�z�{u�����
��b� ?	�%߭u���]5[.�����d�:���"��Da�do?��{�s/�.ũ�I������x�T(6'�0h\Y��_��s��iM�N#xZ[r�6�?M1�PɊ��磋o3>���ٴ�V�7d��?g�JI��:}_���g��6W.����G��I��ߣL�G=����.�i���D���Rd�)�q��c��ӘrF��G��S�-�¡䪵rh�������V��V�
��(�����<���8��9��;{�����U! �����+������[W���?,|��R�~k���:��Ki�g՗Бhd���y������;f�OCSUCк����վ�ja���.I�=���,�ܕ�x���h�1`c�0�
qX��� ��8W E�a>i+��E�R�� # zeȠ����M�l�D Ձ[�����ER��Z�,w��c3"�����@���̾o���}R�L��s�yZ�*��{��L��bs�����)G�Nz�X2��8_2�Z�>�*����`9��c.��)vac���}	9y���R�
�Ā%�h3Ai�v�5�fr�ƒ��W�H&����s�kQa�x�1>��?C>��wgdڰa2�k���~ ���6֏q�i�cnY�`i�7���r�߇̂C���k2�bns�PrX����2>�<O����c��G̒�\��?�r]y��*�/軛���E���t�����(fE�?�_����� g�L?~���%��`Q�}�34�!K�E@TJ�l���O�*��+̯Ȇ�UF�i�ӽ0�n�V���+����ғ{˾+�㔓_�<�S۔W?��/Av��Z��:����}�?=�Ueb���[���A�����m8��L�����p��@��bj�|*�[�s�g��}��(�z�~!Ze��6������V����S(�6n��74���<�F�Z&��İ���� �F�Ie�^�+Q7APem��6��*x���4`*Z����\>�:�e��'�x�� G)C0
�.�L��=�̽��o@=�C����H���t6�� )��D�t{�
�z|2��ڤH
O[1���C�5}��?4�G���'t���bk�rJ	�b�2����<�;@n.�ҭB����{���=�1�S�s$�dÕ���I�=n�9������^b� U�ʗ�4�*
�l�b��~v�a�D	�R̦H%�J��G\��������ȗ�Σ��o�����AIK}U�    IDAT���TSUC�6Bd�1�VՂ���
����?]�ߝ���)-S�� V�O_�Yg�Y���Z"�~�P�)��ٌ���y���������[|��̵_�L&ʘ^Ti��~�^�>FK�mB᪂Dk�6TƐ�=Ov���|�7����3RLt+v�6aY�ij�Ct���u�d��p'�p��Y9%�%
A2H��Y���wi�%.�ڏ<O	�)]��m��=�������6�ˈ+���}���}m�z��w{�������J��3l2f��}�Np�ݷ��˟QJ`%1'���c�?���EkW,�;��F:,[S��������Ww�V斈�E� �n�bOՒ5`��'�C��Q&�%&$:�L-G�]�5���|s�ƍ��k���ۚ����3�5�uz뚖��N�U�jM[9�k��������3�1;�9�*�P�{���g���& gi�:|��Et�څxR�B�] ���%�z��B��D8��?�ݾM��y�_~�����;�$���!�b�(J�"2���b�����l���
�{�����~�C�x���>O�}�	��Nbk]�D��4�y@�$�`���z���_�ٔt��}�Kd�=@1��y|�ƣD`[�:�E.��=�U4��CT3*��ȹ����O{�(��������`��qn�i~8���e�B(���!h�W�w�~-�K�sw�e'�pu^��ݫ0�c@� >{d�1�<��z���߳��/����E���r��G�d�ǔxL��>V���
J[���r��:a���/}=�z�w�n����a6]��F[b�+
I3��g_��#<�������s㢏6�wwޭ2��o�k�s�3���T��Df�̘Q��XN�%p0e� '@ؿ����KE���#�y�o�~�uTg���F�z&�<;RP��1

�	�d4��$���'��%s�)k���}�h˥f�����/�2허��g��e!�%(�����|�޷Qj!?��G�`��{�浟>��}B������ ��'I���VW�Z'��Z�]���*���Rz,�"gS�?z�G�{�o���������#��bV2����ݼn���Ll��c��ƆK/J	F*���2Qq�7���{Xk9��3l>��� D���������F���n4�����_!5i���n��/_F\���,y�q�g�d���t��>��{ѱH�J�[gK��+r7�����l?�4���7��LmșMw��y���L�yw�0H�P�E"�FAPy��ƈ��x�Ʌ����/��>ˉ�����;��N�k�m�1�������)	^BPD�`�)Lgl���IJ�kaq�
���%$��p͜䁯~����O�:�dv��W�{���M�~���-����_E\�N�D[��'t�$K�u%̊,�T��A=���6:����K��̶��} ���Z���V�'I�<�O}��_z���o�΍7�"�����
=�4L~�����t[�k$�V�J0s��JAB�T�1ز�9:�n}���{�_�9�1+E�p_����#c��B	I���~K�b/8������ۿ�/V��XT��}��A��ի�P�P��hj<  x�
��6�,-����m�xibsij�u�?)�A�Y?he��D�J�RK��L�2�$M[D�~�m�!��^6�
*FC����a����W��W9{�a��y����L�$�b��0
]kd}M�}�R[�_���bX���%:��)�'����KLo\EK�F�H�fd2���ɹ���,3�~���p���{��<�%F(DpL65���w�g���O�����<ơ+�d�u����z��H�]�H34�)H'���~ÝW~�{�Y��/~���8L�!�b�I�)���4��s%�_^*�WTsG�-��|�����?��v9>ɳ�ξ���l-IB�CxDW�� 25G���D}�P@�:⺘�|3,��e(C�!�J��q�����w������5f?�>���?Q�y�LW����#28,�X�^�=�1):1�Reb-��Az�3<���!1��m.��{\���Y���üd��!��5߇�D"nC��1g�cc�r�����[o�U�H��xi4D>�[w~�)6��{})%��d&���z|���4��'Q�#�5"�S�+�\e�_���Z������\���ڸ���'	b����RB��9���<���/}�{eu�7
�Z��%~)Œ�ѿ�P�`��(�����~�e�e��3k���+�����_���ύ��B��7χ�jzQ��jR?��;X넖��G���,e�f([����s�R�J��ױ|�~�.�h5��u���v�W�Ǻ��0m-���Β�9�CY!��H%lLRaHQ�*�l,j#d]ӹ7�]-��ߡ�C�~H+�?[M��b�xd�}>|�g\��I�~�s���)��'�HRm�� }�f�cRH��t1�\MО����~���u*�0g���^�m���Ul	Arg ��l �z�
�(�c�Glʌ�r�D��8A�������z���1&����^ ��b|d����4-)Bx���8V�cW3����4s��v]ʅ��n�(!"�@y'�>�g��?E�����Mn��*���_�����l3Õ�����y5<��\w��yIU�Q��i2y�<�¿`ی��_����9�>,�6ی0�i�"D,1��&0�g-
P���ڂ�U��o^aTY�G��p6v?M����3���;�#Ӧ����lt������SOn����V��I�R�R�+kk�?J���|ͯ��R�2�1eR�#�������"}L�N-�u7h�������"ĂO������=cFR��f��ī� 2���r���s���h�*!�D]eQA�h������t�;��t�N��&���@�^�+�JP���b��h��@h�f,��j-��8 .ԩ�%�H���H�b�:֌M����T��IB�M&��f?�E�=��Уm���;�(�LB���6�7��hU��t%bs!�m�v�A���_�N�Eᜣ,s�P(*���Ʉ|Z���=��/sd����C���"`�g�rB¢��$�#"C߷R��j���:���TY�M��P�I�䁛���*\G�Mr�qmU����p
��� �G�@"%Z���M@��C|�XXR�(����C��>�?�s�W?!x�s����8�3��ݨ(���j����TJ����ڜ橰��ȠI-T�)9HIr��s�q�ɥ�������>���yq�B#u��uߺɛĴ::���y�R"�CHK������J�ҁ"xE��.�B�e�T��]�Y�rѫk�Y,��~m)%F)R	���o��H]c�տ���/~�d#��fL���ɂ���(*_�{�m
f����k��eC�������G?O��qB6e��W���:s��o�sLl`6j��B;&Rj��Q�(A�#���f�D���=�8�[��G���3����`��-aAh��56�B�b���a�� ��E��U#��%x����_�V�)f$ڐU��θ4��=� ���a'#��p��O(�&�	��"�$��m���u���׷��$.�g�2E�|s�=��y\w	hc�����)v��7��z¸4LJ�\͙�Qe��>�4��"4���ԡ���`آs��Z��x�Z(t\@8Oa�/�* \�w"xJWR�X��y�@G��H]kAj��(�X �񷄈7��uI4�!@�qߺ��.��	(,a��P��w|X����B;��J6����C(j�Bgb#3�%Ҙ����CS绵&���5�G�}���Y06<U>g�c����ǏQ\����K�V3��7Z۽�y���f����<�J�>n-��_�5���y���g_z	^�����aT��9<`4�%���Z�Qs���u2Yu�S��Q12
� M��r����i�Z��o�!��6���3�7�4eVd5�uSl���| 1��5Bj򼠨r��9�����q���m�x䛿ǛW�az���N��I� 8\�p5$�ЦN�0m)����]��$�³������]t6B޾ƉNDw�֭�n;ʚ�tN�A-�w��[ۆ�x����W.q�?�g�?�%;����
�-ib��K^�:a��B�(�s�9���5����T�>��o2߿�81T�$/k���>O���V)�+��F���u��>��3��j��_}���PB�CI:Qv�����{}���[�k�w3(CmQ -Z'TeAi����l1>y?�gNSPp��9�t�1�$ep���9�2ѵ�.����~qN�o�|�_�O/�L�� �砰����?���J��=2��@L���#�v�TA�
!!�\�Bͬ# ��\t�%Bk�i��r��=◪�����U�!v���ٓ�{.�˲e���5��;��pr� �!h����ӗ2[ԡZ���Bn�� b�
вK�	t�+�ןWM+fʥ�;�M0t-W��M�s!#:����������������F2�r��LX�R����M2���Ee��%����Tv>����E���O�羧���c3�	Af���������u�gVΑ�b�������q�����~�}g��/���i�b3���ǚ�5�d���$ea��DA�+��1���+�����=�͔�_������~�#�C	���#@F댳�y�CcR�s�XT�٪�l||��ۘ��d���4XS],g��-,�w�����w!��۪�8�O��_��n��{�{O�w9��Ϲ�Wߥz�uF�)F\Y�0�~�q�?�E���</I�B��r|��/~�G����z�vz���Ӌo��9�Xk�mA�*l5_;-�ESV!@U���܎�'��BS$�\���o�D�XXʢ������>}��C�7L~�r�4�#�T3�X$U.P*Qw�\���adZC%"�F���~���n��n��Ex�N��B0�s�I��W����_e��%��@�X	�a����}��)��{��>�5>}�EHm���ǂo�85�oz�.�FI�
�R��d����m޷7�h��9��8km���
,��	m@��=�_�ڐ�3�Ѻ��� 1�JxT��w�৯`gS\���3�!G����e���]��J�B��QBHZX�nU��l��aQPD,�d��b9�,XǴ(�'#|�[��l�ʒ�U|�ƾ���6�Q����1u�8�jN�3�ͧL���M��m��ϰ�d���'����o֨�`�FML��gF"p�hn��\���M+��)���?��K��U[������Z��D�zc��ؑuB��&ZJ
_�vLƞѦ���Nb������pNj�|K{U(����`>��Qs��O�0z�IM���d�����rK}�P޴hޕ�
(���*�l�4��FO>�-����y�o�q���عC��f)Ȓ���v�imaN�'Q� ���<�l>�w����l*��1T)���7�Ǩ{���6�bM[;�}fL�$ �3P�9�b��8��ϦQx�G!VE�x�S�����������ޭ9	�*���!;{���J��7�·H�%��� 8!b�w����Ź�%[`]��h��~)]z��Vp�H��hQ#m����w_�抍�ca�g��θ
@�i�1&j�,����{�!&߾jM�.�BH"�����Fб �A_ vDI�vroA�4ţ&���'��d���ɹ��o��\����&�q��$X<F*B�����b����T������C���(����H��9�HQ1߹ʦ8+����o��p��lBB�0��{�>3�o�!"�����`��@e%E�,/��Ƈ�r��&#�����:�<���Zz�t�ԯ ��C��H�ɒt��X�,H̯]����}��:��ϱ���''�!�y�c9Yk�RM�u[��y���GVi���s�
����Eyա1^�u/�g#/��E[�F?-v�КX&zk�� A9�vT몂�/�ms�@m6v,���#�H�6�sXJ�W��3�9���H�(o\��/~��|�M!�	�g�h��ከ���ue��m*8*�ܞ��U#N?�[g�1��>~����'Q:�0Ⱥ&��������뎣�a��R���"���
�z�)>��/`6�|�b�Kb$�{*�Q�/ӟ�u��g����Z \��9�3�5!�\�W\���k����Rd�+����!<���Z����ߋƜ��E\�t�w/"_[d���Į�yB��%��� �0(4��]�������|�����.M�zFލ��7q��Z_�w�=^������UL1֑Ȅ��3W�J�� B�:�,�2A��!����{n��e��{�����[�����d�p�/q��/q4R+�,��Y�:P�;fw[D�g\7�]�;�D�V�M2l�qʭ�?d�֫�����O����M~�U�єX��fe�c�SY�b�O�pEI �"xA�W��3f��������.��<���y����7�ȃ��F7Y#QA���P��Wy$	R
��S��;mW�^J;0�vtj]�=Џ">j�?��?_��>im�#��<��<:���J�J��m�gj����A��M��_��o~����=�G�r��0	�2/(*�.�P`���{x�� ��1qKJ�g0�O�B�\���B3���Q�%epH���G��:�%J�%ũ��%�a��[;�i��"%�М���z�9�
f���������4�hi�52�U���݋�Н�s)���G�Ί�Ҟ���7���>yTUｹ1��5��	 @� 	R�H���E�j#��`��9���6k�7dQwyI�	�$� ��`f0ǻ���<�CVUgUW�P�/*�_u������0$�R��$U��R�e(���z��P��*<M���}\����mr�Qi�L�~�7��I/�O���<_	�qTY�������}N�5$���E��ĭ ���Վ!e��Z��
)WN^�2�������A%��q�խO��0��w�(��:��$�CX�-a�u�c��B>P�R�[řv�x�	�l�x�����(�aR�ar�USo���_<I������=�$ru>��`خ~л��f��� d2$n���VS��_��y�\}�eJ4'?�	N|��h�ܔ�C��!:65k-/s�2�%�
�O��#�P��]��U.=�S�_�I�s��m��G�࣏0A1'�LQ"�b<�W�e��q���X+�E�%U~����ܟ�k����X��Y�y�GJ��]���X�B��P��)����i�>!Q!M��c�T�k�%!Җ0��\����rϟ�%�~%����_�u��!�'��%��_�Z!a�GY��Jf�*A������O8z�&�����y��663�pd2hP���^���o�`���A3�]�L��J��	��i�qWw��կ��y�=���&��{�K��^߼��o����ϴ&G���%��P�K�$Y�D"*gL)u�I_-ӓH+^S��ۇ�b����`J��b�?5��;8�{���ꢕ`�W�)JliV�V��~�1c�}�Q�t�����N-x����j�>乪u'g��r�6�9aC�0<��y1c6�q�3�~�G�	(p�����x���AD�o�w%�xq60V�$�l��A{�*["e8+V�q�t��fǎQ" Q-����J�"��o�X���=s;�0s�
�m�c8p�p�����=�[�L����N��;C�B���F�ޣSΠ�J��b�@H����0�����6��{��ɔ��}����/��o��p��*�]��S�P�-H��cO[�lt)�bo�>���R����q�H��5�jH)ɜ�k(�Y*�I����|���o2�-M��@���w:{'g{�$�l�7�~�7�z��Ì�tZ"��R�9	�f�]�#I2�`�����q���4r���W^�՟>���C�����Z��CH�*Yw�B��f/a�9�6H��82I�3��3r����s�Ir����4���~�x��U�?H���N�>0�I�L�������(m]U/8ٰ    IDAT�t�TJ8�+1����ʦ�aL�uҒ����_�E�\����^��������۪�
�� �y�=
Z�uP�XI h�'�E��[���g(MѨ�����J���:�q�4Ƨ�2�L�����uYI����jMp��S��^T&���T��U���:��{��v|f��9�A���J�` ��]����(f@��q�iY2�)·t����ş�%��;`�h\p��cM�5����j���
o����Vd��c&&X9gv�F�)j���]�p�c��sK�
�5�ڣ��B�*?Z�ΞX7�iRN��݅[�z<1�y	r�(L'�5�ȷ��`���;�>�}���ß�,7>�E2s%%��g�z&Y�7�s���$	"�3 ��$G��TJ��~J�1d"K����y���pw�2�d��G����O�W��qt#E��D�Ȇ�-Þ�6f]o�٨2%U)	l6�L�d;R��m5m��daC�6T��c�C�^�A}��z�Z^V-۞�:8����
!�Ԝ]�������]�s癥��HF3����)�Z�Cpgl`�;����8��	���C���%�QF9����`x�'�(6�}��}��?����1�)��B�����@{�G��Aa#�#�\ ��g3�$ޒ�-N}����:~w���W�1J��2�#�hi�J��{��'�ևk�f����{�t�i�y�R��Xl�xs�1)W؀7�6��@�%�`�Y�)O�s�2��R���	��ń)6���eGSu��Y����I�M��\� o�87>��0/1?��/=�V6@�%��ز@z�H��&*E�)�w��`�Q���L��N����q*Y�}k.�S�4L��iȋa,���V(��*hǢ��@D������F�8��0.̃�a-�`�rIp:�c)'� \Z�q��U��X�����	��R����-,��"�N�B�~����l]ά�lV_��A
����K����L����fdG�`GC���6���f���z�p�K:�_��XU���
!lR_y���})y>�7�O��5�`�Y0V��kZ���}��b|52�8s�x繧y󩟒S�=�ѳwp%M�:a0�h�p�"���I-qw��#�UZ��ǲ!W��o}習L�I�����_��$����Ɗ�r��t�ti������u�Z0��զ1A�"��{��>�J��{��u��q����4mq�G�(ޣ�T����8��-�N��ƕ��S��������'�A�{�s��9\��qx������mN*\@J��8���l0ff$��{������l�K����~�c��������h��e��u�[W���Q�n����i���"g>��W:��Mn{�]w�,���:G������I)1>�X�R��6��[ծUZ���w���[��[o䦏܆�<����� Aj���k}��>���j=c�{���O[Ч�Zׯ>MD�9n�-B�}H��D[�㽯$�~B_�� ^�Z��P��C�{lG�QK1`�$�z�G/�V�8�ߢ7_On��	ǆc�J����ԍ����$Ho��{u_���[��]sl��[��q�x�ެ�R	��wy��?�����t���1�Y6��^BQ?�[*wLj]�X���Mٝ���6:4Ğ{���"�]���{?�����1ز@Q ��'
#��8��c�W�%�	f�g�y_:�{��^��?1ȧL6qߟ�n�ܗ�@�)�b4N�N�d��+cq��\n]�[���^���ȯ�_��A�t�q��j���~6ϱ�4˸�w�gS��r�!n�������}��r�����w�	/��`ꘗ���y"�ԁ�W���&o&N�5�}�Q7����oغ�,�]`���S���TAz��NW�5K�o1�l�kq����;��ds4�$#�C�q����-�P�����S��{���
�-��V����1#������#R}��o��������Mؔ���r�S[[-b��g��0�a~���~?������{v��鶃���1���d�y#{'*�*��2�� �kc���b���:�Y$��T��keC0�K���v k	2�����ck�Ԍ����S��P�}J��[G�������x�؀\U�l	�G�,@h���p�׬[$���6¢;6R���(3%I�r;G�H���$ջeF�Z|�_Q5�%�1�Cd��Rx�H�}��o��c|�=|�k��Cw=��P�u$R8l]��R���e�$�F`-���#�E_}����>��O`��lpח���/�%W�!b"�i�0j���#�]�)�jlN,e>\	��>�g ��?�u}j�����_�u>1���)�(�(�gi2�j��:8�_�:7|�Ç{$���׾�-�lʑC���O(M;O��&N �E�z����t��)n���8��Z������4׋!���7+WL����.�ۅU}�b)��﹫��|O��L�+nH�y�$�L.��[��rR0�����Z��sjϺ\E���Z���;�Ռw���0�8�:r�m��-��٤q���>&�uX�B�
	v���k���^�}e�pt�V	�1��JP��-��W8��pR�ta���c��oIe-�P������~��R]'U�'�V�84!�����nWUں�ʍ�\�5Т`��7��T�\w�=�������®v-�쾿O��~��vLh{\A]��� G�w�y�U��}ңǸ��1ܼ3ɗC��r��M�2bK�v��G����T+&�͋���ŋ�H6���g����F9p�A:P6����H��5Ƅ�a:e�
v�>��`�2��翣|���bo��3_�+N=��\.S
��MZ��sDZR}F������Px�|ֹ���Ή���6�\�C��-n}�E|�D�Kл�t�:�B�f�[��)��̟~�[>�(�w��+d/������|�}홚3���e������6{qr��GN�y�=�M��\�՟���^|	��Y��/Z5_ eH�܂K��>&o��U����21>�>����3-'n��Ŝ��w)��$>H�އ"b�E*��+L1]ͪ��!�K�G����Z��,s5�̆�,��Ɛ,QX���E�v���Ѭ+�q_��ω��W���z����b���=��w�@����貃�!�\�Ң�$P���ZJ��n(~Y��cn���bi?#\�X}D��X8���7�o۠�{��E�X��W��a�}�x�I�|�%���J���#�G���&�"�����6��8������
�Xk���[���⶯"ӌ�����L
�l���{�r�y���X�j�����kg�-P�(p�����+?���I��-w0;~��)r�%4�HH|p��]-�Gp��g�T3S�Iiy�}��������B�[n殯�G?�G�^��,������͞Yh,������R���H���5]ַ�W1��w�Q}�.�5�����6AI�̸�o9��ԗ����U6�ٚ\��/~�/�����_=�H��р��
Ȓ���5 ܅�!E�	VhΛ����+����d�"�{������3Pr����,�=m�q��:f���������r�Q3�J%�N0<y��=�%N��1�a��WȪ�dƘ�O�Ξ�{\O��.��oѺ�W<g�ո�!F������l����%�{;Ӭ�^���ս���w�#�}Z�X{�'�����4�2��	{�Ĳ���M-������NZ������o�!I.��⦈a��[Oh�	�� ���[�_���s��Z��l��>�Q��s���3�/_@�%S%���8�^h]�*�R-�ٸ�^����Y�����z��66q�)�_AO'x!)U���:&�2�n�X.#����Z+�c���{�M��A���
�8S��q�?¿�*#�H����<�?|�܃�	J�����>R�v��s�H+� ��4S�>L9������<�o�����fds��4���ˉ�>�^�n���y��5׷��������s��u�Խ�+��{F�����c,�Qf���8�����O�}�8��{��)���߳�ڳ;<&ߝ#���,cccD�=ϣ�/Bb�Fq�$NkJ��J��8��=�<~�ɻ���?��[�)͜Y/|��A3H��������}������nF��O�/�k�m�8u'��&;o�ƅ_?Mzi�P2�䯉�sh��٨z�*&�ö�}�H"g�*[YZ�7~���y'̦����L/_ qv��+gvqV����"�111�kV��V�/ܷ��規�'n�:B��Ή���;��FV{�ǃ��/erj��.��SuP�د-�Z_��8�vU�}RG��$��&)[I��r1��%�CF'�3�ԂKk������,�>w�Fq�c���|<'�]�[��Y�~o�s��N���|���{����{�J���=]� ��<{;�95P$��q���`Ͽ���a�җ9q��p'�{L%��e0�-&�J)����x����8�AE�rnn���_���0���h6�{�i�P�!F]��򜭶sv��c�j����+�P/,�K]��n][~��8L��.�����4Ϲ�S���{������
?���wv�}�Nn�[NI}J�W�t�q%^�W����>�X�F)�����M� �{�˿{
u�2���v"�fM��"�T[�4����|�W��ӅU��g�2af,�q�^��ۂ+��e��9�%)�� ���&t���uq�Amյ��k=�h�^"�x�lc���y.��&���ʼwݴ�ЎM��ʒ]�[����E��ʺ1w�w�V�Ψ���q�M+h8�3-�U��>���a6�T��PEU�����8R*��Qj��ᆂ8���N�q���l(cD�^b]ms�G*�.T���5),�AB�rR�Xrث��
�`Z��3��>x	/����9���0��z.�RJF��5없�D#ʂB�����M]��n�B��b���s"D����A*��H�^ ,L�F�Sfۯ�����n��1��G>���Q�2��d��&'Qi�}I�w��F�+��[;��G��9^�5��a\�3p�q��`+��
�/��\>c�yy���&�/=Ki������ǥç�`r�(�-���2�e����D����y�Ph��d�k4H�Of��eTR`�#JNl(�>�s�����w^`@Ib<��DGըj��E0��Y��ε����I�k�kT��1X��F�L@���a��)��TG�*X��ߵ�7�PU]�["�F�4�h�{�}�xN�F�����vj<�`z\%����㵢�DHp�b�����?�(���v�E~�\���y�im��9���?((	h�`�]ԕ��J��!)�qH�;b�͐唽b���M��1����9v~�]�w.3��J�Ik=S�u�S����b
���gZ�"v�%^I�M
�fO:��4C"-!��'����{�;tG>����^${���)�[�ܔ�����%�ڒ�NXA�4Z�%;z�o`��imW��P�Q�
{�䈢@9�s�F$C,�,�h~��8������E��eFn�/�Z
�t����D��#������v��Z+"�p��M3F�<�vN���o�B4L�V^h�� $�:��x�ph��h��	��U�J���Dk2�h��/���^��b]Q�A�KrWTR�N؈:7%�:�d)����SJ^�-˹�h���ƙ����ն	!i��$	R٪���6'x��^���=���c�8�������wq�=�`��;8~�F��/1�L&s@�dBiBF,[�w��K��8�������CQ��(#x�7����������Ü��n.��c(�9���$M�̧����AmU��[W�X\�۟Xx@JAaC��l�w~�4��u/��I�u��}���u�+��x�,��6��b�����G����n�h-�`K+�stQ��S���5�;���af�����\Ĉ���a��i����&��l��;�ht��>�S���X���c%�kj	S��ߕ,��¸�\�ڶn�ո�{�sK�����%��y�����w����w9~�4�2<Kvp�h:޷���Jq9l��v�p��	���S���W?������O8��g�f�{x�L�v�y�_Ӻ8u��h�Tj�wX�B�L�!8f%\���<�/����������!���Zi�h���S�s^���E�A�Lg&��X繐��qE9��}���L�wp�ÍE���m`�EK�������+��ܷ8�<���W�U�t_�,�@4�����/n��ZWAo�
]�;Zk�F�|ٛ�dٓ[6dq�C�`�m���};��j�\���y�D�	��7?�SK�͸���[a��>%$���S��ԯ9��p���k&&Ś�	�u�4l0c���f}�|O��uj��?M����{RdH��<��E�_~��w�A=�_�2�}�8�#�Z3�Ph�p~���%�R�COR�.a�~Al��� �R'֢S*��9���3Or喛|�˸�[���_f��6~�]N�9�L���R˾�ʸ�c?i���,��3߽L��O�@z3�.��A���[�1�՝p�F�Rw*J���āvR�>b��@
���1����UL�⽫M=��z��U��!/y�����KO`��p�6FCv.�lFk�����b���x�N�!�e4�L�w�#��'���Yr�g��o��;�5�΢J���C�܇�I���T����{�T���J�Q�9R	�)�ؔ��o��o���l��;.���y�<w���p��@����~;�f�VT��H�qBb��_Z�1p�4�}�17_O�L��As R_P�Ev�f5� h@Z�w�[�E.��!5{�fĄ����ba������5o+�.���ϭ�6벪E����xs��(C�X]������񠻎V}��py] �80�:XԎ��A�!hQ�h�Ғ�g8o�	����qBiMȐe	�b�R���a���UZ��}Amۨ�$(%�O��r�5s�	�+?�g�������n&9s{֣�d2���P�m<���[7�����[z�Jp�U ��rƐq�m���?b^~��l������/�9�=�s�R�"�oI��s��gH�B�HLWB��@(��(!(�g�<�@�<#_0ʧ$�"��@8t=����~��s��cz�]����w�԰�O�Z�
j�8"&�
�cԻ�ֶ�!�{NH�I5l�S���w���Kl(G�%H'BJٺV�yN�
��25���0��q����#�F	r�>�z���O5���iS[�w�~d�VR�FXu���cR�P>����K9�k�b�������e�
�/��(ߧ,���R����z+�]K���-60��%BxJ,�#g���/p��i��o���ϐZȆc�]%��SQȭ�_�(�ǺXw�$�a�E�l�j�������:c���}�����1���\'@6v_���#��S_[/������ԌF�@V����1,��jA��lj���;0��nmq�c�e�ֳ�z�(Ci)M�%�u���@��ٸZ}�qU��!�2��!)��W�c���l&)�4��|���)�8d����()W>�۟n������>[(��p%�W_��?���8cٺ�.n��WQ7����q6j
�H��Im_�H��Y��ʑ=R �w�=o���)���t�p��f�B�L�B;Ű�2����ڰ�s��*� �p+�hR.�u�u(�b��=���C����g.�"JG��3&�^(1*R�S����Á����`�/F�����q�2i���o�l�� ���0��f��7���\}�fN���Z�Z��c��v-�l]�ޑ�`*L� �3J2R�Aa���c��؃x3a��3l��c!��Y���U�����Z�����UZu���C�v��çP�r�y��RL�x�b]��9cq�0�r�������7�H��Wݯ�:ƌ���u�w��jO�<ϙN�8S��P����zy��b��b��v�U\�h��	����;��k��� � �%b<`.��q�7�f��7Q�d|���\.�I-BU��]��}}�N�j�Ze{�u�&�")�S%W.7�3N�v�}._fph�M�}�#w��Eo�Ì�A^�+��׵u���
    IDATZ��3�~ݸ��$J`�3���d@n=��li��'ȥ���W$)g?�87}��L��d����$$
�R��1/�$�p�hf�!���ҧ8/$(���A/��e������&�dt��]ҟG�~oWSg���`w�x�o��u�7_�J����)%Z��1��Ue��Di�#�d>��x�Ep�޷��}�����޳�nbn��~�+��f��1�w��_���9�L0+g�$i(4�����9�6}L�*\t \�D���T�gHgH��}��g���M�i�`�}^�ѷ)/�'������K�B,�����5��Zփ1��΀ēJVP��l�'I�r���E�-���U���zm�kz�F�=�V>����t��Z���������wv����f鋛�)Jd5���A�Ѻ�n�׿��/���y ��[����ܹٚ���˦�������h[ 2Er�mL��Ғ*M��7�4���^���B �Z��+���g|x�`:��o�$���'y�g?f2�&�l�~��!�'s���~wzp��/�g��UM��pN	�Ba�^bH%���|����M~�<��QN�\���v�CX1_u��'x��#5�	H��L�-J��$>8aYJ<J�k���(�E�ب� x'���*3P��^3r��$W�9
��W��;+����1���26����bA�}�����"��`(fs|��԰՗�Y�p͸񻥔X�h.gǸ��ͩ�>M�N�^��?�#�ϿȰ,Е?�ђ�%��8saL���C��C$W�'U��$�b���9��`t����~��l�v����;�3K^8�+WJ�u��n,���9"�a-�/u'F�C7r˧fxD��.nB�����S 
[���S���u~���m����y��U4f��;�D�{ @���Q�=}cs�5N|r��šV�T������Ѿ��/?跾M_��9}�o���s��}�����dHa�/����>�_}���U�e��w���SX/P�������4j�`����1���J1/
6�c��kr�e��|�-��g|�3{�����bV UJY�+|"=H*9����xkH��bVX�N0v&ƇR������s��a��o���|}�D���B����]W���\��[��B�(���=���Xci2����ǹnX�e�v:0�2}�6~_{�j�ǻ�d�LC���9C]1� �}3�G���}�f'!�):/�.G����Pf��B���(��J��S�h���P�#ʭ��Q��V���/���'~���S�����m["�`�_�VI����0qV�`���O'f��S����S���m��}�=>x���;�d#�u��W�k��h���>}B�e�W�ջ/LG�����𽨱gr�����{x
��(��}$��}X�}t��?�仇vf��y.ƹ��q��隵����3^}�ŉ�Z�7��RY�	i�M�4�F�s�e	�
��B��H��Up�@z������x���D�ҍu�4�8/H�S��9�+�
�\�P��>�j�*�)�p����5Ll�3�����
��}i=��&���ak�jT9'Y���Z���u�wf���!o���\�ٓ��$g����^�T���sd�:��R���x����w�1'CyU�k�fBh��L����/�T`=�·�%zD�C	��K����!����O�������oE)�5���CvS�wӦ M]��>�Ԝ��4F��QJ4���ۆ��6�p����X/�B���a��(=�,8�0�����dȑ���oq��o�tɑCg��K���gPf��s������$ =�ȩ%�E*��6\m�d^���+����ɐV�l�eY�!4f�-M�z�"Q)�J^�GiAS	�!�D��"�B������V����h�3IQe�rM,��E��k���JZ�;�u�}w��B�I�������jU���u��CkP:��� 쒄��J� G�ǭ�|/B�� �){0*Q�%�l"�Qv�)z���^����|�����S��>�������m�qƱo������ř�<�!�68���ոT�	t�zu���hT���BP�SX�K��b��a� ��A�M���"��}ʝ��}���R�lZ�&B�N"�lj1�w,���2TީցS��$h� ��7�k�`W���g9r�,���O~��l2@�e��D�EҘzMS`\��6�<��CK�l�<0����k
o��ֶz�JJg+�q8�ک�M�apI�����oq.0�R��Z��Tp�ᩄ$UF&^#΅PJ�@Y��M���t?d_�N�_#�{�^_���(�\���;�e����!�_6��D�������3dI�;�zA��7T���,I�LI�4�yl>g�
f��^���i��#������dY���M�VRs�Q�%���&�O�����JR"0�9fyIQV%l�A�&\|��*�(���z��̝�"�t�C���V�CWJ�^à�$����h��4��j�a�JJ�����p���{�)�d����b�ɇxS8.y�J:!q����?DH�-dP�_#qu��7�`�] ��{}>N(���|�c��f�k��V\ם�>8�!�%�Up뻯�7���Vy{l�V�8�f˔Lf�c���t�S�ob{��'�r��	�>� �c)歗9��? {�<[����/wzvny�I��Қ9�4����Z@�e(��tb1Ó���O����W^}�|�D+�V[4>M���>��Am����Y<�t�l��H�I�$/�s�)|If-��mfWv�ΦJ`3��Vb*!�@�bD���>��O]Xt���U}�\�������I�}���{�d�U�M��
����Z�ݭ��S��/���`���o��T*h�J�PIHc�@��%]eu��/�����$�9�Y���I1e�	|:�н��n>K���L"i�Yn���\z�e H����Ͱ8YԆ����wg�#%��Tei)M��J[��|����~��1l�� [�|�+zLi�Y��m���{��TO����8�����E���m�iˮ�#)㝫\���p���c�}�4w���8���q9� 'EZ���=��X�S�%���z,��]�^�tk��`��a�Ols}:�c,#��9�?�~[un��F�,z�#.ۼ�1�C�q���bl�6��c}�RJ��1�����o��?�}�S$�7(������#�~�}��S����:"������+鋊�ׄ�� /���M�(��������8~�Q�~�+����ؿt�$Q���<9�-ێjm�]�Q,��b������q
�B}�L�ds���/ɋ}4�y)�<}��w�Ed�$�"/� fs�T���%iT�]���fn��k�V1,}��6F���%�֛�`�<��Q>���b��g�k7I5]���a�g�º�!�_/��&���u;B(�{Jkp�C�9�Ϟ�$IF�Ɨ������9���:�wJC>��ʜ�^y�٫ϡ�����g�gv6�,
�ʌѷ��	K�F���֡�l�����'�G��늵.|1�@��IS0�9��_c��O�5�c䈣�s��l�\z&�f�&�vh��}�11QlesZ���UQ�����yCY�Q�LqH�2�y�9^�������>��y�v�����������,�ȵ��{�Uw,�zM!Z5����c��w�-�����׵���UHg�s�U
Z5�x�CPU�50X�D�C1E�g3�Ő�b@y�&���W8��/0�:���&o|�8���1��C&�K��>�sC��qe9k�I�ȯj�Ĭ��z�������:K�2���r���[�r���װ��"c�#�*�����X"�MDS'��Z��؈a'CC��,`s�;����r�Λ�3?�>�D#P�M���G{�0{׾_��t��p"�5�xNW��N�`&����8���W1����b�De�sU_G(��,ttQhe"�NxpU>�nE����>w	іqd��GoE�y�LQ2��2X�k�k�B�XV�.sh!������<��\x�y^�'��E|"��Qv1�Ō����0JGP'&Ye^lXIKU[;� �&S��\Y���aD��v޵��jn�dI��GgI��	{�?���.�o��O<N9�� Ȓm�M�=��qܝ�*�{W}]��c��W�$I0��W1o�{�\��6(f%���Y��Y���ߢ�N\ϝ�W�{�s;E(z�U��"y�X}��^K�-8x��V\%�w5��'	�%dS��ܥÈ�뵻n��_uni� �]W�3�������� �G�伮)Q�A�m��!��١��ȟ��?�i�7��*�������.ٕ�l�v�B�m\W��V�7G6����b�"�؋Z+(�/�w\�;Fg��/|���G�y�\����FZSZ�)C��n�u}�}���C��Q���H�h�a�(�d_���N2<��2����S��:M)��8���ЛZ���E��[��ץ,]E��c�����ܯ�<�ʺ�RF�5�S_��	�㦻�lk˖|k�H,:B� D��5���ڄX:�z����q�aƙ���G}��G!�!��Qf�9Zhyhvm��o�fr���2���ْ�ܛ���l��H5��psC>����b8
!��/�����^﵄������Büpg2��|�5^{����d�1�~����^���m�T\E<ֵ���s�.�X%��@��Z�r�!�Z�dB�?g�fX�4�2��3���o�Żob��ԃs�W�Fv�}\	Ji��/ES���^�x�\�A��wh�_���G}�)%Dk-z����R�A\��s�����>\p�:sU_K�~)��/|�>³f=�3���.�������O~���o$9�����7�Av�<[Z1��$^�)��7��Y^+���ܳ�3;��y�0�x��X�0%�sE��������%s.=�o>�k�tJH����l��5�s�M��mPD��m�BN���5��|(Т��y��[��g�:sz�1����+��.b��Z�����t�Ԏ���zL���w����d�a��s��_֚���u	|��-z�a[3j/��T��.�#��,�\T��hԹ��6��V;vx$ߒ�?,��>,9��/�1��Di���ҵ�$u���]��DdH�)�cnL�(���o?��é3��G?K1�7��*R#���.�0��e;�� �f��'X�xs�9u�!�%<ޕH	V�� � 1���'����d�3<s��>�i��[̬i��kU]ۋ{�����DT������j��}	ǵ�$�@!�D�0��Ô�l�,w�A�t.�����%��.��y�����3�O}�wsC����c��T����R��*u��aQ{��Ҭtۇ��W�>�+����h33ײ���a}�pk�d4�D,��tr�5�b�%�.a;=�u�~�[��ǈcc�r�x旼��`�ʋ���[��2V�&�UD���e��F=�.�RT��fVEy�d�<}'�mwaR��d��ERg�o��R�T��t�������PED�Z}�gCD����e�jt��b���3���C������l��E8ϦL�sp�_V����c_�Z�b��2s�ժ4�1�෪8\mF��߷���d�+��t9�>'�%d�����x�u�9Vhg�����jC)��>o��I~���s�Bzr\ N	!f,�&jI�b!Q�G$�$�e�PJv/��_=��J������l�:PJ2-����a��%�8)eS�O��"Ͼ��ǡu�S&� )1�N9�4�[o������'<�>��M�3�L�8�X�XN��m]g���|SkSt���ocJ���nk|�1̋)�VJ�g$��,���D�26M����+��'ʷ�5d�{9��@~��F�R�ա4�����Vק�[��X%�߻�X�s���>��E2�?QY������U�zU�[���/�`���p4"IӦ<�i���{�D��O��|�Hn<��S�{�_x���O�_��c8�8��[��L��ڱ��ۙWq���Z���#4��y1�@q�C����|�R�x��'x�?&�M)˒�ܠ�4�v���%�s_���5m�7c�����'ｇ��c��p�W����ʣ�Y�8�ـ��t�.�ר�kH����ݳ����k��v�W�^��*��y��&�d$d�m�[""#d��YY��
�O�B3�Ҍlsb�;��R/�x��)���S̩m���1��9U�s��)�bXʠ��!Mbȃ�˅�H�L�0)ɼd�dH� �Gy��F����hHjlP��G�<��sr?'�	I�tء��b�8��@2+Kf[Lo8˕Yɖt81��AB4&�:v9�% ���UM��!`5B����ⷢ��3I��x�q�D塘O��T�0��M��O=���'?�5.om�C��49J�7G.�����Y>"@֠$��m��I��͚Je�Z��&�@��ȌDI�R9j�W')����(���!������$Q�����^rx�W����?�G�7IT�������r2�+�U�%�,�+�qW\Q�	X� �&X�/W��>$Ũ��M�u�1�]��CQ�eY1�$ɐ:�� ���E�^�n�q�`K�H`>�Ըx���E~AJ�: �
��&��� fpʲd��+�w�q��Cׂv�x����}�H�L�4��2G����gN1޻����x��'��p��|J>w�J����n���0/@�H���{�x
B�Y[T)D��W�����X���"�dN����l���p�L�����-O�����!�\@��i��H2D:��?���cB��|���%$D�N$���:��J�^vN�
-�_h~��.;"%�6v��;��jy���O��P暡Q8m����p�ܔ@��5���^�8�#�A� �8_k	-R:�2�����,�u���@D���W�u�����M'z':9R���Ysv�����#����sf���j49"EQ$�Eшl�ͦ�n��ϻ2� ��DdD�k͠N��ʌ@ �����l�)�ŗ������!����dr����>+��ೣ
�6����1�3�|� F���}UU5I�]�>G��ې�s��|0�@��3VR�X�J�4Y���T�=#N5���؁8.��lLq���[��~F-t�}��9_���P�N�g��ֶ1������L:���"l��}>�~ظ
{�2/?���p�=p������'�V���`�!�5#���L�`�M��$E�$���#�:�~MG
��i����^�7��6���-�cv��d'�p��W���q.�]B;˙�.-�9tn{�A���G���߱s�t]:p}���K�"��E$���lF�8���~�J���P��.^a�R��C��%1����	A���G�t� l/3U����K���vC�u����.�}�Iׅr���$���/}�vƖ|#��~��6���޵��e�6�����S2QsNnYn����C.<�峯0ί�6u����hݮOO���QM$�
��f��k}9C�r�(�*���'��
��y�Z�]��(�<�fy��?��/�EEG��9V$��a� ql�=*���s�� m*g�\XNq��G�g��a/\�Z��N�q�Ca�k둔�m�Y�|�K���+O�T����/#x���i�Q��Q*a�=z@����O�y_�.�x����ݙ5�N!�+IC�]$��L�9�q>eaچ6cD�&�-��[!��26��x�iRF2���VB��1G�v�Mc��-M���W�⩯�������sӻ���N��Os��I��-D� S�5�p������ƈ��$��%��;��g�R�������a8s'��ܗx��Y.��,��9{���N����^�`�f�H��9��'��<R�!�i�f_�I[��)эO8��$Q �`e�9 c����g��/���o�̥��9�Y�@rf;�j����Jl|�k�(x�UJ�Qj�f�
��_�t���y.I����D��1�C�0�H<6�!X�H���i����U��ZdLG�����NB}&    IDAT��T{�\|�)v�q�*^~�I�_����TY�3�&�N�]�mk}Cc��4�&v_�K��й�p5�R�R.�k��Юb&�}���}r�g����i���s��'x��83�b�D8�����D��ù2:����e��R1QVv(������{Lo����/�����r�$W�ge)���y#����h��2�M��4L6
�*m"��t ׺��#�n�]�8�����ZD:о��^��8���#�g��������s(���s^����4�CL4V%Z0�T�'%�c�w�(�����\�7�(�9��{������E�F��>ǔ��o~�>�2�>�֭���'������>U0>9��kB�4Ɩ�2���5����$�t4}���TC�D�,��Sؾv��?z��|�C�Ż?�y�|���*�
J������1����x��͊B��hp��P'^�Ү�(9#�~>��]�S��[Huȶ8&u���[�'̬F�
�GƎ�P
����Ѥ��C���F�k��An�������J�0Y߇�z�Rm2+Xנ^�]�`��kk��Q�v#���Ϗb�iI������������/��{��\�q�O��#~sx��l���0="�4�R�3�)a��`���c�*h�Ⓦ�ܒ�(X���I��s��GXV�T��y����>2�	�U�t���9�Xȏ�g�?k�;��̐ l�E�)���N0��n��)�g������k&Y���]Y��"�#T����H��g��@��4i�m�I�s�L_����^��+��� ��xKb����y�`](\L�
Jn�%����˅gT�]����R]�"jb�f��tr��u��u��Lb�q#�A��5��p�
0)B�M�c��J{��������by�k/����`Rp߇>���p��A�H9;郓��7[c����C4�'k1sD��P�I^pv�*���O�7��W��}�UE5�s�ou�VK�hT1�䞙ͬ"Ɨ��ٚ�]��.�Nצ?G���j�ϰD��_����c��)\P.J��l��!��U�yx�3�}idh�$��Q
'�.4�	V�8�x��9���O%��7"� ſ;�9��KF�a��PG�hc{=�c�z�5��c�9���Z?7A�߇#�t��U��3�T��*�l�cW:ek�Y��Sq��~ƾ~k�i[d1�E�`# ;%T΢T�Y˄cr�z�{�F�5{�<ϯ��U����X�U3��_�X���F�P��M����k�Z��f�>�v^�V��o���r����M�5^ ✯b[��@���!7}C�h�M�_K��Թ`E�����0N�m<�w�񇃮/�>�9��M��qJ��+(43�\�7�g*7bz�xb��G�fp�~ƬCJ�>n�!�>�7����z�p���̵K���Nu�U�
G5�e~�{����ZW��u�a�ED;�J*�gSKM���f�	�S�H!,2��
}�/~�/����S5�����9g'����� �E�;M�����Z�i���0�#i:���?>�SĵEr�nι��|]�l�5�Rۊ�i�|g�R4�a���rJ,LZ�M!d�o���U��I�4��!�ٔ�tJ��>߹�L�Υټ�c�RkB_�C��!����	[H��!-���x�f��sC}��Pd��K?K��T��_�_���ݱ��;���%�Ղ�z+�L��p��w�"�.#�D���w�Ʒ]�T��jx�� 2�h�Fؗ9���㮏�ݓǐ��,~�W~�4(C]Vށ�G�%k��Q?c����5�y���*�Y���x䳟a>��x�e���i2�l�GC���0D��p�#� h)�g�ch���4)����������k�U�,�e����+�F%��M5���#R�Hg�}|t�l(}b:��gC�dk��um7�}����x�m�9�T�����2*�a��~�w�y�V�ʇ�H�>2�d�x7��?�F8#��N�=����}�g�a{�3)2��pl:c�7O��O��®XZx�����}�+��3r���L��Y޺�F��4vV�Ck�_��}���Q
Mh����T%��UeJ�6艣��
���2���D|RJA�#3�|L�éL7�<�i�<�s}'ʸ���ٟ{&����Z���m/	Ԙ�ۇ��w��.n������Q�L�1«\ŢZ���t����VˊY1i�|g��FF��#��!�#U&�`:(��SYJa�4ӔFq�{'?�y��ԇ��r_|���|���P�2�eL�d-!Ә��t�q���0�G�7t��=Ԝ@�������wr�޻��{\z�g\|�׸PT*
(}e��a������ś,��@�\��;�8�[Y����ӧz�Bu���c	H��BP W\U{f?�n{�6h�)�� ��Hs�	>�6J�nl���7����ߗ~[	���챓O٩/��\}�y��.g{/����kxX�O�0��1���q�nҞ�7>3)f,�\�.KL���)jξ��/��l2��c������ֻ8�;��|�։]�ǟ�Ci<hg�:J�m��ycB�Τ5�ε���]�5��}�f�5�ٱm$�"7��\@W�l�}fk리��&MG��[k}iek?
MH���F����Z�qm={� hb��t�*I�a��m}��3����~_cL}H8O[*8�4)�1>3�e-sC~l�R����WQ��iǁ]u4��x�sxGf����}Z/�u��g��Ǎ����y%{�4�~�S�S��o��#��4�Zpi�`6�byp8�ه� }t�
��#�e����9ř��v�䦆��p�HA3��ѧ���t E�󰴸4,|�:�v��>]+6Y��u��q�}?�?Uy$���H�,OH�k�B�5ԕO�b�-���Is&	K$fue1�`�7)�/�)D�d8�Qֆ�
D�Z2ڂr.�(>9����uM��^�*Ė׶M�����g|�4��l����\�1<ڍ�H�М�D�Z�5��K�	Ǖbo��r���6r�<������?���QhCb3ȝ�ښRJf�	����Y_v2�q芺�þ�0~ݔd�Z(W����Ø���M�J*��kC1�!+K
���;��������z�e.[ǩ�|�;?�i���ej�m]aı�k,��VT��Ρ\�b��%'��_3Y���V��:��?�A<��:�	�	b���,�(2��>v=��2��� ��eB�2�U�d2�21v��R��u�,P�f�gL3��W���o�\��%�\�pN0��D���Oʃ���V%�,���CkE�g�����\(H�N�:��	Ɵ��J���j�@f���#9�0�8�ߘ
h�1��<��Be���:�(j���L \��(��*�B�&8
�"O�0�g������#t�F-j�Z�Ӝ�܂��L`�Ju|V��T[!n�ut�J�ۘ69j��N��B.j��SB-�@�_���;���KNk�_S�2�d:�q��Rm���8s۽��+������w�*ٚO����"s�(��q���)�m�X':#W��p�A�������uM^��gS�G�#�-,
_�aw!�+��Qg��>ȃ��2��
��q�Or<�P�cd��c� X� �`��8�gТl�`(rx8�������&�������n��i�.�4֟M���L���e"P�'X�  y���$���r�)2M�b�g�d����X�Ϝ�N��SNp�VC�ˌ�h�N�B?�B�:R�{��$~?作�3��o�r�6���5���7$ُ��Z�bq�S�,wLUͥ��^9�l���ч9���9@y�C�'�L(�1v�͝M�g��Wja���8cB���9
k
�`���s��1�9fy�K��9����].)]�ɇ&��n����ס�4Z���)2jg�n�$����P,�4��4�^�n��Y��6$�&�ڂq3W_�(5�EI���D|v��Mp�o�m�1��kɰ�DJ��4A�E�+~���\�<�.��0���?��k�Z�y�5�s=3��4��G����ZS.�	fy�V��:��sG���;���;���g壧)��H�|l6�hc�-8����G�<�l�=A�
{P#v���$٣���%�����2g��5���BgT��Šzc[�N�� 7vu�ك)��U��M��D#�̬!��Z)V3G=�V7?�;7��];��|���IU�,ۈ�!xe�=���*1��o��c��߷Υ�9u���"�h���F�`��4Β�&�y���0z��n8Y� C�J%�5�-@���nhrC�9�}�gl�����̱?���
F�Z�I��Q5���'�ŕ_�W"�NR��0�+O��&FS{���9���aYG)�x�l�m�T;>'�-�gc�NS׊�$C����g������V�1y��������b��(�v�<�
ɍjV2*k��
Ԫ��C�Oa��>�O?sVc��{���`WB�����5;�>��hj�����֮Ɋ��7���3߭%iR���ݨ��2�QU^�H����9ua$͕�'L6�!-h����v���g�s�kJ,+�������sC�8�%~}�0�?#���K7�M�4~#s{W�_�)�<ck�$�9�}�����L��ru�k�|�˿~�Z��V�Of!�|=��J�wð��mHp�7��2 6½([3škE���U!�ܜ������CԹc^���E��"'ӹ�O=X���Rj�b�)>ƴ���,^�z�Xw�Z�>\��b��x"��Q�X���:]�B�A���bl�UB6��ϧ>\�Z�1}��h�h=����
��#	� �"8i��V���u��amC̽��3�A���R���*�t�s�W_���_���C�s��?���"Y��JM]VLD�'ݰ����M��\Y�0]w�ki��k43�ZAU.��
WvY2����	��k���oQ����?���{�����rЙC��K�V��'��=��i����~<�ǰ�����m2W���F�C(l��1ږizA��q�--�\����E��͙�+e��Ic�wƟW:��	>�|Sx�}�=7ʸ6	@Cc턲,)˒LkʲD�9�n=��[Π'�Z��M�~6�(DX���c�����/�#�
f��g��݉O%�I�]�_���)�b�Y�u�5��{?ĭ�}UR?�S^���Bv�,;��W5�P��f�n�q�͵�yߟҚ�Գ܉h��}(�͘Mf+�8�m��?����f�����_��^`;S�Y�\7�ni��8޾7����m0��6eZ�5�oe��7L<�?>�	���'�uR���jL8b�G��=��hQ>48�ɋ	d9Fh��T7DE55{ہv�/��π�Q-ո����$7}��/l�	!�J�L{E��|!QA]y��Za>��θ��OY��"R������Zsx�d6͘N-T�r`�#�,;ڞZ��M��6�/�c1�jq������\}��\������'�������~�7�U,��e��P(��B��dz�PWל���M?dn�v׳�o���p��~}��٘�)��֕��j����q�}Bt#�JC�dL�XBe�������w�ocK���)__��,�˪��
��c�٘P.��w�7�@�pn���IK�e0#�D�0�����n�����f��59g�0}��{��0�z�7������/ٱ��@�QU����������x���k���O��.�3��l�}Xo�^f
��W]Bm'���n��b�����7�����^�*��ۻ�(w)L������ ��?��=��m�KkK�Y�S�����Z�{/���p��!��]�0�L(�"��_3��w:d�Z7ʹD�=;B�!��X1���h�Z�f��hUUyM���I���c5�|F�rTF��9^�����4�Ţd��G��z7�L��Y��Bl�E|��P�_
+�3�V��_ւ�wޟc<�o�X��R��{��q�02g��
G�{��2��vNy�,/��WY��g�Ɲ9���'���:���47�2��^
u�|$�h��Qw��ک��3�F�u�X�%e��ŵ�m�����Q7�F�9�
V1C�R��]�Tk̼Yi��R�0FXS&���1-w���t�Mߥ�;�wk�M�(�����k��m̪l�����104�����?gn}�����3��DF�]I�/�坛uHi<�����Pc�6��� �}��������.��\����E��:�s��IQt|<�8����a�\6��5�޵γk��;�`ɨ%êQP��jr��Gc��[�V�Po<��86�3ۚ3�LؚL�"��0.<��1&8'K'�sB]����1+r���o��c�fc{���Y��ڨ�Ǿ�a���J�+AQ��fY6��Y�Ov�c��d��8�w�e})$��K#�:���E�l&ۤ��x�ŏ�N�k�"�4ٖX���K}C����A+���vd�b�\z���ٳLn��[�c\�.�����,VU8&�g'X�|�<�M\t�a$����8��9�l#�sh��Y�5X�P��3jq�L3�r���ᵯ	��tN�ɝ�m��ǋ_��Y]{c+)P��v���P!k딎aӺ=���΍���ڑA�6bֶ묔jM��=���5��
���W�s��	����\ȃm��Xˡ�}��^��a�:�1I�yzdӌdTc�cZo�_���Պ|Rxa�824�d�萢7���Wk�����6/.�ũfC�����$�a��f=Lاi�Ԉ/��0�1�Ƙ������ʾ#{����9�[`2�⳼��`��ŌzKR�"�H��
�v��y��[e��q-�%�;�;gP��w��&�%�(t�S�aQ8��ʛ����|�3w��|Ỽ��Y^8Ǵ����F��s���;e},��ioZ!�;:�Mi����n��l��G����c�/OW:�B�.�`=h0عf������ lR��r9[C�P֧U�8T_{����	�R�	3��K���yHR�!9�w��__�ۄ�k�;�~>�B�rq>�b����Z���ckK�������mV�K��	�w�79��SfǷ�,����6�������3���hSӦ1�ƘƂᵆ��5��TՊ�5TNػx��V�������_=���j�8w����ATqc}h�$���힖a�wܜ����+2�x��ZV)�҂����""d�&+4�$c2ɛ��>%�����6��,��gc��P+�M�-Q��P�\�?�&�3�?wS����}����~�$�i#�DHi��f~Ƒ;�$���z�c�{LS�ǡ���Cs����h���G�CsK��k�i-"��ﺗ[>�i�=�~�3gx�����_��_?��_��H������=�
SW�c�k�c�{ֲ�%嗵H���JJ��(�F�e9�\��T�Oq��q�8d��׹��s�!�V&hr\E��ɟ/Ҥ�f��5M}�Rg����W�ﲮ(˲ɑ1�q�����u2��$^�]���W�з�q�>M��Ve	�͌@�߼��k�����Lk�$?+�\��ڪ	qd9d9���%�D�TcW����ΑiE�Z	��@m�����P����Ө̠s����p-���(P�5Ue@it����m����,�3�n��C���Hm�V�Q)��2X�i��E�c'�(f��/q�s�PSn��>.^��OqKU2UV3Q+�����ْ,"���%��@D3�
�����Y5�q�L�Мr�ذc�R���2�;�(�G��V�4dK���������;Ǩ�.�ۗy��W�:DdI^.;�Ńǵ`�Iȋ�M,�*(�՜�P�kӸ*�e8�kc�E���Ƅ08ʅ��c@J+���U���Gy��a�k!2���葬�Bi�xk��/�p���њ��<�B�Fg�,�}�h��@��4b�c�vX#��m��/�,Lm�ʖHE"1$�FFM�̭s����� kE�k1��.*��8A�y�	����y�9�F�!j@~�[��X�X����$�J��HS>D�����ׄ�xf������i��s����ёH�Ǖh	����E,[҂    IDATY�\��Z��<��U�J��	b�q���]���C|���5��-����^����	���35�վ�8�D�G��ΛL/´ŉ�!9ŧTh����{���Zh��UԜ����s�YQ_-�Ώ���_s��L_��_ǽ�<RW��Ǟc���#�h���R�:��5�վ��rM`o�w�#�X�qHg��.�:�T�,/0�Rc1�0�t���pz�`b���V�0E.�J9��ʆ<�VG�+�/gq|x���4��(�YEchvItU� �-�1�#���ߏ5U{F?$�������(e�D��OƵ�w�����kH���̦�Zq �.�vt#Mōe�6�u������=����L����ݏ����;���X�+��2jV	N+$��o��pB�_~Mx��US�� }�b �֙����-\;8$�Oɔ���sO����E���я|���_�:q�l���\pz��!j}l1n���K�u�[�=�HHǖ�����9E��O<�3&y<]=ShC���^h��6� ;�/l7렸4���e>��r��7u���c^��a�%l�v����~^���Mr���W���1ؐU.��Ɲ>�%�9k�#�}z�ZC��5x��n�.��3f���kB�H�)���-p��,r1��R�`v�ny�}TԜ�Ѭ�x�7~�E>�0�+�ѧ%����ҿ�1�m-c�m�S6��2�&,qJc�NPm�ĉ{��{�!�*^���W?�!���L�W2�)����c��t��x�O�c�����4�v��wS�ԫ�o5�a´�e�����<�黺<�K/�,V���v�-�Rqs��&͖5���[0_L`�0lF�7�f\��(Di%��(b�r	3i?;��H��ݮ�B;P��V%��>o���p��g��ӻ�����p� '@ؿ��ju#�Љ��&|fBߥQ�	�_ǡ��{UcR�'
QJuj��C�t^���R9��K.~�;��w_��/P��}��'���¥|�+�0�![VLvOx��xӷ�N��R�5�1��퀺���y��H�C���������t�D@pު�׎��sA[i�E�ͨ�:�h�y]��zm/��x�m�C�uN�~�������yloѡ���t�B���fl�O����0�\���%��+؍�(mk�z���9Vg� �d\.�\���]����ԧ�OiʃWy�{���ϟ帚0��ctㄿ|�2F��m���xR��s.��V!����A����竜�-�q�����%��/b._b�s����*�fX�c~��n�s�M���k�!�fYA�,�r�ZTL�B�Ey�:_ds�ɱ񷏷�]�;���^l�a�p�	Y���N:*�G�X`>c�ט4�^~�ZF0���z����5��8�Ƨ��C���싿�7��&��.P�:ͣ_�#�[倫�\�PV5��������Cĳ��+�E�|0�)՜�E�("m�������|F�*�
n>�Cv����7x󉿥�r�;���c��ܗ9?;Ƶ�a���g��J�����Wc���}(<���7��Я��C��p9׉E���[�����!�Y����m�F��Z�kۄ��!���D�Ƙ�&��F��fa~�]Cc��0��/��{��Sgl=|M��f�w�����hi��
�W��:eNCZX�5[�ǩW5��YU���4�>����/�|�2���_��w�`V�L�������$rQ��D�˛���=}\I��ZMhjl�&3d�D��+�z�����(�˿x��g�e�,�u,J��'�25��Xǘ �*��o��G}����f:�l�S�z�Be�l:!96�4Cvw��<�Q�La�~�����]�S��IDQ�pN�����F����z�G��� �$���O^��3�{ߍ4A9	grґ�U�����I��g�����F�sΟ��N�t�?G7ׯ�����E8u'�{�{>�Y޾zs��L�XGFP�c�@o}L=3�9�uӼH�j��a��g ��dV�����Ĉa6�µ���_�����S�O����1���_��� �	�0^���U����g&�\$&�ǭ���z���9����`0�ڧ�m�����[�1�oC���?3v�5�@�I�$!�k���uPk��%��=�n�jcL��}���������;�=����l��i]H����E|�q�Bu���^CZ��O��qhDM���e�H�����86�Cp����:^������e�����L���t��n��?�I���_���q�α��,��u���ww80���s׵Y�a�֎k�C��W�6	�@S�U����l��Q����z��������]��w�͕�<Ǥ�52��󌕫�X���I�ӹ��o#�R*$��"�����C��^h�3�	�5��o��Ϝ��s���p���]�27tgh�>�!�B��K!�4�w
���hёHmB0$y��I[GB�}�/�86���y�@��3͉�}w`�1����F3�y2/a��:ɿ�N�gu�M^x�p�L&�y�)��Ɓ̉���"��\p��ո��bmV<�M�M�P�|\� �cO&�)0�ú�T�ܔ��]�ٯ�{�=ԵK�7�����S��B�Ga�XQ��x֡���qN�ZK!�\8wWm��RɺV�"����e��/�qԵ���>g15m4���^M���3��>�Q��(�c��6�M�k�����bӻ"��#e�}24��wO{��}*��[W(�l��<����\��c�ZYU���b:?ε���{��c�ޛ�v��WƫO|����8��8Xy���:�O���oԛ�m��o!��]k���v5z��u��������>N��ٗ(�|�i�|��"G�
l�1ٴ���J�?�ӯ��dl� ����so~�.�⑌�c:��9EU��
�L�	f���������^�HP��.�<��i���`���
p��8A2�f�t�G�#�$JY�;�Z�! `Z&����$�.P���ͳ2�����Y*�s�lMi�Xe9����3O�ؿ���r�G?�խ���Wߋg����Ų�#�7��+&����""D��Y� $^p��%�4�@��Pe��&F���,����cs�/�΋��do�J�*��w~��l���?Xa��U����ihӵ:�[K%BM?���Ou�}|.�!��PjW�8�Ņ;����/\��Wt�c{J�f����1�z�1͔Цi����}��%�w����h�.e��(A?M�}S�Ji�����`4�	Y����^B���<�o��G�-�,Ϙlg\�+.�SL�-�{o�./��������q�����%s5S`�ͻ���1��6y��Z��b������9�nzN��˹F��ӷR�~�o>Mv�M���_s��癉f�ZQ�5�\��*��<�
"c|g/�|T:4��O��x���������(��)d��{��{�ư�(Vdx�M��Z/����6���x%3І!�l��y��R�$x#˘T�~�I�N�SF1<�u`7}7�s�h�#8(�8�).W�-��/^�K�ȵb9)��#���t#
�3�"`���5	8bB��>��u�O�Rc?@��$�U�d�j\��X��W`�k���1��ϟ��'��w���]n~�Q���:s;���G�*�P�� ��m�Tc�`��k]��#�t�ڽ��_�#V� 5�*sd�����_�,
SCڴm<�d�����i9�~�g{���~�H�D���ƈ����[�@ژ����1X m��;�����Z�Vdݚ0�|�W�4��+Պ3�� ���غ�&��%�|�\�ַ�r+��q��)�	�v\������r�
Y�9ƪ��u()����_�?�(`ge�u�y���͏�����z����E�3��Bx��BI��bI��yƘ�&�O���2�5ĜS�1����|Y��`1��
�w��A��Y�&�Ǘ�+��l�Z,�QfQa7�����ۣ��[}�O�ςF��&Dy'$�|A__��ly��d�PV��Z�'��$-S{�j�6Y����߅I�3�
T�׎QSm�T��18�D�D���2�q>vT�����3��Ћ��S�>��g]��ו����W�'k-Z���$dL�WrB��*�N�ˊ˗^FMrn��Q���{O���a��s�.���fS�5�[s]A�@C����nu]��C� 5`�n�O۰E��Aa�:?� �t���������jJ�ԙ�ǹ\g&s��>�.���Rغ��:y�c7����y��Kc�l�p�c�K\]1Q�!��v?����0�&�:�;\���m`��F������pA,Jm[	�_
<�&:F=�y�3�M��҇;��\��С~|�k�7\8Q��:&&J���ͺ�3�nb��r=�_�W�ȲI�.�s���k���9�$KjL�)��N;4�5R�%��i�?�;b�l�
�������ՇIW��{5��h�)1�'Il���}0`n�(�|�K�Θ��p�ykb��4�`�C	T-(����V��v�\����/q���?tY�׿����������h�"�R)��B��ϳ�b��k�e�RhGK�1���cB�� �5a�,����Rv9Ԋ]{���c�/�O����~�kO~��3O#u�Q�4�
9T��lN��T!,V��`@`N�Y��Q��b�X�K��ujQ���A	d�m�W��ղ�.N�v����92#L$�hŁ�,�3Ϫ �YG.��v ���Z�`��[e!�X�vhmP|�b1.�	ˢƸ�+{�n����F�P�澔�E��}����ퟅ�p��0Ԇ��J�����{��t�Q�����	"����m~��
�l����y���y��%�����ũ�beg�I�U������eI�,;��5��x�A�M\�N�co�u�SN�t��k�O������?�z�nYVh�x�������$C�5��h5'��r���ޙ�c�^(X$.�q��&�1�X�����$Wi»��~Y�kp��φ���6ͦ��𖀡ȃn�~���W��'6�l�Zm�$;�q����t�c�=�|.�5�T�흴!<�7�;C�}O���%�K�����v�
d�@�ɒy>�P[��7C�{����/s���å�\��S����w��Z�x���g�2��j�y߻�1q�r04�� )�����,���l�6�q�3�듟`z�	
Vԯ�����>����Ǚ����m)̚,�t�^�o(�J�6�����;��iq���w����j*-j2tc�<1@$;�I��I��k�ĈbC�bL�������	���S��g���Y�Q��ZY��7p�&�8yI�$���
�3f+���_sṧ�,��.�9v�#,�)R�l��-5L���c�cDoh^C}nzG|ư �5�Tƕ~�s��~�C��P<�(������a^Z.�����_��,�<J`d�ݐ����N}��O�˄�}���z6}OJL��t���=ݵ�5(�ڽ���������	�C�2�}��X�����̾=��&qR���[li��)���#���D�����C�l�|��r�`�����ȿ��)��%�k/��_�5��3�M�Mƌ��u+;�棁8�a����[lk�ʑ�d,TI��1s��}�{��s�a��c,Ͽ���?E]<Ǳ�)����q��<������N�o�p3�%��	.��Ǆҡ��1�y���eY�u�n��1[���W4(o�s�16�5���@tX�| l`���Bt���
ª����:}�ݔ���0�t<��crG0�8;�~A��}�y;��"�
�,�vvٻx�W��Ln�n{'����)������l��� �m=��J:2�!ؤk�_�a���3�Zi_+�֟`�d�٧�D�wg������{~����4�g��4��y�$3�AM|x4ޣ8�.��>0����1��ǘ%g���b�Y�J�f���g�B�OA7��0����,���3*��C<�`㜷Z��}���敶Q¬"L����N�(p�%2��~��g	�fP��`Q.�jE>-�+W�I��?�sN��^Vn�������8x�i��9F�ո��os���I��;�� ��C�@��nHp���7aYZ�iƎU���Os�]�G�v��Z�ڏ������+)�����w�c�}L��5=���HB�mhz���U6�֗�h�Khe�L��J)��kC�-u��Ąt�x���0L��eYF�~�ZG���:���z�>��!	��[;;����?�'Kr>Gg�y���K�Zk�D@ag��J�0;!�69�]�a�`�.�S��-)��I��	�e��Ρ\p��p�Ǹ�{�>Ql����wp����R���-��!�e�rt���w#G�k=M4S:�o#��A(S�����L�s�+��_��E>��۬�y}�����y�o��+O�-��ʊI>�2��߹��֧�켏u�"F�6<q��+�O�6��1省/05�㏿������)u�"՟[� �1@�y��wG��?ӣZ�1�
G�ŏљfl���o]ctL����g���HF�qt�U�\(����4F4�����x��{�=~yQ��/��W�?�|���� b9\��'}�4"E��a�2�����_�+�:�����*�Bt��-��(����s���v~�}���Y�=��ׯ0�&J���i5c�GDlRR�\�����ZS��H]�W�K�& !S� �$XK��
Siuݵ=�߂�Ĩ�KSO�H?Oߕ���p����΢z�����1�Ēz6[kq��FS�%2߆�'A:�!$�ZL_{�ݟ~M7�?wE�_T��;�N��'�}����'�����\�q\]	��	���s?�>w��Sn~�a���/rn����W8�������mW¦�Vc���gL88R8��m!ͫE^
��������_��/g��p��������������um��j����H�)���H']�27��w�b��Io��$-�S�i�m�������Je��ű4��k�ԯ��|��CM�}�-}��Xߩf��od��%��>�_�����~&�>QNi�;=JH��S�G��}z�Z�����eQ+��S���q��~��?�!��Ex�^��_p���ㄲ�ιv�@������c�#l�F�m�ѽ5ڢ��J�䅠ܔ���ř�y�3�ǩ�<Ė�̅����_��-)P�)ui`e���Ctip}GBK��l*�{;�!�xA&��6�2<b"�u�9� u�v.8��F���K��tc�\���Dm�� 4Lv}���Ûͽg>����e�㦤T����$*y&S���D|e��ǃ�P�	��3�W�k��dLjm��-�I���⿰,�fU���!c����"o����'���O���*�}��35+�&��1<�!���:̇^�90xf�_��9�a��V���7�a�p��O�-��<����Z��N���"'f\���Q^���|�9%��\L�Q��d3�M�<Uk�k�v��Νw:�L�g�O�G�쇄�!������g���`1r�Ws�ꆩG���c׈��$e\��هC�_�W)�<�����������_{k]����g|G���S�!著I���Y9��KX�v/����S��y�U�����w��s8�V��[ԇ��GҎ6����m��-�7:��?H{K)w�Ö�<ӬXrl�ѵpNg�=���<���W�ý�f�%�	a�Mp2A����؎y�r�����j�1*%j����a����؄����1,jǐ�7�	�m9��ۡaD�r����@�O̻�x�y�۵>�  tM�cE���}?����%�����#��xI�H�]�ˍ�V�[0����.�Թ���E͊
m���7����\�~��v�����n>����lM��e=�k�w�]:�>1�7�@�?O�*Jtf)�_�X6A3aoU2��تW��ķ�ɿ�?Y��,�-��{���Gq�t� :��V+�����44�M�",MU���U�����X$)V���U0�x4�����lِu����{u��0#��N`�%�C[?���!�;�ߐ@t
���j���_	    IDATyn�tܣ�����B`)�eٔ���^�L︝G�x��?���\<����7x���]���ڐO&���t'�1�\z�s��La-T}Z�~�y!A�M�Q�Pڐ�c�>� �mۨ�>O}����g(�"Wt�)˚W�FR��	��h�����oY�$;���(\t��*]�!<�W�~��8�Z��qd�r��5:/��ХҒ��$�L�1aA]� �ڊ�6�,cʼѼm�l�/����Oi�d���f�c�v^�RJ!�g��9��#G,���ڴ!g���FccpV��Q`�ҟlj���bQ!	�1����*ԖV8qDW�Xg�tA�"����i�>��� [g��5��uY%"�
�Ұz�^����������{�3��S��'�/������Ѯ��
$'�B��\���B�ه��GLB���ƿ'�S��c�L�¬�̂lR�����黼~�*�<��g>���8y�.g�-4�y��1�Z�$�T&����PN�~h��e~]�ʇ�eY���t��߫�sː�T�&��
�VA��L�&��y�j��5q�	��(���z_ ���ڄ � $艄�;D[DY�E�=��-A隧c�N�KǛ�ј��oDa�m�lk!�@�K�-�>׭���1��3�$濖u��pA��U�[?�W��G��@��G��X����I�rJ}�;?�g���?��\���O�������or�\�KVY�9p���xt��>��4��[k�ja��5��!f�ME����!Á����6��rb.dp�nN|ⷹ�ч��^���=�;��N�,ױY�������)�����u���!�V?�5�����lr�2�}�+���kqRD��k�܋�y��#F]8	V���
$�1�$��I��C�ZOw�����>�"�8�k:�?"E�D�����-�U��[�U��>ý�g��5�ZB�@f�Ap��;����
"����_����HB ��BRwK���v�ΰ�����9TV���+���=T�+הk0!�@�Y�8_�1�c����P�E��4����}f	 �{���
;bR4���fD)њ~�[�C��Xs�2��B I��$�%�P�kƪ��d�mbX\%+�Q�
�[�J��gU���>0�ZN��4����5o{}s�G�)n�ܾ��,軖æA���=�r`�x����v��$��wS�t�;�l�=��0H4�,�
��K���;޽~���	����"/@h#H���ӎ����E~�c��8�;�FL`R���g�Фi'+���`������_�ۓ����s}��/�o8Oc�<^T�(jb���I_��>?�}�L�������/.%B�l��ь�/��TS��|5�l	�Hgsq��e�̑W����(�o��9�����+���O|��?�Y��}�����J'SC�{.��.�;|7��r.�C4vV�����s&����� O����_�<~����/��7K��-E�6̫C{eQ��Ka�.Զ{4����
2=��08��50SF�Z+W�-�f��_Q{�����}u�1���=N�t80��b\V�)!�(��Za��X��T��A��BOBv7H�+oh��EN�!`�0�f�<?o�\�������8Us�6w�����ĉ������5����5���˷����x�/|�x�%NN^�Y*�JH�j��)�R����TҟJm���s��\QU��C�ʵeO��/����n�1����>�����Q�(��cI�)�/"�uP�y��.�c��;��D>�g7Rm��)-��3e���o̓�:F��yL�.xU�x�|6R�0sZ���}k4��>��^e��-� �s���:&�ވ��nƻ�+��Z�{��YMc�C�?�F������~☛��./��'�^�9��n�M�&��ߨkX������YNߕ��>����1T[a�pۜ�ڣ��=1��x�>H��#l�>˭O��>�w4�g���6����D�"0��Q쓋J��4��NҦ�0��ikPd�aե���D��2���(�)W�b����id�,���m� ,9�3��.�RF��Qj���5�&HTY��\����I��� 9���9J��01<�j�����	a�S֎�|�ƈ{l���6%�Y�L����B��RY?����?�]G��=�v��_����<���/��7�8A������c�}�t?��IES�~�����(b$.�}�
�Ê�U���-j,rP���6G�*�������RK�8����M��}��2Ե��5Ɯ��Ρ\��y��/��b
L��dO�]jטj��$m%	��<��>�B��[��Tz�eh�Ϧ�]��H�ͽ�V��$���1}_�̍��6u���������U�|*^�uT@��mMߟS�[^���y��b1�9ˣ%�Q�5x�$ؙ�u�p_��%�$0�v�~!�%f$�G1�ytq�����w����E��������>Fu�6K�TZߡ�BLP����!ND,���2�6��ӳm�$(�^+�ӕ%xj��XSJ~�1����&m��b���~i>�9a�����Ԙ�
. ��5N
�U|..�d���X\��Φv���D�G��D>��O9�YU�J��3|_J�Z�+�B���|6�`�YIr���a4�))�0��!�d�r�;^����ђW?�ל>��OѾ�M��C�ŧ�Fw��U� Zm����Z�&~��HO�73_�P��;�r�齉��t�7�=�����7�Su�]��h������Gb��{��!�@�S��4���3E�ss�[�dݞJ)Mϕi�۲��~�� ]����|��>������u�<S)�
��E�_��ynF����GR|���R��D��Po>��H��Z��+2DZ�H[������ �n���X4+:�,0��^�d��wI��V��x���k�1 �z
 ���!7Ϡ}�-��7�����^|�+l�}�kG���=j,^ޥ:W�t�"�>.��1#�~��w�aA����Չ�ԩ�ʥ�$��%9��+��)Ǣ�E�ke��Ąs0\e��b�Mo!�6��on���K!I�	�����o���Ez�@ħ�����~���9H^�w�!��e1�䧮c�;1 &�v�~�V��;w�s�CD�]��
�V�v ��p���/���?�#��ȣ4��Gt�#�� �~�K�g������o1�����#����͕}���Mi̗����.�ﰨitI�g�;G�[V����j������w�I�r�%��{��5���1�ٝg(&s�a,a]_\_��6dzJ�c��ȃ�ar�+��u��hj�]�Q�j2��͕�v�2���M%�9��v��z2�����Ź�f#vD�GUh�0��$d'���̠�>����z��RU�η��W1�(:1B��kC�r���\;�ʂ~]�v"H�k�d.-���k�-���'w��_�����9\:�]H�䍆h�N��c��bg�������jM�Z��v��n̨�ϩ�HW��o���m2WgQ���ݿ��D?'�%���s�^0��ڠf'Sc�?�#L��0W���������Ġr����d�nssHj,�\Q"��N��m�'H�y�lSv���8�J�xw�&�;�@j��T6g�2&$�	F)�
a�^�{BsPs�{_���>������� ��~?���f��
i�X�.XT��LV9�	�{�����S���{lkB�(���z��U���.��uOm���BB���~x&�H(Y��J�����ss���%�q�W��L�~ڶ��&չhe���^���[u]cL5���{%��55�ۧ�7�r���s�\Df��R����=+"9>�(F|���.�{5��Ƒ�$�*\�ؖ�1x���6��);�֓V,I�j��v<..|����T.�7#�%h�<�n=���_����Q��UN���|�O~��o���sb(UE���b�"�c4h����hҔ�.qOb������w����F'�F�I��-۝�ŋpo9��^���L� "�f(�Lp"�+���P �9�'�T���)$��C��G;�D��%ԋ	R��6Ct��M����EE2���` ����3�$�D��UyU�C�ܧj\&�c�:ǫNH��<l�ʩ�y��#�����~�;y�/����x�W��p�fsr������+'�6�5I���ا�[��e�?�<�1G��_�dqo��?���å�JC����Ծ�	����#����_	+Sn9z��=q)�u=
:4'��V�.pb J���|k+\����UU��/�b��]��JfRC*١������Ü�az=���͕9f���"��Rm��g��4��>�l�laε?F�����̵��c!�����w儊�`!V*zk�V�lO90��6�������%�Q�{V�7sD}4��}�x���|����ł�+���_}���f�p���rUU� �,LC/�s=jӽ�a.O�����}K����$�c1�(�)�RE�?f�T�����^=RI>�F鿠���M�/�{>�?s��� (����c&�F��
�@^5H�\��IiT+�t�U"�Y�*������
	�&"���Ởj}�=XS�.�.�`c��J(!	<��Ì�� 1;�`��,)����\Nr��}`p�����5�9��	m\����E�ǩ"����p@�%1Bu]�	#��1lkO�pv�cۛ�|�/�{����z����7�{����y�5�U�ӷ�������
��&�w#!��i\��87d=H�l	PS�����:�2]�*H��0X��.��R�����,����=�@T<b��E�S�C�{W0��>x]�B���wx��&X�2���{��t�h*{����ŀ���E����h�Td=��Ӷ툸����5.���$ԁj�]���뚪2����uB4<q�51�2��2��Kn���H!Y���dM�����)�$2م�Sºs����̓*�Q��xB���|��lP�db0e��=���wy	<���Q�*|W�Ӟ^� t&�׉���qJ�T�{��:��+��]��{�d�#��z���rN}��6���H{�s�W��z���X��ͬYS?�-�w�fs�|���r{���]�5���h�%��ǂF�z,�Bgx�*��Lp�vށ�uo�J!dvC��� �K��H�Uk���<�M�K�P�U�40�kV���b騰T��P��S���m�!nˠ����waNA郋c�U,#`ZϦ��i:e���}��1��
+�yGi|�S	q��-_�Ԑˑc��5���Ч �$J�<E@љ�w�4�&�=��B@����d�3.��S�7���pkk��
�/>�M�>���psL��w�|����o����]��}�s[-���uwI�d���1<��Cbf����O���):I|�z&&gN����Xd~��<�S���2���w>�f�;!G�|��kۺ�_^���;�� K��Dƕ��<8u���?�*�L 7aDw3�ͭcXK�<Y�-���F Y)G�"�|���������t�$ ���d�qQ�w.�6\$�_��T�37���N��&�`t:
�K�}_�\��D��"��>m�,���qS��Z���k��V�*^���G�ɟ�0���,d˝o~��|��>�]��%�gT���1Ɛ	�D�>��W^��a:׋�x���1	�b��P'�ݘhiC�����@�0������ё�_00e��U����v.��*���=18W�y:��"eե��̩٦E�8U��Ǥ
���`_)9��{;�Xz��݈Os����*��yw���$x�ԔUM��l���f��p�K˷�7<���r�=?�c�?�s��q��T[���0|p��LѮ+�0��zw���!����5.	�t�����·]M�����+��D���z�b�M���[��L0"4U���t94��������֘�:��YS#b�V��w�H�2;%=	Yx-5Z�G����>"��tO���������~ѹ��=~7% W_*%�O���o��ٹ���N�>��G��ֱX��¾��}N"�q]����׫�^k���~��y���
�ut��g��8g����g�����3����&�(m��pU�����)�p?Y�����r^s��\�w.x����������4gDpy���YZ�a.��31�o�;��Sx��<`k��}?v����Jq���؅��� H��"^|8ǜU>ޓϩ����h~�Fr,쒐@P��b�DT��Ҋz:�4�h"���/�7OȘ�{��{�ł�)/}����ħ����x�g>L�C���
\[�u� z�}�Sv��9�:���e_֟�M:,�&�������w������?k�l���TR`L�h��E���&d�&�������˃ͲFj�T���������QR��?�%�&�כ:ܫ���N�2�O�W�����Mg����9,������'�r�*��ӹ~��\_����YAaC17���5��$}��O�uQ�?Ș�u��ܾ��#ts������g<�<⎜��5����Y���x�~�Ճ�=y����/��P�~�jQ���լ�|Ps+��W��oSC�M��U�Îv�`ZJ�6m7�m����fv`���Nr���%��~#Ќ�}A{��\w�̫Q#9��E@<E�T6%��Fn$���}ȼ�nR�������J��:�I&��x)Bc��]�X=��C/ۄrN�J���;��a�esz�=��3���?��_de9��M��g�[�|�=��B(T� ���\x�}e�Q�?��^Y
���n�$��mp�!��	��kM�E+���Z�7�7Bo����lRi��,,����a>A�����%!���t��2���}j��P���q?���Ra[�2���x��X�s�ɋ��T��WM�;�v�D��Y�,^x%%6�l�W�s_�G�J�z�އ��k]����镶���,�l�������'�+��x;��p�����O}��g8Zm�8�v��2�/>.�Gю��q���uwΏ�ǁe	�gz��>^4��~+ۺ��k�$��k$v좓�t���Ui����H���yN<�n��R:���9/mhFZ�X�~�Y�rh^�����n�"���f){$9��t�S55�w��ŉ�{�}����|�t/=Ks���۟�-��l����'�d�ӱW9�9fgјJ����+���<#�%�����	�r|�2��]~q�#��`%h����鐝-ivD�n��n�l�[\�)Y	�����ِ�D��=�#��*dtw7w^��8���1��c�*����\\����$�DD�}�XK�X�Z�v<ʿӳ{/Du_���e��em���xG�^��L��}kzB�7�������1x�	E�1O���,�ߖ��Ю�����z�G~��<񡟧�nٞ~��_�}��,����I�>�ͼ�'��]�8߾��+s�F��6��c�)R����*�4�)m��ѠKte��L���3��U�T*1J�r�HX'�+�)c�r�T�;w�Ge�tR�K����(	��و�n�?"@542���j	F��vK�B�ڼA����a�̔R�,Ǡ�X�X����,Y.W8u�����|������x�g��Ɗ��w�_����?�HuJ%1q�bX�= �m/�8�����]�������8�Y��0�o�|�s�,�5�> ��?�p{��`a�|^	�C:7Īw�;*�[�tơ����B�Mc��S���o��֙v��N�Q��mJUc�E%Eʚu��S������t�st�����1�?H��g
s}��/� �w������X<W��~�y^���>N��2��g��8���r�ִ�Or�}�_�e��ø�­��%/��"GGX���eiB&�����D��B,��@1�iE����N��z������)�Rx�~7���:O��������V��}�^8ki��[z����<��� iUh�|�SL��i	R�1�loc�q�ݝ��BN9J"LJty*8�)!�
ף�Q�Ϯ!`l\$4cs��gDm�w���T����4|    IDAT�q3�l�+���N� H{e�]�T�e}z���c��ҩǹ�����%�{�|�/�������{?����~飼������!YU gp�]��/�Ka$/B6���ًi��w�r_�a��"�bNz��j�9\��!ܲFez�ĥ�U��������86&X��"->���D�Ẏ�Eob72'���y�b��9D���0�m��g�\��JJ�ĻyE�.�2����Z0]W%bs{u���Q������N��@,|4z��-��������%�+�;=c�$�����a�V�sM89��|���������nr��/��'������b����9+Y�t�n}��p��]�+��$�����q������\s㝮S�}"�F5��n��D�<UC2��c;�l�5]�b�B��7~L����qtY��4&F��E	'L�rm��[��ҽ�Cv:���x�����m�F�>���Y����j�� T�#Fh�kk��X���#���.����`<�+tQ��<��[tU*��1�S�GW*	���]^��NmY�B�U���m[���я��I,�A��r�Ae����+S��k�b����(]r��mϩ8z�AN��5�����-�{�G����_�o��K���?���3�����Q�ͻ/�+��`&�r �1��%S����5��]i��{mĂB���z��b4�KU}ι�����20���<����� 1��z*��ƺ����3I��#5���p������*1�����t=�"��V��C��U ��YF*TM����"9�yx��aL�n����A�(�S����b�Ns�Ho���g2��q[�!�Y�5���#�f#�4~�8>��2���w9�9�]�qnls㞫_��q/��>� �[��N�b� "@ݿ̲]r�3�Xh7k�׎���~K�>J��c���>�я��~��?��{l�}�8�mN�{��j�fCN��X�X�����e;��C��Q���W�dӚ�@/$����.�>�=H�d%�2f:�?������{O'A�g��{�S��l<�fDpELV�W~��6Dzq�*x�z[j}2�.H<��XSŘ1b"/�#8y���u[:	g�rE���o��Ԣ���9M�+P�$�&�"�eTlD���A%��$�M7S5���|�%��δh7��� I6����ݾ�ji��w��?����B�"\$ �HUa�;�;��uO��8��恇��o|�;��x�c���Q�>|���y�l���O�����sn�=�z�b}f qq���������R �5�s�+%wӮι�M��tf��)�6NGb
��!"���"���,���n�ԧ�L��(����V��6l�g�ES#��c��f��p�Oz�+sgh:��o�����b��^Ƽo<W��LM�[���ڍ���M��]u|W�U��G���:�s�_��3d�Нnx�#�n��S�8�w:���}<��[Y5�o?�w>������,�B닯s�9�)�`'��,M�?���	��~8K0������x�0-� ;)~�)��$Lq_�a>�H��Q��N4�GG��s��%���1�lb��8��
D�*`8��r�@�߻*u~���g�9�C��(n�ΰ!�*�E5��uEP�9e���������G���ހ?Xq�u��� +�ylќ�W9����/�o�>�����WO96��e����.<������#��g~����c��=b�������}}N?�:3�Q��wɗ�<[qϼ����WZ;��2��\"Q�xH�_4��Q�(��o��㻽]c��*��~��5�}�4���Y�	%�a���U�����\�򙫔}pQ�w��\��U�����~���9�Kh�c�#�W)1Ws}]���Sc�����ss}ϒ^-����4�u^:��O��?���{���K������/�ܚ�9�둑�[�S���&�O�J��,��L	�.���_�#c�}89��x�dc��s}�r:f˰s�e�0��1���wf�6�W��'9=��_{�0�.o�#����"M���9�\������$�Ka�PnX��}�x�O��#pn��
>��㠩�ڄ:nw|%�F�`$�S`��7���CL/;�����Qy8j*��3n~�����'��g���}��?ã?�k�^>�ik8>�N��ĝ�H�M(e��C8�5�P5y~�L�j��!N���8�S},�+��S���C[���_��=^-�KW�bv73��'XJH�D6NC���Z��u=ׯ_�O��ŵC�J|�{w�}|�����w��!�To_��+����Ua�,1�������(G���{_š;m\4���y/��ϥל�L���1U�fq�c���z���pTs�^q��;x������	/�S���Ϡ''���g=a.����X��7��%���s��d|���ƀi;>��7����t���/��;;ƿ�]������kB�6��U�-�B(�;���(�WD����i2qF~�.Tw�y�)�ɀ�6�J���W.���I�$8Ϸ��p���S{0�\��v���B�E}�ꚤ����f�E�j{To��w�V�n�
�q,��gwXY<�x��>˿.���r?�6���������~�%V���;hs?"�1/:|p9�wa�\�c�nj4eʿsun�v8WcH!̔���h-HS��A��K�Ng{�K������D�	����<䙱
�1� #*X��41v�q�Z1l�p?HJ�SL5��4��ee�`�u���2��Ep>���)l\��c:s�"_�O	W>�0�����Q�y�j��ݡ����ۂH�!�ǿ��,8��mh`�<��-��k�-��?����0K�_�;^��?���7�ƊZ�����Anon���iH<-B�O�<�����8�jF߫Na��u�Vb̜e2��Ic�j]�l�li���#�ᐷ%	�D�5��Ơ�G��@C}��s����c��-U���J�����	;�#I����%���A˃�;HM�#�t�HY�.�1�`P��`�#1�-��+�U�O��U���r~���t~S)�s���B�TU�&�q�e�n��8���.f%t
]����q�3��y�=�(�׸��{9��78�����)�����e"`ƫ�r��Z�I�W˗龍>W�;=k��V������{�?�3�Z�IE8	 t��&�N�2WU��L�ƙ7��8�
����\U�(3��a�5]��cQ7�������3��
Rd�P�u+��� �e����o���i�cZ�"�^E�p!����}�^�`�ƈ���%��7�ZL>ﻳ��U%�{-�60�7�v��B���~�˯xn>�o�͏��������W>ͫ�_����t��༽â1���
/���@=�o2�1���y_���;��PZ���SB�;Pu��YQ���BD����	�:�P�"F��]���� �^@�Gc�o�\CHm0�s4d�Lһ��T;X덼R{1_5P
&�8��yOU٨��9T���>������&��3�Sk�����ǳۃ��\�Ut��CJ�����h�=��%�Eͦ���{��P@XH��札�EЙO%��\òs�՜�9Ձ��,�YO/�Ϩ�����y�5�`��w`�x��#�٣��x̵H]K�y9��i�>�؍L8%�sc�WJUj�R[ꂙ�m'�K���@ ����������{A{�*�!i�H�7���qT1*d�hr�,�.��K�g�s!6�5t��u��:������^��+��)�\T��r����Cq�#�s����U*sƞ{�-<Nd��:�7�u��pIs�ݷF?���U�>���T�4�u����8����}�ߡ��7y�����_�"�=�Z��-۾�Vf^S�J�Q��}W�w�Me_r�^��f����A�P�q�VL�
�N�9K���J�d���kB��>DL��'u�4� `"��L���/Ky�D̃>�Y�O�DU��{�3��$�Ӽ�|�xʕ���|�㞋��|�!_^���
 �c)�����]���o1�r������ҸN�԰9��0O��ؽ�V0����>��J��)K�1��ִ�zJ��o��c��5��?���{�Λ�;������/rʹ`�a��a\���X���y�AH%���M�|������,�T�s
�S�L����0h�xڮτ]$���cLQ�UP����u5���#�Ӽ Să	\�mj�]�y۱0U��q�f0E1D7�(�V�{�)R���J�S)jZ���ڟ#�1��2�{ .�?��\�t�{�	S&��$�Øɍ�_9.�,���E��])r��SFh��r%lZ�{Ւ�~����_�m����6��������o8~��?� ��3��w��>������$�F�����������ŋ�UI짰aLb.<J]hu�v�1` �^=�)}�&�������p'��U��FxLLt�K�Ky]=Du���Ќ&�b���7�Ÿ޺PQ��nH�	X�2��X+tރ5P�u�-B̦�i��z�ӷѕ���)kP�V�^{��C�������U!����@��؊A�w x��B�4(t::�X!G�`a pu�UÂU�n�n���q�Ȍٕ��4�;�%����'�D�CC�q\�t��3��`�ZQ��-���l^�O�߬ꖇ~�X?����<�3?��^}�块0n��m;6��+��s�z��eA$M6DK�$��a�xB���ފ	����=���i7�%��!�P�v��{OS/ú{�h�15�o�k�7!�W�w�>H�F�}`�!���E�`%�!O8"���]Ϩ�N�"�WΫ<���6'���c���E"�.䵎
��Yo���<a����<���w�631N�C��Q3H�R*�6��'MKYr�r?#���r���Or���7I*�5;&��$H$��*�e�6�/�dE��*�#�mbQ���� a�}�$�`L�`L��Tf7�o	;��8S�6O�W쇖�w�k���ݲ���7���]x-�[r�}<s���/��2�}6�|����t�����W�n��Vغ�S����v�8*�t�5{f�f��*��y>���u-q��ĖlE� ��Dla��X��x7�&&�EUp�!4�c�����wx���,��Bwb(m�eAM�P�h1Fp���U�.5�Y}e�5����˨F���Ӑ�Q7�epl�F�{�;,�ѡ&�,��n@�<Ѹ����T�x�L@�RI���1����	�I%Y���j�h&v �;p9��d�wRx����`�YJN�X h�L��,��h@�F &�n�]�<��!�?�k������O���������z�o���e�����U��jj6g��Y:; ��Ũ�!��Hj�uѱd�2HbD$-#&������Z�DN3�uUUh��c&6UE4؞(�s}�0� ���n:�%��wO��l
�4���9FxKsHi�+[d��H*�����A�%�����Z��F�ʎT-vG�8���kc��MIk3��iӒ)���x������13ل L�zO4Y��r��E����j��g/��R��3'���uQ���@�q�1����^pڞ��p|�����`[-x�yϏ���ͣ��>�u�~��|���Ej;E�S�����1*s5�+&�3fpsj{n9�u�Č� 3��3�Π�udx�;kb}l�y�п�aI�������F[���!��XCek:ߓH[�~`�ƽ�k*��-�.2��p��r<1`N�0c�5!%F�c�$|�k�0J�8���%���_� ��O���k��'s�q��h@Dڊ�&� �lD$p@R4 c*'+i� �e�M�T�s�JT� hr�a�O�q��"�G%\���B��bn��w>�{l��7~���9�����}�����6p�>����,�X�|�R���b�<�EȰ܏�� ��S京V+�6F�
��jL���Ce��e�fr�H��1��ЖI֯��[E5)>���8ܣyi��}��� Gy��ȈT;Ho,a���⟁��@���h��%J����HY�֡l{�g8�r&/�<ER�tn%1*cL��dA!"��XG�p�H�H��U(���vb$�S2��u�Ӧ P�Y�_����yi�r[����9�$��+ǹ��[���XXC�r���]�y�)�����_�������֟������Q3D�L����iТ�P�@'Z��'E|Dv�J^�=8��,	}eK8~f4�ao�T�=���xZ�l}�`��Ӻ(�S����_b�����1�#;��F�/�z*�B�h���r�tP���ǅ��~���8ab�3הĆ,�H5���M*����p'���>�$a��l�c܎2F�%1%3(8�T�+�<_)���6�Hh���3��8@�B��}N��/���s}u������'��~�w�u��Η����Q5]�2����9F�>����R�t.;pÚ�$D�s�����{��PD���YH�)�]@����TU���{�z��a�X)��H�4��pц�	uJ[���]�G�L4g�PGX�8��̉Et+e���1��@�t���}��OsL�� ��U�XI�3C���<�b�e��y�3�׋$�g|�D�*jL�(��Ӿ>��=��G�'����}�ߢ�5+��TF�Wny�{�<��_���������c�?��4�}��t~�/0�%��u�,�x_Ϭ�x�cb��??����{��}	��f��0��`�(�l��w<���3\	ހ�kV�����{P#�~X�rCܨ�xq��`Zɉ�ʾ��iu!�ꮺd
H���09WA��%� �17֛��~43���y�[Q��z6r�AU3�Pp�g�A�:BV�����@��",�0�M���b?	[��h�N�v��x׳8?a��/���'>��Oq�����{��y����9Xe�8(�!��K��j��)��O�V%�8ܳJ�!�M��d5I��1x�[[g�/�*���7��E$d�S���$���(�����Ex�hy2L��⤾�J�e=�x�l�ӕZ��$��a-�}�g�s�	���H+��60<�ޙ�%&8�ӧ9G!i�,K�!�\G�1�;�31>��"&a�Q�̧�"R�!:���t��yI���2����3C<S��,���b슃�!��k�q\?Z��ٚ�ۆ���~����}lo��͟s�g��~�7npG,�M��(��\U#��d�x}�Qk��X��4�cN�Q���"������h�C�ݐ$-�1�����B$i�О�I{"��Hwʱ��sO��n7؅�2!a[ym1�B)�dm�N}R��$�n�/��fU\����:�0�Ĕ��$�1�^2�R!8��e��R�ÐuN�4�}y�'���d";aZ(>/i1튠�D<�%�b����&��e�RT������r��)���VG\���տ嫿��jX<����c�g��p�䌓�'��6G�P�h�Urh�QA�݃����K^�bMEB��� &8��,>���Q�:#!�Lb	[�ǉ�.��a���]�"^�F�LFC�wG�,�Fs*��|UW"���?��6���az9�$�}��D�$� �����	�Y���=#ۂhz�؎E��EPu����e-�l;��@ć��hqWzsQ2<�=}��T/Ս�j�+�<S $�49�;�fH'i�˾(`r�����^~ibH�R�U��g_V��W�]��v��c6�J6���j�x�9���?͓��;���o��]����s�g��3��{8�,�ֱ�1�)#��%�g�6�.F&M%i8�E}	׌׼�?Wa��p\�h�.��'�p������9�!�M��{��u�n��uK#����^D�cب��]��<!� c);D����_D��x���� S��$}����9��|����u���@t�$���w�aHm��1ZJۅe2��Jip'ֽy
ɜ1�O�׋d����IkC�$�ko��{_�W�I�W���Bp��i8h!{�d�Ip[|�s|��]S7Bc��_����`��7��<�V�g���>ck�    IDAT/�5F�/-�n�S�����m�I^�s&D3g%�nl�:�S��2�1�K�;����>�˵2x'ٺ?�f`S-Cpg�9�>x 2�딬��2�#��U�!]SU!�}��L��>���.B�sO	��|7�8�i;��,���=Аo{@uG�7ݣ�8�Ü&-�U�Z�%�q�	n�.JeR�r\2�d�!��S��Ma,I����� Wc�,����2�0�!y��rY�A$����a�D���X�Vll��~��x�/�:�?��T�
'������}�y�=��.��>�1��p������0��2�\�qDѼ�����~�C����ٷ�L]Y/=3]��m�Ʃ�:v�mx���a�~ֲ�I�P�!�ee@m ��4s�$�����������`���M7Hdl6z^B]��$JA��_��#��8!��I&,yb�U��ݻ�ys�XZ�kVm�����>2�탇@b��L��d'}"J�hӽl�qg����.R��&�=Y�{�E���6�&g�S����?�מS5X��>����O��?򛬞z?���G0�wy������?�鰦�����8�����]�i�=ڏ،	�àE�Ap��A��,����~�;SE�r�w!>���n�
��ҵ��	��p^�b�kf�2�j�C�'"]Fm]K}	�&��D:39�a��8�W^��8ϯ0t���q�)A�H��S@%�Ü���7&��B�2B���a&lBv�ˆ���WÌ���@
]-�1MK�&�aq���b�\Bb�rJk[M)���1��ރdҚ��Z�}(��^-��Ld�i�}�~a�����g�w9\\g���l�9|����_�(��ѧ�6l��M���ǰ�?Gs|�f��y��k*w��ah��=����9d��`2��v��@�C;��4�}�^I!��i���8	C:-��t-���g�b���=8�:	�͘:�k8�s�����F-J��*�D��Ўb������wo���P��H9�K�ݻ��lԄX�F1V2�mn�γ�m�ǐ��bQ�h*�sTbq8A��m�5���l���m�t��/�eTpbS+!L�B�-Hv���!1ь1X#��% $ӹ�S:����� +a.a�>��W���F*��V���v��xjS�cD6���h�� H�ƙ&�撮3��`+Bc,���W�,V�W��u^}��\��?��#o�`q��O��ݻ��0�@���(D�:M��T⁕����^�Pn� }æ*oi��-A�'W5����zb�f��(�(]��z�a-�[�]�(�N�#5�WʶQ��c����x�be8���9b�l0&��[�^�M��pC��>l9�kV����c�ZX��sf۳4�5�C�P���iX��n���9R��r�*��56͂%5�v�M,����X�JX�p��͊fU��
Z��v=R�cB���`�ϬK�<�p�5�n����	o��mUQu=X����p���s�X�ΖK�s��ؚ�R0-U��9DW5��Z��{*+4�%�z�b�IWs�����~��Vh�s$'�Jue	a2<ueY-WتAհX�jO�<�zU��RA+��9��1l���5�1>h~ꊪW���������h�����+6�F�	�l���uSCݳ\W�n9fA�j��a�t�:V�`t��M��U��Yha�Z=Gt��Ji�%eƻg�\������]R@߰��ط��7���>����~����W^��ѻ�쒍��K��V�OS�s� $�Ӏ1j.��G���ꕘb�[�*��h$%��h��52������$͐,svӕS��.���S�����~XմW1�����RWUp}#]���g�d��x�3�P7uTH
IN����Z��ưXԘ�>&�lUщP�#n�9�l��7���~��l}Ge�֡��"LjX��`��!�w5�+T�����{���,GS�@���ı����Ud���q�d�d�������>16��`��e��KbV��9��Ɖ	W�QY�c�^==u�1Te�,������5̭S���;��C}�1��-�z����x<�	�"<ſ1Ґz��V�/y�+_�?�#�ڻ��#��6n��;��?�w�p7:�e0IyD�+�@���� i/�>�j�jY���;�Y��n��Ε���ؚ�X���Sy���=m�UŁ�<\��D�����,eɲ����j�Z�-���%��hwF�eU{��c�;A]ͪ�0����nt��ܲ�r�����ۭ�ME��8����y8ߞpj�öae`����ᴷ���-���u���W��5V��h�QiCMOc�2xo�\�����!�}��>K���a�*�Kܨ��p`�ҩam�"��>�u-'�1�lg�[0��hI'k��n����%�kײ�k{�v�ϕ�o��5�m@�yǶ�,�q�(��5��5� V,�3H︹�u�]�SYZ��{�m,�k�����Y�#���Vjx�∗��4昅Z �5h���[�Z�����F�|vJG�rQ��5��S/�^��]��dK}t���ܵ��-���im�����^a��4��ǫ�]��]r}���d�[��L�8"/")�^���o`���y����W>��_���Ӹ�3����.��v��U�����x!$�
�[)	4�.$�s4ĩ �z76����}�:���ޒ�%�BP�x�w��˵��a��ϟ��"���$-UX��=\<ܸ[70.�YJ�)��4�r����x!Ŝ���ʚ7�ʘ�o�&7>�f.�H�Ub�Lpw*��U���}��.'����
��hc�u0d�V�F����{�`��	i�+{ONY���!�T��f�́3�!R�x�s-�kH�P[�áV,���gk�]�w����r�_E�-�m�����/5�(�v��L4'!T�"��B�T�">������;�I�ӗ��cO���O��wZ��2�}�#�đ��e&�D^#�~�(��0�c��%��oў�bũּb8x��x�mo�t�@*۠F�^�l���D������w��q=�ز>?�z�kܹ�u�x�[X_���4,���9��1�[��s�Vv��n8��*/~�<�[���۫9x���������5���7�������z�5��q�{���醍}y�}lzS��9�����1�ca�;��՛���78p-5-�Y�eQPcYw-���=B�p��94H��ځW,��pG��+�׾w�#A����:D{N��m96K���2Jמ�/<����c���L�7K�4R��^a�;|#��CNձm[����1g��;Os�6,�����؃���y}����b���Ab3�E}���ZT��k���RK�,t����+7_B���uH��.N8ඩ�����Mc-��;���t�7ի��b���P�H�"EY��%Q��m�������4�'�A# @�!H�Hw�N�A���nKjI�LK�hJ4%��H�S��*�����g�C>�s����`��](T���=��q��_k��2��(u̦�бbl M!�5��
�X@o���fbbY��D�$����c3IiI%(�$�BoP��*!���2�s"�+j�p	&pZ�&��,L�:�fv�O;K]{�^����*7wn�,��2���:���H���R�%�>�p�]��~W�SzW|��@� kC��20�� �i
AESKλk�]�ѷ��4S��3g� �Y1efl���_{��V�O�J�Q�ڍ�0�х��ߌ|m������u�H0��Z&��2�cϼ�5�h��0up�K)�y����x��w�kv�Έk��D��;�VS+v�w����;M`Ή_#��pԮ����~JD��=����=��`�>Ό��o�� �$*�x��������ϱUt{K\w�A6Μ�tC�1u]S��%��Qĸ�P���)�T�N�ŷ��f[!�.h~�{�a�`�����I��Ïk���z�cu֯�ΛgW��R!Z�`����m�?�'K\޸"��K�N��7���?��=�(y�a��HMhc#������[_�2k��DW:QJm�(�>�N�Q��!"bc|H���cp��TU�t:	~W[1�\����'(��{�i����laT�z�M�E���I�ׯ���CF��s��*���>>�qY��N�[�5N�FȄ�F_�fo�&� �C��/���kF����H�KR��v�i�M�\��͂̀����x����f�����ӿʡ� ���Ғ����'R1�ڌ)�x��o|����c�V���i��S.����x�/|���E
�1>���$J��ls���;�#_}�Ū���!�~������:�:�K��DR	�f�Y �C���&}v���#��?���G��E�d$bv72�C���^d⸜�sR�ڢ*��$�x����.;O~�~�}��܀��u��3���C�"��q1"����0�*��|���c���;2)�Up�g����k��=�+g�w{l�����o��*v6�p�[��z[a�2NȽ���C|�4.��n�	'��<�hs�Z��L�q)5�'Q��[���a��p��^�3���������Dƈ���{��Μ���7̎񬜀Y�5�*xw�j�+%�{�l�k���4�+��P�K��$�g?Ecjه��Zh���勣u�{�ՊfJ��O�fQ��bߕ~7�A�B�����gS�*�N��8����x�Q��|�3��Z�UN|�2�z&�����$��*�)�R��"
�]1�*6R�Q�#8���^��|6��+"2����pPW�`��ą�
z�H]�,Im}��q�����p��+vg�@���X��N�,���ef�d���1xy[{}�ͮ��$�;8YS����x��?�yW�5^'�
Q�A&
�C�D��� ׽�!�Q�JJ~�%u�\��ja��?p=khƅ%�%F�ʠ��jHE�(�X��-�R:)���>����#�n8Fv�0�Ê����\�Hz䱥s"������6�{�Dy朤�I��ㆇ��]���1y^��
c!�
g�=���^���2'�p�+_`��ߥgs�q�.��#l�g���m�R4�m�	�ep��[Np�#�p� >�D2y�	����Ș�X�Z�;��'0x�����g>MH1�UI�S��"ѩ���ٿ��nEEem��!�8'�"8�?4Ǹ����3��WC�$ê�[o���c<#�BJMY�(�㰯�N�}N��E֎�]A�����w��r��c;l����Ǹ���7&�K��U%���0�`L�򉣼�ɸ��UTT��!�"K���P-�ʭ�7}���>�wd�^Rk�cޢ���|��D�ʋ������kꆦ~���=�װ�g����w{��qJ)k��q��?�}FyNT�)�}
<�� t� �Q$J�A��N�-�m{>7�y�}������:^@YW�ŸHN��{,�	��ڴ�QM����प�-�5�=��'��v,��&�t��&��Ț�<��̃��!��0I�k�{)v�om$�.׶��zw[pgLedP�B�]����֢����F��Ch3;�{��6 ,t��6����n�{%_DS�Ux�-�}�VTZG�C�D �i}�Ak���!�8|���0��Ek7��_I�q�Қ8�"�����	r!)�y�F��n���K�:���[�*A�5�nn"FC�͑� 
�/�*�a9�I�l�<m���3�c�37J��B�&�nq��;6�t����6X�&�sF�
h��	��,��.�(2�vDEA�i��C.JֶΓF��D�vl*�T�Ex�7�s�����o}��� Q�Z�2E]�II'r�D`,H�}�H����`�F�2��u����=�o�QU���{�-�(����NY�՞�j_���&!���������|��8a�6I�"�',�c���Lmu��p�}��y�9���̓�fD�xr��p�Ϧ������f���H������Z��w9��{P��2Z�O0u>F�sh,��K���*��9p��M�y#�C.��W�a���c��{��}��%�O?H�6Q¡]�9A�0��K���gy��Q��ɛ?�=	���ۗ�"���(��gkjk�Jb�b0�FF[Fr�(��MEu�2�zIԃ�B�ս��}s�я�0����5�|�*�ͺ`^8��D�d�n���~�����M߯���VY��s��؇>�(��p��IT���S�WQ1`���s
��X����0m�u4��'.��❵��so��W�̞ɻ-����B��VlW;8�Ȥ#��$�^�mk��B��E�5�ub��8��
B�]���*GK��!5R*L��N%�J⥢vm��m�Ԡ����W�k������i��FnL�E���^4��Z�p?!?=+����*���7G�>����AŅ�PbZ��
�%X����f}+�'ӈii:gޚ&[Ρۜr�8����e�߽1������b��(왠�����o�����vMJ�𔻆q-�������mNm��Ds�B�e[��UDl����B��	���$>����Q+M�����qz��@���yh��<?���ꁋ�x���n���m�y�\^~��~zx�ҽ�s�(�|�-�5tY0N�Al��F�zG��	��͆),��,Y�k�V�Dc�
aj��ﳝ�_Tx�!9�t���V�l��MOl�f�A�TM]r_��jd%(rO^Y�QD�笾�"��U���e
+Cuĥ����C�<�!t*x��ˬ�?��3*o)��C[��W_��VQ�A	u���:�	�4�	����x�'�'ۋ��2���G�� 9L��]�C��3o�.��.6x��Op���sHjb�+��	TW!㄂�$��B��Hm�C ��$ғJ�Sv���ء��=�C*A1�d畿"�=ZƌG�Xﭾ�'�/�6(E��Xs�����aEG�]%,�S_=OU�$cL�4��{⨇�}Lw�[`���k-Ϭ���|�]F��C�|����d��b<B��Q� �R�(Eu��ŧ��7�M^�c��1�ǲ�A�2d�I����+��5�X��سv�u��ŷX}�5E�ˈ��}��>��t����d[��f8"��Qol��.�2	�����g�m�^{�*��e�<��?�Q��<c3�WW�6Gŀ/)7s�A�C�=�	�a�(��~�����L���ݫP�M�5�d�@ʾ6�:����	���ڔH<����&MK��p�2��JBL��Y$���K,���U/pZ㥦�zX�0x�����U�DTXQ�S�I�RN�����!��M�e����d/Կk��w���Z��Y�D��Ѿm:�Ӭ.����ڹz�{I�I��+ŵȺ�~&,8���Fз�R��V�����~��｟5L2�l�4�h>T`ӳ�o�h���]�����y�P�I�o6�j3f𼈦ߝD���R�k�Z<�$9)�ux�I���>R�ǎ��������_��_�w`a��{���k/<q�ܱ���{�]��9�z����l^��^yyGhb�{�7���b�<8��,�j8&�R�^Ba,*NpڳQm�	EڅI�/���a�RzNhR���YT%�Gz�qV�&s�h��`����券~�7��CV�z�e�B���(�(�#7q�g#�-�,]�܁��1~���8��r���8�/?G�{T2�h^�qV0*+"�饚r��|���wYs{�ko�'����ĒHX9�o|��ͷ���ͩ�c,�m��@J���u��p��'x�����Aݍ)�C�1QY"���}������}��s�!�l����y:�K*��&�C�;pm�]��[r�6`40�5�DJ�S�Y:�.�~����d|�,㲠O����X/-Go���?��GU���8<��3�K��دr���b��Ć��广����`�A�6*�:x�?�҇?Ψ,�z�xj�ށ�������2�%k�<�O|�z����F8�8��)*O�;���V�ޤ�p��6��-SD	��[O��,ʄj�<�=�8��*c_')R�#7p��3w�9��    IDAT-X��n��ӏ~��j�+O~�V���>�'��o������\|���iw����D�����ЯS�s��>�ￗ�m���EV^}��z��a�Q!�V��sl����]��Rn��Y{:2�+�q5VY"初A�I*guM�B)�Xz
�g�n�6��F�Jj�P�!#�N��`�l0O�밝&ꤨ,	n�|D}�2ó�^��6�� �Fh PR�\(5�1�UlӴ��:�V��Kr���	����/.lo��j���(�n�9x$�3�yϖ���$��"�("M������0��}�P�F���*Ip}�х��@�2!����s�җ���2��X���
�
�x:A�'�O`I��+�Dh�)|���e�����t>�8��2��:�A{i�GޓE�p�E��!�^��`��dR�f��ܑ	���4�jiH�&6���A�(1Px�vo�?y�w�k�7��_z��g�]�Ж����y�{��_��9�/��<�u���%����ya�C�Do`\&FE�oH\[�FH� ���^ �.8�{�ڔG����D�����B��
hɅ&�Ա$qc�vh�b���[p��)�f;>�+=���(��k�x��t������(>�xK1ԁl���j�,�����1���kɒ�l�+(����c�I����.��=����Ě8��b�x��Iq��BTھ��61�\�x�9�`��M1rH���#�R8�0~���U�r@�Y��bl��l���-�Pq��~����u+��{P{�m��HK*��K�p�)��7x-�UD�;F�iɐ�؉Dr��:Cl��D��r����07�D24�H"��2Z�6oT�����c�,�����Y:�a(��ݎ��ȑ�<��װO=����U�XFf�x�5^��݋���c����Q�c�������E7�Hd�܏ @�1��̛��Wx-�츈����Л�p+��&Gň��P�Ⲓ�+t���&h�r��O���>Oq�:CK�KL/"�5��^&�2��__�:ra4�SG8�����:��ċ�n����O��W��W��әgd3�0GiA�D�>N8�鿇\:D968x�T�'�+��
10L2��S_�,)O[@e��@m�$j&���s��Y%@	5P�Ld�,6
е4T0��c�0�-$N�H)IRK�Dƞ"�� 9q��c�n�W�Rh��J��cI�Cm���
g���Z�m���D�C�`�YW��B�T�h���8��EC�>5P��r��t!���pg��O���97�G� �O�
���n}H����˓ �I��p^Zk��B�Y7�h
��8נ��f�y��28�I���2Ӥ������&AY��5�����.���	1j��럇k��م���sOk���:k=XQ����Qds�����,���r}o�DK�ǿ*r5�]6@S��M,�v\dS���5�*J�뚾����a^1\:�y�,=��׿���/�.��>p���7���:u���i��2���.�Ҋ��
�E��>��UÄ�;C��Y��l����h���͘M���>�w:���}� �exJ�q�RE9۱���%��8_C��1�5�(��*!���	E"�Y�Jx�zהzĎ��)\(�G�N@-��ak�����F��%㔠rM���T�B���MrX�F)�k�k����S!�'I"��C,KV�o����&Ne�DR��Qi(\�V(� ��x�<���!��k���QH��2�jKiǁ�I;�XP��->�S��Qe*_R8��%��6�^;�ҥ����Bj�h@�:�4"W�&W|�ʥ�,8K�&X��8�$Aynn����p�Gn;���E��UP���T:�p���C�+~�:Q��}'�O�H��l�1�h���/p�gоd!є�+!����^�!~�r�%^���3>�c�$,ت7���ƫ�нp��c'1�&� m��\D����/g�����/�VW���+c"�I�Bxr$g~�#��/0�����tek�>�j�;�a�Y��d���w�.�u��6������i��5h)ɄB��J�V�Qw'����9v׽���2��ҁ�I+�(�Έ�(�W�*Bw�ˊ;N�`�r��g~����T;ۘ|��F�*�R555ƙ@>$RJb����'�@���4�cԘ)^4nM��>c�V%���P�.���g?cy��9h]ծ���� �q+�ӝ	#�M6�>}���o���^~wP^{�O�w�@�禼ح@>��b�k����w�y���3ʡZ�!p47V;�V�����bB�[��Z;��H#p:�zd|dt�g>�ٝ<����ls�|�w^���88��'�ٮ�R�+OS����>���Jc���������v�l�P15w����;��8�>���-V`���#+Rt���NPUa�rS��A�kЊb��v�,����K]j���
�G{��@E�-�IL��S�*K���נ������iD�IZ��K�1"�@G8�B]
g��!tH����	9�Ьc�k�B���)A]���U5��X+QB�ʊJ�8'������	JR�{��eC
��!������1���&ւ�[���i��-t�s�<���S�Z"�#��)�%�HQ;(�B�y�\�]�9�::�>U�J5�F:�T0Ϋ��e.%��O���������"0VP��\���[ly��o�s�C�|�]t���A�WT���/x���%����^SJ23�/�K��2f�C���r���FY`F���i��:K4Ũ��3��'�-e�#L���}��g����
�F��$I3Jla�D�	k#�w�T%h����:1qՊZfO��6�7�k���ٽ������0{އ��=�=EY2?�ǌ��ܐf��s�&n�;?��ݏ�@GԖ�J���I/U�����P )0o(n�������P����Ս��yš��s��g�y�������%�=�?~�= ���	ʉ��Z^*�����3�wءH?%���Y����ݲrw0�ޙ�[S7����6�R+���I�����؏��7ȫ������o�o�}�]�;i���3S��ɳ<���y�3�P®���%�g;;���]���jj�ZZk��i�_��Mn��^5�J�W�V����u�Y�����_��Ǣ�'����7h���/>�ԗ����痾v�I�z�p$�.���F%]�Nǹ(&�3s4+�w�kyD#����^�]��u}���(S��;��.h��$�Z��qc���A� <���q'�w`	!#��Exo�h�1y��)Q�ol�\J,3t�֠�ǚc=^(��H�R��Ho���?�r�<�uh��P����0���1&�F�OjԶƋո3�s!�Ӂ��<���@���e�qΰ�l�yTةKMF/�4��T� ИXQ����u!��ܒT���������Hg�EbqJ3�5��Ա
T˽���l��}I�ua���ْ���,um��멊-����yK�<�THd�Pc˂�˂�/��|,-3�_��9j�p;ی�#�	�I�o��;��GJ���wp���		���٤�a\�E��j�Q�uO`G�s�d�{�����UE�r�MD�4�8Al��-R7�@4O�-ua�H���*��d�q�����øNL_D�5Cj���U��N���vϼ��v��ݛ�vM{��<�9���&�Qd���PBS�)ä�ܽq��f�����r������&����5G�����0������ϭ^8�*�d7}ⳬ>�4W��s˒|���!����M�΀T�0+��*4�8� �B���~��\য়��
-u��f�'�;��s&�ج���ό��Ϛ��@��zv�g�m��x���}��,�Y=��(!�M_���޵�E��mA/v[����g�L4��k0|G)��x�0��`����8��>���m��g��/����� ���]����gs�Oax���a4�v&�"dTx��;�m�	�)`�E�]�q�����I��eEl�I��KO�
UaM�1��� ��8f����c�D�S
_C�!�Z)��p�蟺����o!�b�D����G�y�n"�s1�&$u�t�(Q�IaJFC���C,#�PTΒ�Px�����(5�;���U=9d�u-��vA�IS��0����v!%��Lx���/#��4�1�����t�]�NF���T�1O:�Q����g��c�˗Ht�lP1��Җ���C'�v�25�8&��T���{2��;dYOb�q7C��;�ֹ&.FQ��xgɲ�K�m��DQ���x�stJ�]�B�:�R�B��UW��8�������\9�㍯�#rL'M�G]�!�H��VH�pnH/��E\e$�>ȡO|���e|5$�^�����^��%��^��EĚ�ڣ{	�h��vd�yVkϰ�����ȣ�:|����oS��:��D���2~s|�%�{�w�����O�ҙ�K�n�H� ��ȗ������3�Bt��z��_�h����O�����S�S�o�����������rgtSqDV#�9Ҍ��,�69��y?);u���݆;���g��U&H�>s���-ں:'�o/����%��>�?�l��771l[��2�:�v�5{�nu�r��������'Z8{�����fj���Z5��R�-8�H&��5�V3�{:Ғ�~�d��neÅr)���|�	p��kv�[+T⨬%
*Eq�-������]��5��Shw��o|����_~��-���C7�&��&�ϾET���m�ۄ}i��g��
�IQ���B�0���B���g����ۭ*��q���ct�E�� d��5^�֒��xz�o$,P�%I"P��kF��b8d`,y�I���GV�kI.-uO�[y�gƗ��Qc]�1�k��0փ�����-<I��(B�	~���zh��D)�0!��;��O�;Z׏RD�F��a�)"�e	P���ﳘ�������:M�����B�qs�������
]�xы����W������EɆˉ�<���(�>C1��,�y��?Wvj�Ń\w�.z�%�('K"��#���
/b����C�a��B��2����ZT��4�K��b���xL��EDUz�H�1l����s�bH9�$����7���~��.s7��"W_z���e��P��4�f]L=�����r�N8��ǹ����u=�:'���ݯ��7���9O�#(�%�(��Ұ������X+,��9���9|�#�� �&���l=�4��K��&��l��z�&kM�λ���T�m����v��j15�hҐ\ңH���an��_E>���.$����r�҄��d}���Ο�=�x��� [?2�����{���E��)|D+EgϤIܙ�e6&mj�5qC�us�?fR�)���n��G��{�I)h?k�O��� �%��G���~����a��ҳ�Z�g�t��}�V��T�}}�3����T�6���I��:�M͞��z���x����Z&����_��ƑjrO����0���P�3��Q���|v˃�tߗ�)���?���k��]>6�4���_}������������W���ZrhHY�U3es�{���\ٌ�P��gK;�9F/��o`��Xi�ӘHgx�Gw������,-3o��c��V��G^�1�),i*B���t��5z'��SvjG�-Bi��$�кg��`��j��!=�0'�c�^�Sz�P!��[�U��6��9���=�dQ����x�����I�A���Y��Y$�nbX\��*���;���Yl���*����KK1�Ȣ����K.�1��P� �5&/0u���UʲCZ��I 9��G���r��>�\�c8ޡ�=Dl���OFY
��'��8)��@Z�/U�o)|^�P��Ұ�T+\G����>Xe�-ҭ-��K���6��;\����8~�}���A����<*������*�i/�Q�T�^w��Q��q����,w��/]�L�_�����3Oq��_Ü;�@�P]QF��%i�DIY��q�S�T��Y��C���ǘ?p�am��o=Ε'������<i������}����"��f�����gsأ{����I��R]��7}�Q�O�����d����?�����J����a_N�����{�Px� C[���4��������!=��Z�bZ=�5z�qy;3�{�a�C4��{]#{��:5X]k47���L���1�UK�낛aVF[�;��u�K�xS.�Y~7|>[;{V�ٻX�����T)\H�l��[�b��3A[ja��-��=�w��~:�B7RN�&���uj7��~6� �����Y�7�L������ãk^����������o�\������N?���5d~!(IM?�Z��s��nv3OZH��M��6+��ܧm�tP�^2T�r�ހ�`��[Kt�vn��_��{��1��C!���f��>� ��2ok��*g����D4�O2��t#I\��r�5���Jjj��PW/�/�����"bOeJ�%�#b�%*
E��ň��b{�^8�u�c�,u]���5��M�tzX�0u�s�uDK*#A(�.p��v`�F	��Zg���s��_�w��	�զR�J�	Ѹb[<��e��-6�/���k��1#�#|m{�YZ$���S�!�9:�uQ ����N}�ȃ��\�X\��ͧY}�UD1��;(��c���x��g�J�D	�IJ�SY��Q�)d�p%Bd(k��a��Y{�u�:�B1�:{�}���n�
����ddQ��<���'������Qɼ�0�1,���oRc�^:@%1ۣm6��������K�a3��V�p0��y�_e�ų]\@����1*�7"b�puNg!acT���}��,}��~�B:��e�>�4���'ī��&	�C>*���2�j���������b�O��F��8'�`yc�x�i�=�Q��'�����/����я�����z����lQ���z��o�8�U��5��N��ک���nJ�lyԩ�4��w�71#�f��k�M���\��ȵ����-��V)a"ӌ��f@׵��fpX�5T�5��R�-�I�5q�>����.����Hi*g0��GH���kZ�M�>E����d�l�� �P�Ϛp��P�^8�JD�Xbl� .�Q
τܺ���D �Lh[k݇Xt��BXGVzw�b��;^;y����;-ԟV����������D�����'o�|mĠb1�Q�*��X"�x�"��Ƀ��cm(�j��i�`~@���mn�Cy�=y��֢&m��Z��� BR�(���
I�$��|�1�N��qX%�]I��PY���ۺę�>�����@���d^0:º!���������sxS"�N�������.NH��@%)�s�d �mR_�T���*�ga~�$������@^s��Ӽt�y�F��I��!I�G9�]�5[$��ʠ��.GzO.2�0�$���A��J\���k6�}�\�����\���C�^���%��4B�R��q<���B2��dkc��A�$[�zI�j�z���R�T!S��1^[|
�Ze���7W��E.��<K�;"��(};,�D-0:fю�-
�U=�ј�#(E�r)5�m�A�Im���0z�/ImF������v�,�e�/����Av8{���:���;ԑ���H*�a]D>V��z��>��|�n�(f�M�7���7x�L�\�ʷ�;a.��1�5�9�����Sγ�?��G?���}��G�9IU��	.}��a�z�O�S�xH�<&v"��=H%&��{]�{�Ť�;�w3��ɇ8�aH�&�w��GA�e;l-�ħ>�����I�����m�?�����?�����#��K���ӵ9 jCE��"�U��^�Z+^H�$�ڄ�+���u�*d�D�FK@8T�v�	.�^�0���hr*��q������UѸ]m� ?�kk��k�/�� ��9�B�d`tRP[A�z�B�X[�g;��Z�i���mΟ�lv�\�sh�n���)�a%� �V� L	�F�p���U�)���H��f�}nۗY��Z�]������ dl�(�    IDAT	DM���<e��t���-���&�p�����wΜ?�/��Bv�f.\z�2%lV���M��݀T@U���s��q��W�8c�J�ܟ��=���{���-�h�����C.Ɛ�V�c�#�1�Pĕ#
���l�s�����7������i\� D�Ě���FY��R�xo�bM�DaC9�s����t -N�5%U=&r@)�F	�l��1Z	Mm,��"��
�JP�5��&����Q�cz�Pz��(�QQ����Oe�87t"��3vʊ�:z���ի��
΁��(߶|�Ra�A��H+bl`�Z��%N�P�R�F��A��M���t�=~kL6��s�O��S�rjp����$Io��xH?��>��O���S��Rrk�ӖaY���J�[E	[���غDT��bЉA�3.$���D�)W�u�1�Qwҥ9��q1BǊL��!���J��êd-�r��p��?� �6C���������_G^�H�k�RG�I_����.����e�u�m���C�p�c?�YX 3�Snr��g�x�Y�+c�J�
��	��5�H)������c��'��qBG	޺#!p:N�>7�u����?�t���/���n��_�헾���N���.��2��y|Y`#HT06�1X��E�hH�0��NeU++�u5O���Qq�%V��~�i��J����?3�@���ֆ��& 1��� �i�0!�Y�oc��[G�쳿�Z��>D\+�m"'����S	C&<��D�����d�Ƅ�����Rre�f�vM���S�_����]�@5�X��9�=t���$xoז����7׭�G����<J%eS�$�P�O��,�����B4�G���2/���"h�3a,���a��}�_K)0��,HϒsD�,Q�(a>I)kC^ٺ|���7x��_c��š8�(
6\�w�'I�T#|��s�/���69֕X[bMEm��҈@K8�b���D#���K�;7�z3o>N�E9E�Jh_������*(F�rH�0�DD�$R$�#\�����`$Zh��"FTW�L3�
(RT��)ǂr�iÜ��IK_V��Q3H#z���Qt��!�I��D
�(B��"�8"��,�פJ`�JJ�$c�����?����*����{�'˲�����{ofV��U����<�@X�(��$H�p�V(�Ѓ�:���)��� ;l:a���IE�4� @=��檬��t���9��{3�Ѐ1pGdU�ΰ�>k��Z�B�>'�قi�1.�[}x@�c�(��s�-��ak4"9�q���L�h� ���3�s�����P��9~:����w��Rmm2�aIbp,J=����:�l�N�;1Vgy�/�'>�>�OQ�,n~��o~��>�G�o���f�b"�aXVl�)v`�p0���������*͹Ӡ���>�'�ē���_d�u��7e��j�d4ap��p�C=���ˑ�w����!*K�x�1Y��D�9s����sW��_��"��[?�!"z�Ƶ>:y����y��HN�f��֪�׽�7jrQД�����2IU�d��q�Ǻ�ۻ�;~����`��׌q9� f�δ�B�걘�~\hk~cTD�B8Ǵa���nW/p=&q\��o=Y1�oyZ���\�W1F�	Jq���sg8q�En>}�y�!�bqEy�:�stc�����fu���r���.-��k��z��y��ߺ�ȍcW�4y�/����>������ȣl�� ��&Ng�&��Y�V7^�@�1"�,��SK[��H̺A�ʱ���F��e.u��7qs�%v�t����P[�z-��nf[�nL�ٝ�@Y�dN3�18Q�g>o��o�lN3�P�m2QI�1��kL��@�H�P�j(p3��ll�:E���A�0s�P
��=C�P�#�(����d#L�h��B�F�8 hA�P�%���8�s����-s@�X�QS��a�$�&®�!�� �I�`f���d ���=�<�դ�Uӭ���Q���Mīgow�kWw���ޭ���}��@ʬ6ݐ��TpE��1ej(R¥@"76�m���G����Q+��g���c��lp���};���N�8q��_b�C��3��S�����~�����!R�aC#-��*�U��Mٳ������ϛ?�_s{� �;TE`�ɯq��>N��������/W���4�5`�69`����(���/b8�,rf���c_��O}���K�)�����sbʝ"�Xc#$t�����)�&v�r�uC§�M9!5i.y��	�>�:�=��"��^���Ƈ���w�����{��>�!4S�	P7q�^F�\��^4��"��[���_de�A���x�t�?>\�C"w2 �Y�}�AY9�bd��L�n��P{��Gc"�e-��E����0��X��zLq?�X��E��Y�p#���P�ΕT�����ð��a��q��9�l�*����<۝�o��rH�u����O�f��ӯz�o��+�?�ȣ/<@�}
?�Ŧ�9;~�E(���Z�wq�L�%)�1O>��6!��3���]W����O�>�����c{P�'���g�����0��0��y��>�3�K_�"����J1E~�c"�^$+��	�j�XJ됶�fJ��/�(�F�뚦�����Fe�{]03����#�H��=^������u�F�L��k���Q�E� o :�|�^���#
��'K��ԓL�u���0�H��4wc��Hʔ)��
��5�j�)`��$,^{�'���/]�054��^��_`8:��<p������������N�������c��B��f"z�[�������]Fi�a�a_K���x�#����]�3#��9��t�roN�yo���1z�[)f�u�"��[�}�ٸ�2%�a�S\�|�~�9��+�&�fʼ�RĄ��i��Ʌ����#��6���6W��&�|�/�>�<�!��2�{
�j���p;L`:e�m�7-�;u���A��L<eI:�����7���>���/q�ڤlQO�fbq!`b``�:��	;FƮ�����ݸ��t��k|��q�gK��'�M��鷾��r��?���)�{��`�O��/�/^|�^=&�M�hH�갮<����w$�s!�����so��,b�ʲ��r��=�酣�q�+�f �܍�H�k[�n,��m3bBS��qݤX+���;�3_����h��
���#�Gb�6���:DT���k���'N�g��34��$�YZFK���I��h�A���~B5Ǻu8�^���y�|�2~ۻ���ט��f��Y'�R_}�2�EH��#�U�%ѳ�������!�n�u�]b�r�
�;m�nXkIQ�Ƒ���ւ�M�2�ؚቂ�����>�<T2z���M6_�F��q`��d�bʲ�,*�"�b�ÉA���R����di�� <Oe�����l��Q���؛�*���x�[o�co�*���8�a��L�k
������	�-6)N]���N:��M�J!JC"F���u�{�[�N�.�]���0q��_1/Y�/�^�ۆ��uI���R�B.y�~z����QPF�R;W��dTV�n>��OͰ�q�]�@<}���S\|���8��gnq0S�HڻN��"�>�M���6��ޯs�����ÚL$�9�
|�x���s�bNr5?�63L}H���h\|����2�6�KO�D���ࣧ�x����{��8�"q~���V�mþ��zy��w�<o��s����c�mq�ɧx�Ͽ���+Xw�m�:��0��D݄�N�x�,78�mFox~�#����	2�r�{O������.'��xqFj�������35�Dhj|�qDa�?;�L��g^N\�N�n��WUQ�> �Ór���e��7���~BC�ѿ6g��?��b��%anr΍�)l�r��Y$w#��w�{��tBv軚�eE���?��]��kk�0.8ꤾ�!��g�Q�F��	�Rn�p*�I\ѹɥ��~r�x��1����U������/~��Nwm''RV��>6Xg�U��t���M�xnJ�:��DX�r7�q�/���\�Σ_��W���| �r�U�P�N<�V�'<N����S�_���%Μ��jk�5b"�V�c�q�G��Ү��0�ƴ���G���k��U������:�,E��(;��u4)�S������g��op)Լ��=^���&����_�\g�>���f�H��4s|�	�S!`L�{\G��a�f��8�	%ab"�q߇~����n&���i�"���� ���m����K𿣗/Ѩg>�2<3d4���i�����7���.�y����/a�
h	�D�֞Ѹ������?�v)4)cA�mt0+1�e��8z,�HȈ��_|�4$��fFJg�h�rɘ�Jy�d��K���?��~��x?��!��#�f�g��O��)�s��>�i^}����no1|�kx��{c��R�B�#Tۜ{�u�a$��������T�]4����Ë'a�<l�����[O�cvs1�̌� g��^�����-��un?�u6�����~�x��|���g��P#�a���I��}���n����V-ÊI3fs�p��/0���p�?g^�f�m����c�}�C���&:���x୿ �����L��$�P�e���~�34���8��Zn�)�;����^.�r��.����jPDL[Y�m�.\x�շ�����~��&|���[����x��.���X �iI��Q���js�Z��8�[�xT�[C�G����\꘻����y5e���v��퓘�4sO�Z�A_w���1f�������භm�^�W]gZM������!"I�N�g��fED� ?9dv0Ξ&K�h3�����	�n%�o�UR�NѯS����E�@��3<@���V?��Oye��v�]�c)���0&A�5��W��֕�"#Ar2�S�;�i�䨫���o+���M��$0��w������P)Xd)av���s�Y�5/}�	����[~��z�;��l�j���s��e�<Ʀ�~%`LKKi�B�)E���W!y|6��"�'8��7r�=`�US��g20��	��Q]|���܀i
�pHAI����NΦ�Aɬt̊��y�a��2O��b(�PK <���4/�٧��>K1�6���,���Qѥ��YՃa���l�D"HB�!i�H����QZ%b	M�$�I�O�(��$��Ol�5� z��	��3ݿI��g(�.�KL�-�����a������ބ��
��M��&en��}n�k<���p%a6�ɿ��cx�����#���|�k8�����)����4"���:�ť/��~��y��!ψ�8u�w��>� ;�):��s6OX^#�g���ҰI	�mo�*����S|���w�iN��^�������f��-��9BI�9y�g.��j�0	3<#`R��c���O|�8�pj�uOѯ����A������9�����\	�Ery��`�����O��G����������'���?d�>�]�@�.pa!康da����1�]>^Z{}�(�����.�V�uq�ŵ��%��G��؜��F#6O�"�d������e�lJ��$�X0JM%�&��R"��B����>��l.H4�e.�cG��2'PJ�p�:�9���H�,	���W
��k'��[�v}��zRH��V�-�ZX1 .�=Իˉ��8g�i���e:��3<��.��'4�a����x���������2�sbj(jGr%14�|E���N��dr����4(F))EQc�{���w����K%��Pf�'�3���O������2x�)f������f��[@�=���׿��=��{/���wq��/s2��-�}��l_0z�ܼr�Y�)L�9�mqlT�9��3"��G����k��k�۽Ω���9M9��Q���F8��xLQmS׎{Ű��rjtI�����ܶ3�������ov��$­=�7��g��S�?�4g'���i0��TXL��4b-�Ѭ��d��h۩QI#�Fli	�������()yv��ő��Zʀ-/ljd�ҷx�3s�;l��}��8�Q38��-+N���n�Oxƌy�/~��*�9�1m��V�d¹�M��0�����'����(Ԅ
�3��a��q�8N�)g^�(�Ҳ�5Z��-�E����or�����>[�n�O�K�N��5g)�4�{7np6*��1���0!fdP�$j���
�3�rl�#q��F*�@�5�møQ�D����i4�y`�T'Z����b�3��]��,����&/t�]�	�
B��(Z�$�Y�e��Uٰn8�������о�BN�b�Mh����������*�~Lc�����Տ����5�j{9H��[�\Z�$�����;����ζ���2��d:Q9v���M.����hsh�ҋA[�YL��BTO�jk�����I0�� 5�C�>��l��$G
Mn�e*��CC5��/�45��:$@C"Q��vK��'|�[������u���{����`��%9���8}+����,'X��JY*��G���e���BaX������mmRG4�9�b˲���Ab��ۦ�rm���N�껵����'����#G��������P&vwo���ϱ;�3���ᗾ�;<dӕ�:��ߪ̤F)���d���{�&ݾ�y�ӟ!^y��gOp��_`�[�y����cs<f�`b�u�e�9��D%�"�P:K1o(Iؐ8|�)����r�[�1�ڠ�3gFp���3}�;��uLc�1��4���ͯq���3��1l@b�U.�L��`�3B����>���x�SFs�&'
�j��>7��B
	��,��69ve�W�2m�ln}���_��f�|<��g?���yr���'$e���F�]�������Y^���p�w���n�0��q��&\����y�9���x����[�}��%4�ٻt�g>�G�?��ݢ>s��
q�`o��c_�֭����p�k^˹ӧ%�s�V8Um0�|����_���2�y�=g��=����_}��g}�3�8����z� ]�x��H҆�#'��^��ߒ�7�x�n_����9SL��-�f��AN��L��?�Z�O��(�m]���'���5,0*�">2�����Lj*W�ʂ����9�p��}�_w��7Ə�>s\��yN�:}�}l�<��8��d�j���,�:�.H�KN]蚮!L�'Y������FZ�y̹�a�6lK������x��s��m�DcLKa�ן�7I�����d<�}�,�|.�4]Ag�*b������w�����k\��l�G����c��z<�(��Q��TU5�}�����#�G��JMڟ�;��xá�U8n��N�j�v���Owl��>M5� ��mw��X1X�0	J#Ęulǭdo����!��0��Apέ��;J�U�ެ@cV���!�#��N��b2=d������5úa�(>f�
C� ��#�����U^��? ibxv���)w�0��c>�-f���҄�(>6�M�u�ACH��E
���ʂX���9���W��/�}⛘�c:�ghqI%�w�{;Ր�I�(�M�y������-.'r�*$FH7\.Q3�)��[���M���Is��J�i��ѧ�C�˔���S�$8�e�|��<��3P{��!�KC*�I͆TD�9�	&*�d�䫟�矢ϙO�(��"geo9�N��o��\}��_@�#���X*k8��ev�Y�z�V����@��9[(�ܾ}����f��2��\$pN��D�I�3~�Yd����a�j�b�(7�"���ع���+0&�	��Q$N@��R���߽���ѽJWPMw�����T}���_�8��8���T
m�Q�� � �}v���w���L����N��q����O'x�����Wn�}wx=��8'���&1KP�;E��]�3f�/�F#UI!Q�~F�2��e��R-,�`r���M�jf��w�%��Rѫf�(Y5���    IDAT����+w��̎���!�EY�28�[��:�]'�h�]۶�v���4g[��AW���R_W�]���7�h�2�p��V$��������1��c:%�������Uw_���{\\�5ؐ�4M��G���wC���6�pEٛ�%}W����,�$ �
��ba�^W���{6�y��.l�
6�0��L�G!� ��9�j ZD,�hT�[Z�B�B`�p��Hb�:�~�8w�b�!��-R='�,�׭��KU�L���bҰd�RJ��z�ޜJPjh
\Q�B$�����آ" ����k*�ICjn��!&��Q��"!�t��kF�-_��1�@�he�EUK�Σ�'?�h�f�׭��$�l�9V�(!MT&�Z�P1�!aK��F���n<�e�u��>��Y3���� ��w���7�u`8RX��t
m8n�p�O�h�bn]M��Ԑ'KK2����\~gK�)P�ך�f�a�h���st8]lS�֨���t���]�p6���p��H�c f�04��Ec�h��-��;��K/p����ۊ]T?��9ԭ�&L�@"���a��K����	�%|̃~pBBC�t6���HUr���zh��\��W�fF�iF��x���h���$�2�K���\-��p�/��HZY���G2�7t�s�!9oL��#FZ��C�u���k�4��l�����2-Hj�:�C/}E�f�ѷ�
�Z�*�"�r�H�(<��=�1^(�E��~w���}F���.!��F-�.�����{�������h����ݛ�/>|�����y���UD�ɓ�ܙ-
F#j��0���e�%/w��wP�ݾ����ܳq�M6����J�1*C��DT
B��N1Q�Iu���}�XGe�a:��8�� @�SY�j.����	1�l�w᝔uCeI���F�cs�*u��F���Y���;(I�Ш�V',Mm	�P��#�k�C�1IEYRb>��;��MC��gƹ�11�|cH-���saeI����1�@�lf�Zr��i�{�Wŀ�'��1!yl��� Ua>nh�b#�g�:z0�qQ�U�(�#QbX��b�X�8'���hy4�2����J�k0D��d��y&&+Ή*�@�a�,�*W�Ϊ���1Dt��s�6��B�·V�%�H���%a�c��XN�<bZ�+	!���A|�-�0)b��S�7�����r]���7V>pH�u�yB�����gSUA)|\�*�s���uo����-�����4�ُ�l@i��ٲ��J��Q]:"Җd��x�N�s�w��N��<y��
��+��h����젮��S܇�������tH��[�~�X]�E�Z]YKsj�,��I�/�����rcݹ��tV2ˉ����Y.`�y���jh�(<�-�����?���Y�?p%~���eN=��w?�/��&�(���ic�1�b��7�k�e��â
�=����z�!����+�~�9��rP�!�Ф��i�P�!�@�x
g0UI='f�B�MdPLE�z��4p�
�����O#b�����k�&bj�
4�tĔ���)�B¬�)"$��i&\�D���Ԑ<Z�$q��6e{O�FS�	s�gV�"&C�$R�PRUhTB5X2L�dŝ��'����O�3�&bmr$��R��e2��Äx�@������T(Y�
,�(u���\Ye�"x���a�H�BR���.��k��D�-@"6��3	�*��46�Y�M �JS`.*�G�d,!hC�u3gP�&�40�>��kLĔ����msU�*�X31�f�`
�B���
�qV���&GT#B�5lr�/_�QW"�"��h��Ǯ!�Ǎ����Q�Qs��h�)S��I����Χ!RX�5�$4T��Nk�m���G�ٍ�kۑ��s���ި�)iEL�Dmݛ�ém2�B���AP�ļu�  ��J^�J[� �]������'܂y�x�����}ȡm��(��j�h�:�c�BLkհ
�{�w�/����,(v�ovQ����L�w"+�,�^��'�f<+Կ�|Yw>�F�ݾ���K�V����Ԇ�O!��.f�9&)�q�m&n��s���^Q�ie���歵�RľG�q��N����R��d*@H��-J��4�z���*ےɀ҈�:j��X3ĕ��sj�)�g@��=Dɐ^��hgrj˰@���Iur.��ր������Q��ZdnZ�i���Ȑ&V[�R���CR���)n�-��B�x��$���cH�u���Xr 5>���UqY�+"cta`��ZF�
wQ�i�����Q		)��aTU���מ"���ihNҘ���kc�e��la1�����F����	)B�hH���:�8�1��S�D��W��̢�x�ĀG��b��(���F^ D����04�{���X�b
�N�h��L�NP�ih(���[H�{B�>%H)���ز�4S��W��?�Gr~~j.}�)R��|Y�$PWV����}���su籭��E�*��7���+�;����+��ж�m��Kj��O��^8�-�^�&ۣʥEx��<tQ�-L/��� 3��^�w��ލe(N������UY��BU��]�T<�2�u���!V#�������<�p�;7�r{Y�rt�����RK��F5m�r�v�H8�o<����:*�C��@����.�����;T�gK�g�w���xx_�DQ���?��|�-s*��xWf3�g�&y��0Z|�U�}�`XƎ��}^��Y����v���A
�[{�M�	u=gdGDͽJW �e�MR�pܞ��P��$�hľ�G�>6r�<���3\Y�>�Ĉ)@}Z�JP��@�XtF3�l�HE"����::��Oi�V���º�D=�1N�p���s&�	Δl�6B^'W!*�(D�-pN��s C����	m�&���'�+{<����A I$�H�
���an�SN��̥FS�>�n�4tX���fP�&�a#Xh�y3�(
6F#b��fư��M��`�`���el��(3ߠ�8W�B��V�'f�)!E¬�J)J�ڣbp��)˘p������DR�2�ZnˆT���b���R�efrY�%-�ēY�
�i�TE&XjR��H�u��Q��W�w#�RU�M��D�l��kޛ`�}_���[�H~�8%9p�r��&;;o���S�нqg|��kNl���n:�d٭.���
0;��"WS�ў>Jd"��*��<O��eǞ�:֕|�z.eO_i�1��>����U�&�,�-0�U�2���ة�]@�`�r�����$]vaJ�m�8cQcH1���D�}⚤i��IJ0��ӊ�t�B&�i''������[�c>Fl��:{r�ߔ"�DD
Dr�}NK$p6wpKm�����1,J���{�RB$.>��(�3fD�Էq�_���<�����ql�e��x�r6N��&�7��s���l��ͱ�D��#�� ,kwI{i����+̛�i��P���n����E;�v�;�*���m�$�ɒ�*�6ֶ{-�|B1��i"q����EΜ}� "U�	��o<_�$��g%�T��4i��,�5fd ��]"?��3������ mZk���!��L�2����_���߃)�xJW"�}.}���=�U�Y�4`��zƼ<���]<=T�������)Jn'�R\XSGr,:�U��ڇ�%�Rf:ˢ�a��"@�<�@i
�Y�J|��=�:nϔ�[[���&��wѭ��i<�,[')Kǰ��ao��7`L�&ŹANJ�])�A�ŧ�\��׀� ���ܸC��D���uB���Q��fnd��BTC��y��Ts��GeT ��460k�P����Un�UP�D;#|�1���H�1�el,�(
�Qʘ1���e)���6l�y��q�[��{��� 
��}�`l��H����;8Jːg����{���\���!��
�O1���ߎ����Ƈ\�Dl�̪U����Y&�e��"�J�\o�|&���hXP�y�n���%⣂���QST��ź��p�|�|ܔ�-�Ut�L����5e�c���ڐC2 m�H�٢"٨5Tq�$��k�G/��"DM��U�K�|��i�bH)a�=���� ��ZA��0�'����묟�<,���2՜Q��.��`�ya2��wq{n���[ά��|߆�r���ឿ���Mu��o���$?����jj��4���,��-v/_&̦T)R�cN�u�5�7Hg��R�t���e��d&T�	b�DT[س�_,���4��FM�A��
B��r�KFb:��}�x������E��q�������g��@\��Z����5e�l���JY:�������{�۸��8��Z�!��^�:S?!��j����r���=W�7�eAU��|��6���XG��#ƮdhQ�n=DYd�D�R�i�4��Fq�2��N�v�t�`}�k{���u�m��c��8T5C�k��eB>FFܖH�q�AT	�WU�19����y�&�{]����,�^�cL�We*����y�?�ۯy0g�&5��|��w��w�1Pؠ ֺ�
���T��D��)�޽�?�{�GMy[O�ko����<}4�ò���& �|2g{c���?����b�{�?����?��ƀZVy����{�Dv�/�mwS���gŬєrC��#+�$���˶@������K�_�~�ر�^�=}
�G���)%4��Ik�^BB�@
z�zF{w����R+(��	u�����?��P��9J����e���E��C�Df&�.���-|�mǳ�kHH�O�7�ݺ͍��5C?2o�?9���#�?���Ƞp��p�;��"2�cD[v�eN��x�Eh���v�?����i7~'���9�s��a}�t�����0Yj��AQL��cZ�C����U�Pnm2�k&S�6O������]E\�7�+���5+d�(��h+��>E�8��`����A�s�s�f���Y(�3�Ulq||�o��f��9w^������W��`�P@[��z�������F�F��7¢��<D����'�K$�)B��uC=k�M�i��X��+s�aZr�\K��ݧ�Q���3kY$_gl_���F�佒Ĵ]������-9�B�in~$X2mr6r�}`�
����ќ>�ޠ$�9Cu߽�Sg�EA����޹M��m�
��5���;n=W��ů����#�4o�1{��V�:rbTq�{�8{�����x���8}*|l|����� �J�w���^�Ik��6�2�����}n���Gs��a����C�1������N[�;�!��d}�C=
��"М�nDPY&ӭ
�la�׻x���5kq1	}���}�������댆�;G獚%Z bZ�9�����a�bw�=�@�C�p���>��}���������Q�?��]�c��q���%;�?��u}�)��]�
�0�5Hh��bK�`�%�IG�h����F^�TX�`=�f��v��
,�G7����[��%Ze��0�"	�2�<�A�i�̳��0۶rl��Ɲ����g���1�#Er�y/u@kJ	;�	Ed;0�%�>��\n�8㶸=5��ݲ9�9��a1�%�,�-��ۺ��'�4M[t|9Α{X{o���5E���w	�w��B���F�>'P��)���@��WB��1Bݐ#-RӢG�gIDr�k��Y�r�pڭ���Ψ/2,�P
W�� ��/�I���a�����ҳ��u]��>FT�96��l��v�P��Jtr�sDg����Dڪ��%������#�+����/�ݥ��=�!���QG��w�p㫟�W���c��ql��_]����A&���j-��yQ�ea��U��ms+�Hr��IA�d<cH��){�=�(Z��=�_�IߝGo����bǍ��%��	�-3`j�Esy�t�k���s�0ǘ�2�7����ȥb�N]��Z��N�g�,�2�`����y}�͊�ůw������nd2A	��DRj'؂8�Y(��\����Co�����7�{�������,�׾�,;_�
'^z���L�P�Ν`{I�	%�.�.+�~eD���b�.Yj���uY��+���]}^��m�����Ʉ9�¶js�Д�8�FL�3؛�綴�-
#9�Z�c'���?�H,�mL��-[cG�0P�L94mR\.�1NIMn��bHuf-KQ0��,KF)Q��5i�}`ot!��OW�t��q����|{�����{d��Ҝ�$�h�Q���c�ň���|�+q'Nbc�v�mU��i��oC/!#���v��c�R]ܯj�֓fedZ� ��ܴkIJ�rФ����&#�u�յ�Nz���S���;,�Ո���4����!a:�0Gbȟ! ��tɧ��GX4�Z���hN���F�F�E �Ξ:�ϡ��s����
K�<֜�t��K�z����o<��3�I����;�����kz�eHx�T��j��q(G�M��b� �C��֧y�rɚ�8hϹt�R����[��
`�	4���^�Ӓᨬ�#�<L�y%H�P��po��xb����
�'8	%�&�h[�ߝx�\ޤ�RpZmK��6c=X}�gP�Rae�v�ם%J{.Ŵ0����О��$fE���}�vԠ�)�ш��2�
�_{��O�1����RU�ZD~�e�܏8B�i�9��7��6n|��g����5"Đ2u��ԧ�*zRfw�J�ގ.���g&�}������[�����W��;X3E�y�ˇ��6�$%����E ckqEAH�lx��	�/�dr�S�H1��3�I��LVd�&��[�
h&��n���|�SQ�u͆�$�`8s�L��P7�&&ꦦ	'�Z��q�nz/uHٲ��e��XƎn�w|Z�X��Ϝ��em�hM��������0z���8w�89`.��$��s�W�ˠ����6��`�E�_Qp���=�fi��9=#�{��n�P7�z8�9�e�M���9����QU,&�"4���=="m��甪��QT#��dh�n ��z��\�ݗ2�ܕ����q��/�ꑻ��X1�~���oh �"�*#vX0�5�7O39�e�k��w����~����~�����?�<=��w;/>I}�&#hY����F��t��fi���ޝ�X(���eI�&'�J�	ֶ�ĝ��##��G���9zc%<����X�u�����"]&(��2d~�iA�{������M��'?�	�R�vlkһ��w� v)`�V_����ߨ�(�v�!��w���>���e6�,h��]L�.�����5��"l$��j���9��w�����?�y��z�/E�ٗ��?ܘ�����{W���_}��gW���Mf/=φ��[O�ㅅ�9�>CF	�Ѷ.�ͷ�N� Ԟ2�^3F�'�mEW-��GM��IBAN�\]�e�UC��2���S�D�4�BVC��X�q�f�Q�qdmc�����2�R�o�k�,;��(���X650}�[\-n���4BFS�O=����h6V�Y�IK�t'!�2_,?�����P�#�4�;�bȥ����g)#wX�u�\in��!FH�Q��w�����g��8k�UIq�:">�|��"x��BZo��ѻ��y^q$��M7
밽�k9��-	f�װ���
�H�{:1-dCH�@�!JA���W�ɥ�B��{��9n�)1-�x�g'X���߻�Uiz[�̝���T�y�8<&D��QC=�f��h{�_[��ﳧΝ���zfwsj�-�I$KTLEp$%B�Ȁ(F (P�8����{�XF %@�`æl���H���f���Û�tΩ�=���wթs�}-Ŋ
��N眪ڵ�^k}�w}W��C�Ϛ���Pݫ��_�!"�����ݿ��CG��J�$�&H�!W!��t�ؐ#���ؤ������ⶍ�T�1��7��q>�>�b\Ǜ�v�Sζ��N���k�O�sh]*�
�p��+�_�#2UʬF�g>x鼓���&�����x�rX    IDAT�b�<��}�y`�����Q��H5�L03�>\�0�MN��I��$&#Y�S�JR�7[�tA�`qw���v����מ���?q���m�����{��ι/�5���{�s���y���m^���xO��������:���0����ɖ�D�	�r��(�U�0ARSF��9e� �6��'QSe�b�R1&�P��1_��A,�*DAL��his�jw� un����+�[q�>�Ѧ<�YN�\�'*e%��|ۭ:����Sz/H�w�2F�%	{z�׿�e��濢�kvU����Y�qqݳ�7W�PJ����Lw��|M�ѐ��1�<;�n�i��0>��|�6jJ�hb1��,��x�&+�)c����TMdyx���%��J	�)�Ύ�H�$HFf��s�c!nHz��69PU�o�2�oK�"�")F�9CxTcN���	�HD+�٠5�Q�i��RUn5�Y�o�3-A|��5UV4��@�Bjj�ɪ�u��.O����ṛ�yd>���Q�Q�'��tӸ�Nkj*Dt��8k�+������[���o��� ���Zn��?�G��?���_��k�"'K���U�j6sJ��L)�&	�q��C�Q��I�LQ�l5ka+�,L���r���Rx\zg�?v=z����m��5�~��Dh52�s��(�Qv-��F��	$l��2�o2��@J1�$rĬʄQ	c�B�����&�dŨ�]�ǜ�B4)΄"4%�O��T�Q~麦g%~�H(P�UY&Ԙ�T��mP:����x/��)Pt������g��Ou���,�饥1WQ�����|�k��cҍ9���|z��0t��,��o|}��_�
�9z��n]�����퀲-*t�n ���@���W���M�i�qD��2.v��{�����I�D�y�TE�gS�q�3�"w��by!I�֢%�L$Yϩ��v���2��Ԓ��V���h��hS�y����
���5I%����]b������z�	�H�.�1;	Q	RTDjLo�c��ː4+�q��3\�E���ΐ��<������x�{���a �-G8�9��~Am����:���7�#�X,������J2J!����u&�$1���Z��&�QA%��P7	Z"�Z�> �Ak�u��֠�E��$��}����ۜ�C�}���m��	_�x��N�&��Kv�|�A��(�(�&��[SS#6#V�
�JkE'�%K�b5u��C
�oS5(�@�re,V-�ɳT�HU�f�SUTE]/0VL@���Ƅp"�]CRx�>i��+������j|�XհV��si4q8E�
S9ZS!VѯN�>kߓ����&�CO%̈́es���v�u��B$
Y&�lx�*i��1���gd�'����db���c "9������2$��8�(���÷_������s�w������������������y㥯�OX������TzSU�A;����D�DA�8��,%lTU�7�T��l�s1G�ر[a��F
��*�����!r�PVŔ�TKJx��Mq>3qN�r+ڂ���I�%k�hZEr!�a"������.�㔍>{sO��%b�t�/1��Ӟ_}�>���M��*R��(���H1���� H�<�1U���%*�P�wN���?w���t�0G���\{�u{�>��}:�EQ��(��;�ս����]���z�/~����ۯ����*�}�iCǥKX�.I�N��Z��~��w���oga�4�"؎N7�-,��0x3'�Є��&�C�X؈�5Zvw#'��b�k0�{�rUQEM@ʽ������`[BLT��UZ�C�]��@�z�:�FE���k<R)- �I���e�����ݖ��!�����1Ri��B���cT�`׎��@�Ղ�(N��T�f;)0t��X۰��ǥ@W����E�+����t} ���!iM�mFU$=v�J8Zt�J��ZE��K�����5�$!6K}�1JpN��
�^�l�E���Z�2x�hv*����&|�a�c!5��%d�*z8&ƈ3�+��T�z���gC����·�I4��`�-i�B�L	�9��;���5������º'&��,�.��O�:�	X�(�r올��DT���RE?1L�IB$f�C�0�Y��1M��KC��mK=��Mki���G9�A�J'Ŕ6��nXӶ1F�a���&�����cZyd����{��w�q�&�;A�3��,�U����x����p����}���_W������7�~���u�������'�n }�B�c��\It�4���5V�@�f��.�S
�k�q���������m�?{�x9��I���a�h~~m�=�����a'8}\�Ș�+�G|���W��.��� ˌ	��N�l�s]ޔ:���م�O�,<���q�D/N%�K��(k�ÚI�#:�r�V~�$��;�N$�}���U����������g�x��O8����߬��Kw��u��oN�n�����o��W_�C�.�D����n~���
��un[�ѓ<����[�|>Vgg�y�yy��7EV&������3�K�P�.�h(�[��~�Sv	f�5�W���Ի����k�P*�����X�=K�3'غ[q�G]d�L)}S�rG�\r����AgɟU?��t����P�����,V���Q�ϼ#�ce�J1�5��)O+&v*AU�^7��� �h-Y@Eh\�Q�n��t�����@���$���w��`��c�Vd�80�i����;>��A�(�k*�%��c�i`�9��]n�ȐZU��j8lk:���xpH��fĔHKO���{���#;u!�ƞ��%(O������������DPˈ޻����zRJXW���%a��ڠjAiO0, �1�^/�]C��S1���v��=֘���ɍf|dG)jrI�U��w� ��:��UOҖ�*z�`�wr>����X'ϲ�h��m��qڟP7�̀r7BI�Ka���q,[V����4Z�]��}�c��>o}Ok��i͍<�(sb��V��s��7�����^4��E��L��;�U�;���tz�O���S�������7HGKl�)�1��&������>�T��9w�����^���0���6��y�y��)�W#Aoc���UA�TA��9@f*zނ���>��h���=?^�"��1_�CiS�RvH.�!���$JW�� ϝR[�J6����HibS�s3C#*���C�T)�H��^O)c���d̿�ޙ�&2A�6�;��7߀o�p��5���s�y��.~��v�=[�ſpU���y��_����}6�D�~҇�/�8z㙗��3��ηxP"t��^��=K<Y�<�ӄ �$0��'l�r�F~��Pۿq���{�6�y��3���]��D0�U���4�&b��*��mz�7ۧx�Os����V��_c+�v��"��w���Ǆ| 9j�چ�N�n�e9m����O��>L�,�Ւ�r����^���?�NZ*D]��������7��S���NX�=����Yv�@ rǵ�|���>��5�Z��w��]��~�}�"�����Gy�ß�z�!�)� !Pk�DX��np���w?�ò>^!�%�[op��os.W*��&u=J)�J1X��MY���=�8W|�^@��l��5�n���#8��}�������Dv��4�$�8�4'WD?�!.����6�!�9'ި��O����$ڣ#N��j��-�_x��R;�3
֜���� �?�΃��]�EZ|�[���Ap�PUBw|��k���U;�g�9��Q����Ԗ�`��0,.�C��t^�"�c�M�b���DE ��]����*�[�B[c�o�>܂������!1�Y=�Z���x}�[q�D��()��JY�7M�h������cMݖRM�hKH���<�����T�E��u��{ܿ&$>�ߣbe1�	�Bղ��Hi�p��?�ś��>��z6��������R7�+o���+�����y�׫�7����g��+�>�j-%Dɶ�j�IU��������pt�Q%oUŁ��$`Ή���J*sB�%�c�s΃�X�s� ϯ3��Xg<&�H)*�[o�pLF:Ȝ7[�)�D�a��K���1`è�<�?���q8=)䞺Z���ez#߿<(6@��H�ӑ1ݐ˲T�$2�7�lV@1�s/._�D��Ǳ!��e��hrc�--{NV'��H��Ex�G��@��C��'�~�ٻ�;��nղ69RJCǲ;���u�;�	wnsyX�X�^����?:$uP	�Ez��/��[�~ףW'Rr52>r+��m���(���K6�9��Z2>ϕ1�4���V��K˱j�y�)��Gy��?ϕ��˩�,�M�22�Z��.x�	�-��heIX���&}�*O|�<��_�3°:�>}����������ߧ]�1ڠuC�<����_�w9�*�Ԯb'�r��n��
��anJ���S?����ٟ"�������w<����?z�.��^;���ӿ��\z�Gr�WhJc���!��T�Fb�������?"}k9��p�U�7h�HңTh:�X���8����O��aq�AN�=��k*lJtC���ZN�x�ן�׾����
�wG,*�`+�b������/�G\Z��ʩ�2Q2B�耭j�{�i���$��>G���]]�[��a��ʕ�e�zz}�#����������b�"C��%�F[R�"CB��ۯr����n���o�z�(�zX�A�w�����D;���|�o�M���gI�c�^2��ᇘ7Sg���_{�?���'��۴Iѧ@�@���V�"T�x�ӟ���>�8�*zT��B�=��u^�����⁋��.n��Ԗ�oۖ��jl���0�Ҧ�u�m�Wrf}�	J&}�-h�L�r������H��N�mE7t�(�USs�����|�=��o������_����>����P��߽ټ����������'�?��?֝����9~��,�z�/1,�R�Q2�<!�M3)�@U����s��ض�,�%�]�����=�tL�n��G��(�0����3N�h������6��NG�G?#�� �yϕ�@�2���IR�}3�,�CP����r�WFe��Qd#����-W?�ޫs$s㜬l�Y�#��%qL	h6�q�EǦk�D`�����x�yĘ�G�`�U�V+R���m���}�l�@=�-��}�`�b��4)xb�!wV\2{z���[^{���6�{,q�����8�Yv�b���zd�r.I���v$�G�ܓoq�����Y#��r�g�"S�S����0p��>�q����Ņ_bq�"��N�mU=D��´C�]ͨ�g�$��"C�G�.��n��bo�z��D�p}��^&V;���� jE��n��=!RGp:��^i��+��U�<=��]�-Ƿ�X���F�7���1���ʒj��As�П&����5�4�
V���x�k���8x�w}�a�������vL�v��EZN���'�d�]�`.]�oi��a�n�|��&����������k�����왜�_!<��c\|�	����*�emj*	V~��-.�:n���:��k�΂$
�jRR�̓<��'���Op�Ϡ�H�O1�*�[g#�B$��{�'�B�����~�ݓ�$m�2P9E��O��O�|��'�ͅ'ރ�|��Xu�"�&��,1z���޳��j�&�?Z1)��e�j�D,���|���%�ʢb�D�k ���~��x�����|����r���\�m&W	lBM�ѹ����ENOO999�2���@)UHaې�|����iMO��r��>����4:������gO/`iX�v�b����W��O^�֏�j�����>�k����~���1�籼k����ɴZ=�>��ٓ��/��ߵ��W���w9z�%:�R$j�j5�6`�Q�ޢ�AHw�M_�,?ځ1����-�:��j��l���4�j����P$S�ϋ�a���5Ϯ1��m��T.p���w ��|�gIdrH(7**H��u3 c��8"h�'��Ű��"
��TB�X��o'��f0����P�%�5�s'$M5��@a
K�D��>�4�	R�L5�W�Qj���1U��}��O]D��q���2���t�]eQ�C�A�v�VLn���,���^ᜡnx�9]���!��� Z1����co�i2��g����l~/r�6���<����7�g,�=�QH��+�1�o'�<������O}�Ԭ� 1qɵ�Zac�u��5��>�@�霯jv4���_Q�Y4�ݶ:!p�z�Y:1y����(B�Я��@��ҭ�Ǻ��W��ĈE��%��$��b=at�g5)�S���i��`H!�k����ʩ����
�!��;�S� \����c�x�+��?<�?��[��x�����#?��<� k7ob��^�h��u��5��@��$�9�z?W���|����[���,t�V=m�q�*��TzD[\j4!�`:B���ɿ[ߡZӐ8�wİ~�a���s����-7�naRG�0,��4�E��2GYq�,v0.|�c<�<w����i�"�k�����ǣ��i����Q�w����^���6�0b��v	�tDE���㩏~����_}��Z�s.��QP^��p�P�H*f�7�T��*U\z�x�����У�prD<9FV}1"�PK�[ETFIN{��k�f�0�Iڴ�Ós}�|f�g��XC>+�>�ƕ��cX���$��%�ma��Nw���~��%���������8����u�=�Uu���}���2��%��orx�du��OVK�W������OOٓ���8h*��JV%[�@��JJrZ���k��D�}�1J�<�����K��KÞɔ�\[��n�?��m���A�?��9k�m�*9�5VP(��A�1��#1޻�o�ob#[+��4Զn"��L0��M'LŞ��An�=�1�w6�t��F�vv�сP:3�sz ;/Y�S��9����q�~�?�m�+m�F=���Q>��%g�"��X�#�I�ԭH��F�"���� �Aeb�Y,�Q8]FH�8!�!�1�cH�R#k�F��������^�s��:���7z����G�&~s�P$/�Z)$)|��͂t�2?�O<�臼�M��Kn���;oA}����w�ikN5D����z�j�u��gV��ۼy�m�,O:v����(Q:�R�G7T\P{X*��k	���&�t�c�Bz�u�+�ĺ����*R{�K
�:����TҲ
�$�KT+�hT�q��[�rw�zg�����}n�Sg�!q�>���{|�g����t'�I(�2,�y����{��p�o�pq�Ry�,WHߓ�*D��]v��}�^�������������u�ђ*�8z�G���\:�t)����Z*�i"4��KO��I�:��5CwJ|���k�XKoq����G8��U��ǧ�6E�Mv%�p�
k����"�ʥuIs���?�Y�����wn�O;vm�����>��~򳤽]^�u�������a�D�g٭p�zX�]vv���	N%X�ّ��r��)��$�g@3`�����,R;5ڃ��O�{���3p����&�|u�>��,wYJ)�t�GGG�q�eV��C��gS822�g�ks�6�次��������d���CU��@J���X�Y�ĉ(�M����+���?���˸��_F\�`/SM[[N��\G��ݒ�:f}�#&!u�5�>Ѵ��Vc�RJQIpؒ+�A蘇��qV�@Jt;6{RJM�;����(uWk�Q��n�`TM��|���"C{�Z��7%B�φ��Q�v�Խ��*�@\�)?�!d�$O,�UV����6�IV�d�UmJ�&p�%��c����B��$T&7�Ц�L�H"�mT�92�'��h*��$b��k$d�nI�Ky|P�����#X(��G�#g�r��k�#�63��3hhb�,��U��U��M�	儔<���5$	i|�*e'h.��H&\��rmmdD*Z4���ʊ��.pN�v    IDAT�TrY��4r��x{ږ��}͛�2H�_�'jIÌ�$3ORJbI�?ź���#��|��~��X��1u]㗚Z����7x�w�̭�~���ta��O���^z���t��s{�����7o2�:b�X$q�����B��e����m������bҳk*����XKM�,���h��
�j�`1��x�F�9�qƱ�
�r���{���-�|�~韢˩_q��'x��?�_�"�4ʲ�V�ء�����p9�$�Q���nh16辧m�.�g"o>�%~���GV=Q*}�}<��_D?�A�rE
�9%��=~�c?�W��\?�Ǝ�H���?�/�]��.�����'�K���c�Uo}�wY�їX����:���6�	mױ�G�y�s��`|�T�Zѿ�?~�+���k�Mͣ�������`�`� Cϥ��|�����I���ܼ��~�Iv��pg}Ⱦ�B����:׾��i�w�֑��K���}ܣ��Y��څ!��t"����B����0P����4������_���C��x��;�������O�M��քe��	^��F'�9����Q)@
��!>pr|�bg���s�'�ڶ�o��g�n���3�!�
0�ͳFk���
�FD7%[A�t�T�(-���f�#�L���o�4�@Wu� �0�q��c;V|$&�X��
QBY� �/Qs'�q��褚���)�Q�<�9tU��,����J^R.e�`U�V��"}��DT�s�@��\&���@5���&���|��uQ�M*sj�G ��V�
��r�H�r�j��g��1�����F�lT7��ǭ��1/$�闊��K�a؂K���~`�����"��f��Xѥ�~~N��
�,>����-
7��M�-ͼ$ #@ܿp�B�+m�9��G;��\�%E�H�bܘs���3�٭|R>�Mfg܆�d�/y( ��n����n�2!�2?�z�S��V��&�BT&Ed��R�-u]3C�Я�����|��?�΋?�z�5�!wbR*��T�F��Ի��R�"��8�L�(����p0��h2*RUFi$�ҋZc���I��S<)���Ο�	$(����2��.mZ�m)���E�CL�������7�C�7��o~���H��3�KW$���ƚ�Z��Z[a�&s=��d�*�!�s�:/?�]���%��i~p�7�k�*����Б����q�ؽ}�| =G�<���	XSM�[�\����֍������'�^�q�O�6T�A��`�^f��R��wD�h�fu�o|�Ox�k_���1�v���ÞT�s�'>LG�J�Bb�`�~���%��6->�Wz�薪1�8S��[o��s�D�y�6��]�J���4O<
�`k�R��i�^�hPP*o�����k�Gvh�� G���ы����Q1p�к�=�~���]y���2�FU��6�B�gL�	cTFQl�!sɝ����aoo�F��:�M�b�������{^08��z��h��h5�H"ab.��J!�(
��a�f@�B�X��/bH�"(��Ȉg�����C��z����E��'�1�!y��)�9�,�UDJ�_�9�i<տţ����l�Y*豺g�tDlRJHx�1�E2t?��B�!Rff8�ߺ0�0I6u�
��]P���M%v4<�YԘ �#V��5��[�H0�u����L���������DR�`�l�)�)W��1wV�x�[0�L �\�Q�S2�$���\�|���cy6}�K�de�j�ȷ���P|�旕���[���;�(O*w�gx/C>?�:>��nCVw�U�����
?yװ����{��z�t|Ⱦ��J��B��M��!�Ecꊝ�ss[��Q��(��R 52����`�<��(k�^>2(�Pv���\��;@"���Y���Z�Җ��>ׂ[�ڲ��t�Lc��o�^��u�&���8��fQ�P���MvZ��>���G�t��SWC��}�E����ܺ�7^|�'���ڊ�N�hQ�UC�X`��)���N����Z�,%�UZ�@Z\j�X͢s��}�)P�
���K.4��}��~��'\T��$���~��o����8K�#�0�Ȣ��^8�OYV7`������w	����D	�"��i�%�@8`y�����p8!�����Vo^�JS��E���Q��N����Tq��G\n�b+H�����{���'��/���n�vQS�
�Ae�mI�E�Hh�P$bt]��*��8�X�����v��`�6���W�6{��<��Q�V @���k� �����9�)(pɧ�����n"m��:5f���9"�8�� =`%���0�������Kv�Fw���p�6�>:�YIu��R�4I�Vk�exs>�y������y*��w��ԋ<7&�Z.k����J3)ޙ�\g;�@��	7�YR�v�u���1�1�{$�1���ne��9�?z�M����q �P��a��٭w�M�s6��:�R�-�a%BT��/k��V��J9��9��a��E#f���4ϓ!��������dU�ŒF��ilG����l�d�o#%�##"*�H6{�zJE�7�WN~{f���Y��v�T[QlJ��)������XЍQ�:)�=���
vFy�a`HMv� �/9��и�f����kTh� �8[H&kNF��7�R��"#��Z�Q��M]�R�C��%)o�7��6�J��yIr�e���M)S$����	��C\�,\͢q�8�f�5�0xH��CݒB�DЕ��M� �����E��(RT֠�=�5���IF�ZW���u��I�X�s��fI�9,*!C�&	���k[n��HP42����ؤ���	�a ��.e-vg���G�I���
gֵD/�\��$U�2�@2�XM�.X&����Q���'�"���<FI�o���|���}b�Y��k��Q�S���Ω;�J��ҙH�e#�:Y1�.-u{�7x�Ͽ̓�r�C�$`�:���x1"!�E� B��oUN�u�un���M�����=�眵|��F����(�O�و|�]7�Mnh����C��S^9�����6�Dn8���F/C����M��U�Y)�t33���@�InKR9���)���Ƌ��qtf#>��s� ��j
����-���S��e�O�t¼:nn+�69br�m��������������zk�}��ōO0i��s���0�n.C��0JM~�R
C�!�〗DT�.*�q�*1�u�)��D,��'`t�lT#�ʔ�[��|EH�	ʙ���m~�������ܢV�D�����S�]�2�EΎ��$N*�xF�e��l�2���c7"!������N�Y%AFgM�u����I�K�C�~5�ڱÄ2��3Hn��Z7I '6�[2��j���C��X}�����uu&1ڈ��pC�����mB)R��f�����~�s8�r�k60����Z�s�����34�rg}�:U�*���@�]c�"n(TD���:kd��0�D���Xa��sw6v	I��:"	�ѯ�)�j�1
�����c,2K�X,�s[_�]�q	�§�ђP1����Gb�u5]7�z�惿�+�V/��V%*�%f�J�5N9���j�{B쁄��!*E ֧��!�b�g��Ћ&(CЁ������s�(��g=x�"#:2�=#oYH�F�61:�8�K��}�ָ8p�>��@k�Z�L�?������hnB�P�P�׬+�1b篿�4�dn�C�>�DEs6\��OLJ�yr0��ϕ��3qiz������0n
��%�r�qr�t~�#|>�}�����]^xv?�*㩪�����L��H*.�~B)��Bb�	���;��e%�.CØ���!�!Q�����<�����O������	�ua3�0}��oR�*�(H��m������X�'N��u�}3�bR"Ā��۴:Z��K�hw+�5��5 �$"eJ2a�(AYP1{~��r�bXd����Sl�^��T"{�Ȭ���T
̔6�4L3�h�����l��f�j�!��:z�J)J������ڞz̡�^:���~���Ҭh��l��b�!��2%��y��%��i�VI�+��-:j�1�{�y�"��)�1�G�Y��(4l]w*��T���ᛜ��HZ!���$;ƣ��
�/(�~�e[1�	2��_c�%J$�rJ'��Ԣ�'D����%��TS��u_��!��� ��N�CB�ߓ��RYTЈ�PUD���*S!�!Z���� *��j ���XD��&j��K�c�H��d�L�<�1�c]��A^��-��o-�����t]!uõ~�}O}�z_J ��1�$F��AH)fE�����~�Zx�1 �gR�kI�u�<�q�N͑�I1�45Cף�&Y��T���^錒�	`���6d.D"7��i���.����fK�ĤP��nj%�&�p��^h�aYh�Z�y6wQ�6q�D��A��z:���F��S1�,�5��!��rJ�]Q�l�"Y�/�Hbێd$yT_���k���s��6���W�������$M{��j�]�|"5J���:���s�8?%:�|��0�yDFr��Vӳrg�Qˌ2259�1WsL�xҳP���Ƙ����6y��;�@�H��E)! �"!h�������Jal�x��Y�Ltf����QU�mkԐ#�iv�������Pe t!z���\��0�G���,0U"v5��I��}�����+�mC���go�R�����d�ߏ��nW#ObL�(�w;og��y����k�k���o�M��`l���Ҩ(������&E�!ԮÇ�4i��T���C�D?����֚b���l6��"HPJ#�*7Re�,�
y�$�T�i���prk�(��<v�rh�������diS�2R}��&w�
2����)d������
1�J�i*��&����$$� �Dw�f����uĠ����J�D�������@�2ԜB �
S"�q.�ɝ.s���-:D,*�\�c&/j�(�u5��CO
�ֵ�Ҹ�B�')O*����#�D�C�V�H�2�S
g�G�@`P�p*��P�e�ם�d�uF<���={f���܏39͢��1Wi!e�b�	�p��h�r��Sx�zh�kX���֘�3�
$��J��}l�&��g�랩�k
���I��э�=���=��2���STs����Q�{�HI{D�a�7NKa\��J����q(8��}�^���3`�p�6�h����6����v���X��'��6(]��e ����΢��|��ђ��7���@��t��&�2�\��ķ��w������!�hn��si��
CH��>�д�D!mrm����uE���dEP�z�����4Ld�B�p��U�^�h�1	�cfJ}��or3���LD^Dh #)��s�d{b*Fv�B��mn��ЛY�y�Ő
�f� ����P"^����4��
:�9��,�ѐ�s��6�E��t���vbr��*K�!)�$�c���\�dF-�R�R�����I��q��F�ژ��͝S�ƪ̸Oĉ<:"<�F��T���M�t)�w��bw�v���1� ��$�$���O9�w.7�!`#�T��ʦ�@[C�#ݢE\M�*�������=��&>@kjS�{hl��kL�U$�i4C���_,P��6�$B��K�29�<��$߳z��B��c�Qc��h���G2���u��C`A�.Bo�N���8�tͮӄh|t �nuB
�=1���c�w�I�+h	�xj%�*�7�k��E����;,�3d�#�`Bi�����[C喴CP�ڀ����j�!F�z���i�Z����ߧ�x	o-F:i�JVM	��E�J�aU�S���bn��W̜�iG��.L��1��[!W��(2ߧJ%�]N�뗷*������Ԛ�ύ#�Lه�U'Q[�w%M�c)�6?���m�M��9�Y"b5��
{���JJ���~��*B5��!D0��9GJ�{�h1�\�_|�}ϸ������K��ѫ�#4�]��J"S挕��AѸ;���9P�7 "t�==�4)	C*�D*�|�ǘ�̑[ހ�Ґ�ϐB��2a��06�Nl�Y�d����)Xg2�W��A�e8���;O\��i�BR �r=���ͽ�D'����Jg>KR�ds��=媌��y����#���J�@��<��L�֙�c�"��c4܀DGB��l�h��PSA
��Q��?�<L����ɐ��X�Mf�h�%/�uo��s6D������-���"�H��/oo�#K�����,��y�ں��!g�)�iJ�H��$ >�I�z�����7�P��Z(��������t�twM5�k�[w������xDd޼�B�neF�G�v�����o�A>,l�$�@�9d6{峠���4m�aCv��y�Xx�g���;b��RIRpő�GZ@�5̤:��D�9�z���h��m�)"_�c~Y`{`�GܔBz�e��P6���;nE��7>%�H�D��F��)�����H|ʢ�x��3������� Y��J�h�P�ќY|ķk-r(<��� ��-!xJ��ё_4�qCU�=�Uk%� F����HkZ�#���[�^q{3�/��.����Ԥ��isb����v���-�^���]�[(ۉ�)W"|�U�}�����̰4�-�i$�\���!G698h�0|�9��������o����
�b��hb�\^�xq�Sn��qqӈ�g���sڵ������0����'�q�k�����1S\�yze)=u�!���Ȁw#/\��K�*����$,)�j����fr�x�e����b�w�e��+_�ˑ���,ё�0���x�;˜��<�1��o��`j�]��ȩʹ;.�����������Ù�n�����T�i��j�z{sR�Ɗ��S�su��Z�{��<�?�&��Z��Ҝky�RC�g��Bk���rJ�����B�V�U���HA�-��e"��~9z�~k�r���;�KH�b"Iv�IH��U T����W�As]pN^*'��� X�3�pp�$!�c����i��=#��
N���n��A����o��d�6��qq$xSAg�qJ���nL�Z��@�1�;��R�E��F�
�����'l6[^�|AM��fC�2/�ݛ�>R�9�s+�)�\�tт�k�,goQ��aw���ܛ�������x�R��W�A�k���}޴�	�x�oo��M����w�
p�����%�4tH{�lܖw�H��/���Y!G�fƛun�Ҡ�֍>��Ѽ�kD��=��f�2/ٌ��3�܀.D��!�>�n���7H�q�a�3e�e#0�B��"�"4b7�a�m��������"Yf�)S�̜�"��&��`��֙�Ҙ6��7*�r�T�eF$��Orf9����Ss�r&�?�]Ct�Q�!nF
�Gz��M4�1ւK	�#�zT�W��w)�R2�m�o,_СB��$ZQ$��3��������\��������3�-2������?`���>f)%R^|��2ĉ�y��?��<�����:��[�af�|��F|���/^EG����_a��!U-�#c�Q|ʹV�!ס4D#18\�*��8�X]rl� ��y��R9�:��"��|�U_�(�qB^'���y}��"�_Qߝ��c����|�g��_�C�Q�]ù�k9���_�F��۩Z��'+�y�֓{h�ٹ֎@:g�ޜ*s�Öò���FJ3O]��r���՝uOϜ�*���um5D�=�̎<7���:���������	��.�brF�[7ǉy����A�k&�}�u�w�j��s=�n�3n'�i��I���Mu͜ǒ�ï%v̛C���.7�͎F#�D��1��g+gy���BKc)���:چS������ո�]�䤬�|=�(��3�BZPWy�C��C�s2�]�_�O'�$��Z(s�����!�BB&�|���iL̵�Ѧ��Ћ�����OD7 2P����J�P�z���VHe!��
87j��h�P$���/��1m�D�[ F#��T���    IDAT	��Dn�bMh���E������L��P������VR�OU�b(W(���TmK/+���H�̕���X��R�nwI	��%��&��C�.ʆ��%i�vxm��-���e�P�Ԗh� ���Z�aB�1�BKKG*-4c���Cpa1H��H�	�VQ*��@��q7%���L��}�U����[b�F쩞�+�.Ľ2��8��GG��7ҋ���-��)P�)��y$�Gj��WR�4������㎱���"D�\�]�)[>�)�eI0Y�t��[�ꩭ�'�PO�M�ZijUE'��� �>1��SϠ�պ9N��q�9���6�lzL���=Z�������A�)<�%����My���5݀�1ҧ�N�;�u���עG�-�Q�PjcɅ��	!,-����+.�#�%�4���5�U�Uzk8o�ٚ���9��8>��:��׻�}�ݹ?V��s���'x����V��¹�=��:��ʉ�֔���l4j�����ĸ��곟������};+�w��9!zo��#�O��o��> ���;O�c �礔�Rq]P�n];�NqZ	���:����y�����꽝�J�,����x�o�n�����E��ﻟ���kn�˶SU�}g�T"�e�FJNL�:P��/���#���yn�gi��-O��M���~�Ϟ�ɇ�Z;���>���Z���5J��e�Pm�hL�X���T����������}^�uq�\Q?����g����\�@+3��5�RQ-�h?Um/Z����L�y)�M�0È�ᘯlj� �F�Fi�3,�e��b��R
�9�!r؛d����G<��OUH����]�U���X�zp)��w�«��Ayu��E��z�W�َ�i$5G��h&p ^������ʡT��
��T�5�񔋷�~�>?z�){�:���ls�
at�1]sq���F���ea��7x�o������(Z�r�����}���{E�Q�b�LKPn������ȋt����)���{�ʳ�����p�A㊨�s煜�EM�YXJ�UJn��L�0:���L I�����
��c�&��	� :C�+�U�X	�o��O��G�Nܜ�Q板�� ��m��������F&����������܍�ײ�7��/�N6�絓��?"Ъ�P���*2z�*i)�l�;?Rj�u۸x�蒖�^='��pѥp{UwUݑ�sj�V�:�X����"���_c��z�{zIj8�3�o=�}A�j5��u��q�&z�s��wBc����^�4����e{91n��jқ�U��V�b�ά4+Dh�iՔ�L~ձ6 <q��b���4ܼx�&�cm�c��ݣB�����#�&w�a�=*�?�ͮ7��u�	_q�5���Kx}»�C7�(�����M�7���Ŀ�Ϲ��jtN����<U�ذ�-845<���<�����w�/~�?�*ף�4+���C䝿�ٽ�.���e`N��]QJB]�:׎�[4L�Lq`Qz��v�9>L�J����[��W����K˞��l2����o}��>Dj�%ze'���s"B�j�F߅>������HpxA���h��Z\@|o��:3ٙ`��^2�\�R������0m��|��9s)�.-�����[��R
�J������m��k��t[���W�%�W�B�n(M�U	"\u?��zN��
N�n���=>j�Lq�G.�/��Vn3�*'�~���}��I���q���o~�/��مK&��7|���:`���,�뛰q�q��7Ҿ�G��� 8�F�%��)�֘�t� �L���7y�?��y����Ң�:������p�X��w��+�5�0��G��r�� 4q�a0����$b�ɚx�U��R2�����hGL���9 ���~��Z
����E^Ϗ������j��Ί�5�iԳ^�E���79zf�T�:=_�;"���&�`�z�8��#���iv�Hn��m��U-�Ξ�*O�>bw5��7���{�2��):_S$�p�xG++��S���:^'��آ��������?�s�7Vhǈ��q�܃�wrV���=U��<�W�I�%��BΉw�{��������Y�S.�7P��}!U��T�lE<��~ֆ#�4������	Q� �;�G�=%��>)�!���z���GO����}�Ǒ���_�v�#��������}��I��v@s�J�&hT����O>���{�+���ɓo|��g����m��x�og���Ϙ��4t�
�%e�o^2uU( 7_��O���o�:���_%�n�-!񒋯�:�)r;�4�w ���	�0������/~��h�/q����\i��F.
^�ԛ������v���uF���Z3_�Rs&��͒H��s�f�.�E6W�}��|zq����r��Ƒ������[���0ni2�5<��׿_�����������,������ۏ?"�f}�=^��I�q���N��(8�|�W����xs���������?���Oٌ�O��?�w��=����?a�����B����=�����1�9CHz�"�p����S��~�g��IQ�(�.�|�?����������i1B�G��>o}���pK�����G�0Y޶�P����x�?����1n�8��Ѵ0��\3[<T�]�`�J,sk����Lo����"'��Y@�e�ۗmo����j3�k��}Dﾝh+
�@��tU��2������>� �ڀ�E^;\/�c:$;�9_��a"�b��^+(�[C-Q�~�)�.7�t@���?L;r9!+�Ѵ&�AZ�X�x$a�ms����A_�N�/��Ѯ�~挡oнX[�5��ЍT5(����|<�E�M�̫s]��4 θ��X�
�%F�)�<��f�#q��I�L����Z�b�xg]� ��'PR�a�i���_���rb�ݲO�DH��}k�H��cmP�������l��P��-�xh��{��&��]��O�5�v��'�}��e��8�r��ݔ�닽s��Q���	��y����:����bb��أ�!*��������-�s6n�&����T٤D�������x";.���Y� na��:�SBQ�af6&�)_o9��>��������pkI&ĒR�Cu�S~ә����(3��\w�^��C��VZP�-*���P]����1���CCD��=Sl��O��������a��o��ʾ��&K�'�����F��\T��b ���'�����ǟ�RX�5v^��5��	o��>n��Ⱥ�Z"��i8,�h������Hm�)N�Þ�����'\��_��o�� �N<_n�hQ_V��(Q��ָ#\nɢ�mA<qYx��������xk�m��_"9eR�ٹ����w@\FI��*�?�ea����f��J�����U6�3�J����*KɌ␢�������w+���p�v��o����/��k>��ȕ;j|��|�E��E��<��s��F�E�k�rV���~�_vS�U@E�;���=�
��ݘ��8������ȕR���еM�ٍ��˫--^|��z	p����F:)]�%{-��3�F��(V�z?�r�z���i�u1��qM8�U�;ό�EFZ֕�~�N���Dlpg5��g#"L����9�-we�@Ή���w�y��-^���9�^0�C�.��8!-�ی!�w�<�)ĥg^b8�����"�?���x}ҬZ��'�OTO��iP�ky�7E���׾�l�?��S,�����s>��u���5��1Kc)W���O����x��Ox���wx�k�3m�,@��=ڟG!���x���Il��!:�?WoF��5?���'W�3����]!�Q2Y3���,��q��X��������;/���J�$ejɔ%�<%�� Έ8�FX�a��E�L:�b�9�G��]#�ǉ��D��F�2pR��j��Ƹ��e�r�����0z؎�9]��G���O�oʿ��/�5�i��x�~a�3e/.w;�����>�	?������\����c.��f��?������������ʯ�|Çƅ	Ke��D�0N�\�B��ю9F��l�O���W�?�[�����!F�\癋�dyT*�ژ��SԓS%o_����Ł��=�'#�ӈ���ÿ�?���W�o�y�U"l`p�7J��ѳ�4�D�.hs8	��[J>0[|�hK�A�v��h*�=O�}����u>��}�;i�5�I��_*h=ٯ^vk��w�SQ�_�|?Ԕ�|��ߟ���C��E��At��u�ę=�oWZ������f����`eٲ��-�Nj:O�S�"JO?x�i]��;[_�����5���h)À��W7��y=KoT5R�6#n:'���(?~��]140��y��>�w���-���>p9�������c/C��h%�`ƢS'����V�)j'�̛�V�5B��8r��b5�*6��^={I:�<~t���1��W����ih�	s٩cP!:��XZe.��G�6��m�{OS[���>
�l��"�/.-�!�E�
�w��c��7����V�~����מM����U�fѹn��w/�*#��;1d��u>fΘ�j�pT6<�h0���O��ث��Z�Jw�:D}$"�{������u�a�w��rF����?�������6��:�w��Mp�)��W�q�e� �8����?��w����'vߝ���-���,�O8�k����Oqs�� �C�Ej�&�|��/^��~�?�S��5;/�[e��*������-���P�HnJr3��OY~�CBI��1z��}�������������4q��g<���PZ%�G��x�������w���e�x5|R^����?"�����Kc\f>��?�>�����?e���PB �"u#���*˼g(�����c^}������mD'�8�j�r�|�����m����&<�� ��:QO!�[b������߼ :����������s�����a٫��u>�昞σ��x�{��v��r���Dɉ&a���?���k���������	�y��+�hU��ߝ�V+������ǼD������������\\0��.sV޺�r��#���{&	��qB |������W~��x���L��w?����b��,V�� ��������\<�u��0j�H^0�1A�b�����4��E�+�f�	w���1��;ST�$���91���g�[�j�~��[���˓��6��]t� X��f'&����0�V��|iU8�5��(���a�h]����+���d��`:��N�DON�T*JN���%)�A�����Z�Gz�i|Ņ`���� ukYx3홮��P�Y�z�.2�ڎH�&��;����?�=�bd���n���{*��m%1��j�:Q��)�l
e1��������jI��z���ڼ*C���W�n7l7�J-������W�x�BʕڄF82E+�����&�i@���Z-�ܩM#]���*ռ���6���4uq�)��=��z$}>YW����'�yO臼�_�ٶ�����{��u��,�,°�Z%%�T���wb�J��Ȼ�}���1Ҷn�!.`B�]?V�x�KaօA�����_�����8d�y��%7M�8R��=cb�iK�,��U61 �X3q�si1�B 5�t��f������5�)sQq' ��S��(���9������ng�8q��v���gv.RnMhŗ��\s5�D��[�f��6�H�[s�������s�,��d�a���61��=��Q�j���1��)r�!2�	^�H�3p]�X*����
.7u��f`.��?��xZ�on��]�����Ы�������s��(�R��T9(���]�PepB�q@�,P+bPk����W��̣ݖy��4!>}�!0��㶨S������]PU�i��[�tA|�e�1��fp�Zx�٧l�:#Ū���s��3�՝9��o_�������U�Ug�j�.�������:��7�_�/߯�{mn�T �����~�~p��vF�[mO��;�:d�	�k+W�I��S`Z,��Mii,K1a�q@UXr6�,�0:6�@e��oQ�_g��FFM��L�	���ة�'�!@����e�xk������aI���g����WU���&܎�[r�a�q�����ɷ�A�Q�Q\��M��3�6��c�x��-^����3;�\�io����sF*�"�<H���4�7{Б���0��3iص�n[sW
RM>Z�l=���%0��'=��Rj:��é�u�p���qx�#?a,���]Ǟ;�g�����)Uz3�S����>����������{±;Y'#��y*�����m�|(�S����.Zz��)g)=2��W�c.��� <ǭz�ɤ�$
/�k��U϶A)�	{��L����˲�� �K��[kA��'Z �4mv�SE�.����".�V\̈́ D��4J�t�v>ࣃ Rf7\���=W�Hj��!��zIrJPpNy1?G/��fN�J����0�����@��ޖ�gCu�y8�]�h��oE�zOOp�Fz�1�4v�i�����)-�a�b�c��Ak?��nSX������	ڔ��F���]#93�A������g�l��H���V���yk��xo� XӡRL/�f�_��q�T	���p3^�U��a� b5�RjcS���9��J���_����f��glǑ�y���46�3L��U�c���%U�g��juV�r%���A	�	α�C� ޳Yc��NT�:�w>�Z�G����U�'�~O�9�:b|D����sJ��9�ֻ�q�z�ۂ��e�Ϊ�̓���vg�E�]�������}�riһ`�E>gs���ܹ�Cp��	%'��X5��`]�1:CT�RK� @N�Z*�
�������s��cٰ��=���ZMwv�>+=��}]�*�4����sZ���|�\ί�吾�ٓi���/hV㪱J��.L�棂
���͈� ��"�e�qL��0n�ˁ�"M��hT��\v��ֺr������K���e�b4A5�U���X�e�681��A{�n���F�������@����^���9Ϗ��w~��ϼy;}F��O8E���ؤ8r���Op��d��_e/�c�^�ڇ�j�	=�Ph��L4op�o�k
Zq�C�b��A �@��e�joQ���"�6�6f�v�z��di
��xP���ո �adlR��j��0������1�*�Ԁ�!�Hs!W��o�ugi.�&�ò�H\��O//�|򘋋�_|��g�y{@o
ZaOd)B��\�������@k	�-����D<T�/8�pq�0]�����8PT�(���Oog��	i���Q',%��#8�|)͛&�8��ni���E������qjg"\N�s�V�b��+sl��{4?�UJ&��s耶�G=���s�Ł�<дr��A�'8ӹo�����٘�gi����8���7b'y��RΙZ�aڒ��4E�0�X��1��09i����l�r�ŭ��� �j���9�����3��AY��F�}�N:�)nܩ���b0�O����<���8��Z��ޯ�k��d��q����\ɹ���@�f��^�Mb�Jo��x�j�S�TDgr��HK�ˎ8RZ���62āqp�m`��ymR8�b9����D����?�h\߂+�+��,���Ya�vl�Rm��Yg�v����6�9���x	(֜c㱽��"�8�:,��j���9�~k�pXP'l�-�9/�b�r�\g�����{H��eZ��_[E�������a��	�l�]Qs\�q!3�&���l����'��u�������z��oJ�2�}��|\}}���W�	�?�h�J��k>��5hQj5Czl%�J�6	�w���+�)�5���8m�
�*�C��`������8g�(��T7��"�W�bP.Gj��d�Z��t�-2'f���    IDAT3y6q@�#��S n��f?��B�F9�]]�|@T��JTK���@¢ޯ=��O^>�˟D]��-e� sZ�(ӆ�m&��f޳�'V�jR��&���xҾA�Vє!���%��X��U)s}����6S��؋3��0�@{.4e\U�`�JM�.\�RN�Ω��Hk#!'�Y�0��;Hw�E���cMK]�&\12(�fV*%%�'��<��z˱�v\� ���?x�(��"��2�%(5e\�h1���)�2�L�.�b�#Z�;T�;\���v��w�7m=X����[�����o��i�*�찵�6�G<-:v��K,�S�<��nk��ȞR�pJ&��q�P�d֏|���y���ˡ�ڀ�;u�)o�G����p�TH���HU)d\T�ad�N��U*�$���#�-�bך�FZ�qc�Er�l.6�&��7�
�zc7m�}bV���u�4����y\'�y͎S�3I�<�Z-8u�\Yk�b���>:�[����h7�[�"�Zŭ7�\��$���X��H�VZQ��1���`�V��.\ ���̤f�����a�`h���EI���B�!���Hˌ�B�ik�pJ&Yh���J1Q��������ܝ{�H)P}���{kj�o�ݽ�}�o��׶c��Ϝ��xY#�3퀳K���z��w�����k��BBt���`��<�f�;N	ZPi�V�-�Ur)��CD�G��s�}�s+4��8f\�N������s�i�r�J�vn��8ǒo{D`Q�2�~���aAZfF���H���$��QS��7g2�4��4�§?�!Yl��q��������?�q���~���L�3�ʜ��W\$�j��b��C���R�76[�^��.b;8��L��x��v��P���%%'�7��4��kj56�qHP��SJ~A<�������=L�g+օ_Gj.Х�+m��0 7@ȿD!�h���֖��-��G?��j��S:byr�-��т��8�r�H��3�w\��(�:PiH��2(.Ѣ'���J��i90��q�֮���E��������=�sڣ���=w��g�P�q~^+2�ϻ��-���(����|_��;)�A#՝��~Y@��vcus:���}�T1e���>FTzN>���＄R�W�l7#--����>YW�U����m�!�,kQ���ZYrb��w��R�䅚�UαJ�ZZw�]��Q��m^:�pvmb)_SM퍁��	�W��v���+
qN�f7@��g��9w��V�܌�c�<kj\��f��2]]�,ڼ���z^��������Nxh�����0db�a"�LM��U�I�ȃ*?�D�T��b��E-�r{3���v����z6�׬��w�u�ih�h��7}}��Np��d���A礗;З�>)~����s�sbײ2m��,�+le_���>�����+��w'
�!���e�؈	��m��`to�Xk��a�x�(���;�A���V�8��?G�Ԅ�y&h�hJ�>��0�TJ^:D�gd���^^�]#���!h@�����ь�?�F�2τM����F�]g~���=��h-
m���h��S�k�}�1��w����� �8�q2Ԥc����rN���q���G��K.�^��e!j#Dg"5��2�),�ď|thӖ༕��v$��8K���k����>�n�َ�Pg�Pc*[>z��\�Y�]#'��GU��l�=��X�K=N��~��0��=�#y9[��h�P���Gk!���j�~S-T�\1�$+��P��)�,� �5ѪJ�.��y���|h;j���������7U�#^u
H���u�����+���2@kK�:�x��O�s��:�IM�Zz��:��6(9�vߏ��Y�.=�݈Wؗ�;:P��׿#��*]�&k%�d ����M��񀋅���[��o������$�kn�ڬi��c�~�����C|��_�0=}������\i���N�%[+�O�Q�j���#��?�g�=��{_{������4�WiX�������u�jzT-�8�R3/�ox��i�>�M2�J��PGZ�Y�W"�ŎasA�������yb�-����w.ނa�fk��B]GQL�Mз�v/��@=w^����zop��v}�������C�{;�.x�5{�y����*Kz�@g��M��Vt@|�(�!���{AKD%��`_-��L?6rQnK%00� %�Zeh��|�<�ޛT3xV��]'_y��N�2&e�,,bęV+1�x7�RcVB�h���4��!ѡn`����$Q�ȸaPG)�P�8{�iDŴ�W���X�<syq��rxyMI�|���~�>zƷ�������	� �Ţ���P���Sa���V��ŅRl<��:�(2��sW����4��{�|�^��Uٵ�d�͞z�Y�b)�q(.8|sԔ�aKN�J#��8�[F�\W^�⬼`�B��*%-V��Fi�z)T��#c�||[�yyŲ�Bo�-����M�k#�r���%�K9�\���٫1����J���E �#�^)ޱێ��zs�v���і���~�m������z�����Νx7g�6Sz<��^0�w�Ȝ{�s����w�-��z<��J�ﾱڜc�y�.�T�� �.Xt�NΩX���q.���*��8F?ݡ�qxuC��!95�lL��nlڬ�M�/�VR��6��͋����0]�_|B���ޛ���6�t�Q_��B����Fz-�u��?�zU��7��y��'�~�7yY�j#/�.yY�W��6�d,'xwH:B��F�*����E�ӄje?�Q#�4�����u"`b^�V��(��0��r����Q���%�fK)��$�����z�KRŵf��5'j)8?��r���[oQUX��$��s͢U�Hp��E���Ur���4���@km��ޡ֠GE����9���s�HWW�
��ǽz�F\R�n�P�v�L/?A���=*�zB���x��9oz�8���=<��-�r�t�)u���jF��G��pp��/���E.����ʊ�X�#��Ѹ�F�u��I�z�zXZ5-�q2o�7{Quh�'��O]s�N:��aT}�T�kJp6~Jm��GA�^��{o[cG�����9mW*����Y�4T��1����霂+�$F/H5��&	_�3�,�T�����v�8	Q�y��l]�j�FFmf }0'Y\c�<~���x�Q���%�j�ʛ�8�:+}o�7��XR�g�k(�}����@��u]�>�4|���|H��)+�,�u��=��7bU��ֆ�@mJj�����q�&j��Gv��ԺPj��%o�n%��1�Q\��f]5;�fr̓B��:�B���X4'd��6�m\j�̅ZԪ��V��3���V��Yz�'g��k��f
d����N|��D�Jw̗k�V-'���kK�~1��u1d���`����~5R�u05�`����s\Q�ڃŪz$��J?7�B2ʺJU�if�,U�Kq�J�72���:��;��Q�$��{HD�lL�R�̭$kgެN~����XpZ�*s�0�ĳdX�FN�Gk��b���-���-������}�;c|Uh��w9+�zZu��h"V�OE��c��V�lc�9�.���^�������k����{��K��k�?�W�?�n��=cY.z�S7��NQ�����M{��F���׭r�����ݑ❩�Փ>�8kLc�F���^ZY�䃋�10ω�^����l64g��;謹`�g�!�V3�v]ET+/�x�n��bsII�r�hCo�lQmNq��a����a%��^�A���m��:�	sꝰ��t���|��2���&݀��9�2�z�9�'︡mL���=1՛f�H�qk�%��ȱ�c���q�w9G�1!"0"$�t7�����;'#+�r�iV���5b�wMq'�C� A��w��Ĥu��7��Y�أ��S�j�~Z�t��=,5��j�-�n��Js�1R5� V֔F�LS�������'B` W��L�x�n�����'�Θ�k%�)j3&z3z��VL�C:򲖺�g���,���H���Nc�����.�TT��+9�`ZQ�K���*9�B�}l*J]y0!�HK���;�sj�j�^k�u�'�%:Rͪ�#�(5���硘��e��;�\�_�)~p�spǱo��5��9��U�lf{�C�Վ�{H��t�ֻ$�AFkJ����br�ꏟYsˆ�YY�ݿ���~ޭ{����_`w��=0�YNc{��|����)���`�Ɏ_�e�gh`kJ��;Q�mp�*h�߮C얶�t�6�zq��9�����1m" ��g�{�N�qv���v�e�F!��q�۱"y��iDs�c����}UTtm�R*�+-J��u!_����1��b6�������������O?���o�����<�֬N�9�T��u%(p&M{m7������8�m$l7��k1o�K/&E{��0:Gk��
��3�er�y꒸�3�43��q�@�4餌��3G%�LI���������C���Wpո��t�����͖$I�,�ò�����K-�C� x���?��'D��Y�����r	_�Tea<0���gv[QT�{������r����f�r���D�QD�a0"v�<�7XN�4uF��G��s�]�,�a��3��؄�����0��ݔ�k�.�0!s��d�6�7�E�aF;�os�mJ��!��x��x����Y*�[A8�:w����A�6�)h3�;�9`�:	F��(����hmN���!�qs��e�f��D�hChD�-6tE���g���`G��\��l�U��2nD�tj���j���ϧ���LZ.<�7�Q+��P����O���3JJFT��ٴ6Le�����Cbk9H�0�]7[<�Y*�V�.�3��5�P�������tla�rX:����1�^�}'���q(;�Ӑ��о�sv���ș�c+9�ّ�w>K
����tO��^�ۼ]d�1�1L��0��Â��bF��_{2>��On��c�Rb6K���||9�J��P-F 9�_�,��MG>�e��TH�C�E��6$��}0J��H��YmJqTN���yA9��>?`�#�D|�g��;�ZWX�v�X�I1bb�Jc	�l�S�
�b�u��f���Tn�jľnI��(��MEv�.�xX��{��s?sh��S����^����Ϟ��`ju�VU�Py686��r�ũpN'T:�զȝÅx9����[�f�Sz78�/�&�ղ�1��l��Ư?�J{��p���P��%�	��C ^"�wR4(���l����,�[��t����I�Rv��Á��2ڐ��lm�0=Z�t�#�ﵫ�C�`�9����#"�4X���x�����2O��%3+�kY�<�P�)���Yt
NZi� L��}�Le��Y�p"c���߬���i�j��{T�k�cb��"��jrF��_��b7�A�
 4C_��6RA�VgAV`<?���i� ؤ�ٔ����a���6��Z��5�ua�y?F�ʆRt!uA�r�"���&h�ZPQ�����<���]��P���OI@�?��Ð�!b,�ʡ�{G5�-M&��6Ku�T	�S�I��G���ű|XU��Y����րgl�	7arg�sl�!.gk�G��~�NA�q�FW����I�������X����Nn��!�r8Q ޟS{�5X����ƙ�e�|� �m�:���;ym�8�������yV�!�r�9L��k �2h��ż����)6| ����ʆz�=�s�t�ْ@Z���1G�j��h�!��*�*��Ļ��#��}]ꊄF��]��c�B�V��Vj�x&���s�!/���Q���l
lu�|Tk�%�#�V��#!�m���y	<?=Үo3���G0��xE9��m1ӵ�$�8���eA%�$�U�f�a��xM�(L��ӪKbm7�m��L�'�U��T�0���Zk'�Ľ4�
�T#�kᵿ!����m�vc+�pT3 )%P^#!X}��n�J�V�����r��/������1�����Go�6���V�3���B���o�Qê��C����!F�!�5n����\�&$�[��jd���Ȃ;z(���y��o�@�l�`�|��X�a�t�X#23*m{]2�.%������0���b������2 ��CH,9[�Y���2���$>>y�{���F�Y<�R�	h��`�m��MYͥ|{G��x��d���#�<���r���'B�kߪ9��Ս[]Ms"X~SS����һ�I�͠X�!�N�@��J���H��G�������[����9vOI�s�_pg���"##���c�$�>P8�3Q�\i��@s��9�lpk3�f�2�����d�iI�#��FRFZyAe��wvR���Xo��O� ���°rV��,������"l����s�e��3��{ޯ��(S(,ؒ��,8~����D���Y����Ltڮ���9sQ��}"b�i�f#�kb0/�k!F��6g&��!
!e�5�uk+-M�7�SB{#�Amo��I�}�p]�NeSj)h��xך=i<=�8�DVE����9m��3��)h�Z5boy��]N�P�(�%�P��bS��\�߇5�A>�T2�J RK�u{'�L�����<���g�t���+���9�0���0�s��˼�b�\���������g��3��Wֺ%�b��&�����(�j�F�H�Z�K�n��^�<~��~yk;[y�ݴ��Zc
���1U>핪cSF��Vjm<>>��Bo�u�lxdM��'�N�.#imdGf���GԦ�FVs�k#���>�HH�����~#�;�S�&�q��� &$��饅���%}��f�]�V7� �h<�m��:��tmwL�m����`&�:!]i��Õ��%���1Su�X�1R5g��u
&�;W&s:�T}�T�g?��G����a@����C��[5ti�-2��CF&�N��Mے��m!�k�Y��;	r&�Ŝ�w������+�?���_���C�c�ڛ%c��f��j������<�8?d$)�(*�X;�{�@ӌE�m��0z���պ���Gg�q�xO�(�L����J��Q��ڇ��{�Q܄MR̐��v��y����:������]`�~���Ӻ�{��M��3v?��}Ԕ� pu���@����!�N��0Y�Q��|8��r�mT�3�UwP�!8�'��x��)3`i�{堾vD"�����9�E�H��¡R뎌�fm��gQ5��![ 1����3)/�/���l�7�k�68��F��ɤM��Z�8��Vr��(��R6���bB0�����D�{Ta+����� ���Y)�"<=^XN�V�`��Z-p�ބ��^�{o�38P!$n�Fi�ǧϟ��]���<`�t��'K��g���gIHİXoj������������G�T֯o���D�c���B�&#�gs���ڭQ��x&�X6�5���߾�ť����G�j�f8A��bX8��`�u���-�(E�����M�l�p�V��ƨ{M#26h803c���9�U������R�A�}�6G�96\�m���ё�F�N�IL���
ֲ�R&�lY?5cd������s�i�g��8|7/���,�gG���d)��[?)h�A��t���0
Q��u�V�ɨ{�5����Pw6�Tzx���0�ʘ��{wiQwnU;9�C�:X��ޯ{m��.�L�'��˯|~~���o��o�o��������`�w-�u��.���R$=���;KH�Ţ{6���dpd�56t��ϟIKFc0� �io��� �N~�Z���؇��0�!��W9��a�,����Hk$�,�;�iPH)��Q�	�@;� ���q�6��r:�{���N�vuv����n6�.I ]N�� �)�H��h����e�r�;E��y��t���=ɚ���m�F�s�N�����6����k��T���X"a$�Rl�n��@�<��ўqe%^�ۥАIO�.�<>���|���'����%���j��RM���&ք����e� �ZnV�	�%�{��a��8ؐ��J�
�b��    IDAT$�Y"�,��!r~t��mu1,�[�n	!�I��[�ݻ�$k��-q�*�N'��|����(�+�13S�Ds̋U��9�5VH��C�P�
����	io�7�ߕ�ϟ�<<�����u.��U�"	�^Meo���T� \�k�xy�j��w�9]N����q��Y�N�7��m&	l��(��4�S`Y���X����\Ng�uֺAJ����DR
�`�؜9�zb+7T!�̦j����xk[ K����3y[�`�CF�kxK�#_��l-��X�f�lP!m#=26w.��k���^&�AV�uj�o-*$C2,Sj��`1+yl�L������|8���(M������'�vf2�`�1ͮ�ḅ{7P�:�1���%;�i��H�YT�p��w���h�&��s���u��@�p�/���D[�+uNt�5��HZ��`��A���t��;_^.���?|���﨏gn������m+��+�V��,%���/OloBt���ݨ��$�L��Rh�wٚ�C���&��&i	�4�
d�!)JU�]u�U��10�F�9'|m��HM��JL�H�<�j��~ə�[�3�Q�d�4�.�W��B��L{ ��g�${0�?ޚ%b���{�J4$`+j#�P��%z�L�]��R_2"V�Ӯ�_㰣��@��=���;�ټ��&Ԁ����f)K�3,��3끎��%�s�ڏ�����v 2����1#����1E9�����V0�z
6��K�]��pyB���e}54gb?g�VC�:�u�6�͏6A����ҭR�:��=��\i}�9&2;0r�<Ӫr����b�pX�]@	���T3$I���2�Vu^R���
)�ty&�2o�_Y�_�a���K=�0��Qnt��@xRj�V9W.�;Y���������w<�����Ͽp����<c�	hS%
'J�,��(j�����ˊ�;��.���򕗷W.�D\2�m���@��
�P{�U�jxDͼ��~�<}~��r{�Z�&������X�g۬�r	FH���46|�$�j-b���#H!j��Y&�j��Ƣb���B���N���r�!�en�	�� �Ӵ��e�p�u��R�7-�V3r�6�귮��I�`G?�WwK�����8a)r̬ňJ!����s����$���?d"�B1ط�|�q��%˖T���>�Lǃ'�5�ҝ�m/6-�3�`s�1���N���m��u�(q��c�ؖ�8	RU	z�`��Wv?B��Io�*��G�s����׿L�\{g��V;�(��fk+<=��ӟ�˧�Vn�z�CR��b��v-�Zhו��2�l�nׯ��g�$&:��- %�I�[$�i��"��F� ���� `풃+�X���/���Κ?d�f�0�1T�D�+J��m�f�2�ZmνT��9��h�
!�6���}Q�z�(�hF�=����+m<����]!iY���)�u#��|D|�Z�d���$Z��2�N�MC��E%�H����:�Hi�#�$�}2fp{P)�:�g?��8:c���?�J�A�T}p���^Wyk����=)-�A�@�yy���5�Nc9�(
��9}V/������/?�7����e}{���Fh��9�8�.n׺�i�����$7bwm{C	R����nW�JΙ�t�z�x��+�2�l?���?��?���o����k-�,�P<�:�jc�<�z��}��@����n������K�կ|���I!�MuT������UE����M�ZY�:s������*i�MWգ���yV�^ot�ʷ�~AKA׫9b��U�#�32�P���j�e}���x~�p9?�B��ol^O=�4�P[&~�K;�#�4��0x1���ە�ϟyz<���B�m�:`2[���T�����@��u|��00i���:ؐaŻ�4
O���)e���|:���ҕ^�y@f[�ȆB���(E{��ӲCkGx��ꆮ���!��a��e�ӿt:�CՆ��f0���b$�LΙ[�~w���ۡ��N?%���u������$�}��l}
��֦�*����>Iy@�@��ݏ���r�1�9���y���2|�?�2�c|����!h�#��,�)Gj���:��������o��+�Z֊�kkH��QLV��]���iaK^�ˬj�\�wB�.jYM	Ѓ��=�7��1�h<��J�1���{��?@A(u�HY��u��9����{���!��\JJ��,�C�9��l}��jG���M,@�vӎ�u�� \�z-�%��Q���t"�ض��%��N����I�m	��l^kC�<��Bi;5׻1ޣڜ�.�×m�7�T��ujܗ�#'ALJ�C�nV������z��;����9_j͈�x� IvP��W�G�d6�����1r[�����\�ty&���yp.�	iS��Ѫ���H9��[%�q�8�h{-@�eYP	\o�+1ejSd����y���;Nb|������:KcoOrg0n����u�b��'���@�t-�fNKF4�B),�]S��q�:V�#Z��aU����B�!ok�!Lݮ+���t:�������+/?��C��by�q��qw��&흹r��x�+��J�����'^y����Emԡ�'�.�,z��'.|�Չk���)+'�Eٶw�m���n��Ƕ����{���QBV�6�d�pc�����8���D�"��d�񕸊���P�0rb�� q���&!L>°���޷�t�jd��|�0F���z�!�?3��2��<���̐���>6��׮d0!̭(U+�6+u�3�k^�/���wcī��Af+�(�$w��c��Ww8wC��襶a)ѻT�~�L��u�AΔ�TTrlB��Ht��G?KL�^ho_�b���ĈS�F'��rC$��ڄ[��&��BdM҅#�K�9=����9�6�Qa���@8eB�4Bs�'�}ks��AN�#'��urwF3��A����~m#!�'�뷯7%#�T3A����/�NB`{�3j�Os�2$+i>İ���#�G����~}�����	��f�KϾ�G��?"�wO~��=�#�����C����#S��dw��CJd����n�*�b�ǘ�v|&��8"b����[��Ֆ-��N�u��n@'�@:_L����ƞH1�{��B��3E�����I����*�c2ތڐ���Z"��eI,y�ڽ]?�%PC� B<Qk��v�	q���mE����_�������J�@P�8����:?���V�J�T��{$ʒ���Ј��7��F�}�Lm2"M�����9q�q�0A �ԡQ[�/�ÛV#����?��G���[����Znܮ+�6�Zͣ����$b���쯷����S>�{���"�����bo-���6c����L�ǚW�ڵv�ؤX�J�6��_ޑ�<>-�4n�m��¾aǵ+���g�J?԰�����{��2�1��_�V4�嶡���N�9���=��n�ʣ�ѱO֟�ޫm_���N�u�����ٟ�m�h�o2�0�`�b:H��EH)z���h�h0�r�����b����><��48���ӘK�%���?1줿���}��C��Mb���!HQt��}E��$k��K��Ih>�����A4Cjm���|��Z�Uʆ�319z}؟ɾ�bd-�m-t�HNTU{FR�������O�vEk�5����^^DWNQ	�����pS�m����p!xy'�D֣F�DW��4��
����Q=�>"lл����Ő�Z������2Z��J1F�)s?��Y�F����~��,��Hc6���'�yю���Q;yQrzv��Ze&a�8�l��� ?�r:r>v��\�[CEI�I�Y�$H!�5%w{);��sH� f��	DB���9������`c�h?
�}�!]�2�Y��"�$'��4��|�dR�p�Po$:� ňF��Qӑ���dZ*�7Z��1��uR�=8K��f��*�������w�|��rb{}�����ѣ)��n~a�r�l�l�Q�fmv]i�WL{Ɂ�ǅm�L�w�Z�i$�W�CV�8�L�:u-��M��KB��H:t)�*4j�:���S��o��/���|���ߨ[%��Z�94a,���C$�`�f���$Z+\�WZU�ϙ��GzXY��M�\_~��.��;j���U��DA���U�@N�N~��{�a<��қ����-���(�ea�A� `�8Vֳ^k�K�ݩ�f-!ð��򏤔�X�r�dfV��%�����Q	����&$Hw�+x���	a�;f�m��wZu��B�_;
>�l�ɸ.q�7#�Egm�|n�_�}���D�!�~��}�����������[8֣�����bm��v�P�3�H
�NQ��0`�����QkUT�!��l��o�f�`��O�
��7nk#��UZ3����O<��|���+�ۛ�y�S�d�:d�]�x[�Ѵ]o���4'���8�c��G����S��?k�s�8?�� �������+0v�Wk��A����e1}��5�d:{���:�]��?�H��6�N�n�f0>��u`W?�`���K�� �:��=P� u���Yd�>GCzԵ �;����A��!�8�/���{t߽N(����fɦ��]Iq'�R���7��?/��{��&�-��1�h���J�m�vEz1�J����l$��yp1�AE�O�쉃�V"1g������H��VMlkY��'.��������#)/;qu�w�
mu�֩�ћ4��J���x��f�wQ'�=�ޫ���5����'��]����QSM�����nd��t���_~���O����}}���?󰜦$�� *iD)��K+�E+)�ڸ^oT)|���|1g)��Y�E�^Gq��7��?J3Gc�>�9�2[]�����8e���)%9 BT�;����5k�È��'t9(C��y���a��Ǆ}j���۫xvl�ў6����`������uO�-�5�q_U�*��m6����g�c��x� �F�c[�)�)0t�9
"�όu�����j��"�)@��X�����b�7��yL�Sݯ�~�������7��3��qY��uܯ�����]�~x9���5b[�c�[��ڽRZ�Uw"�3�`��ef���7n׊��,��7�=�#��+�me���a��ݠ���j�پ5x_)Z���Dw���$�N3pb�w\�N�_�����ZU���͞������d��%��;�`�@�	�	���oc�Y�%:Y�Z/G���`�RF����6��[�J5q0���S�	�^Z�l��r@�ܴ�}r�C˲LG3����ahb����c9
�xA��/D���2h(���o����	 ^B�62����1}���9yڑ�n��ZV�"q$5`2ϊ+�Q�T2lU�;�Ǆt���v��g,�@���rZ8ga}1�L荭T�c1z��y��z'������]ń��S�$�Q�-�s�&p����1DZU�V�CJ�*��?P��J�Z�?�99t����K��"�/��3O�?�^i1�_oj�g�]Q�֟���x{y�tY���"��X^?��=G� �nm�5XF�=�^5Rk���P�V;J���i��8�hl�!�c��Z�v��GAw�s<(��7�I$FXٶ�M�9�%��l��U�.zW�7��9�ׅǿ�u������-��;:ϱ��2HJ�|<��i�f��p��w��x�w��k�J� u4�>��]��}���P-�1�:����xDo�׼�h�����(�=G/�1�<~-������%�������>݈gA��]��y�]�TV���˕�늰b����9/�.�����L�X�vۨ[!���|F{3d^��ͅN�
�y
9�il�}O�L�u������w�+ԚM����m��UXNy�B!�Cz���]��m��7�HG��cV4�1C�]���K@��NPk4���@$	�X#sRz���ή�[�>���s�>���%2��D���<c�W�h�e�"�-��F�5ǿ{7�E4v��|BD&1�R� Ot>Q
5Y犨��Q��G�j�w(���zc*<��O�%H���R=�:���fB����e�S�JJZ"!��XWC��u-�R�)�%P��΅����D��D�nY����~�v�,��I0ښ���J���]+�����4$$䠼�����z�"��~���[W����������'���o���<�B�$����`���,KF�ZP�I]y���V�<|~Dc"D3Z
��F���,\��I"J�+!$.�g�Rx���`N��#0�@Uw��y�d8!�y�3�`~��У�hJ�������Q��V��S��#�#�3�>�Y��d�z�^�!��a�����:�ޒZ�h8�����d�Zf@#>QK���#�=�ufo�M�/�L|�=�p/A�h�[�u��p��!��	199��m�D4<�W��C�~_k��J��r�x_����弣}�׏W��}�_��L�����S_��6��3"9�]Kq��3�X�7������ڔ����oN<<,���w���+��|�Y�1����SS���P�2)���ϡ�w�X��TADfr�}> ,1�LD*E}η�ѽ<d�y7���q �F�#0�=?��u�8����j�}� Dw4Sݔ��$��z%�L�f�SJe]iZ��i��Y�e��-Xѧ�uߓǵ�`�(����zi����˾�m��1�c�
�y�ﷻC��ج��6�A�~O9y�����8�7Ė&�ب��l��$I�s��uݸ�������������b(��!�q��x��u"�3`�&��Z��F��O��Lk���NZ`y8�{!4!&+7�W#=^҅Z:ۺB����jU�$��\�3/�e��2����Y�Lal�	��`��ڭ�q��n�>�g�=�N��G�1ҥ�����]��ң���[����Z)B����?�H������?Q�o\b�l~|��xZ�(���\΁��ޡ�B)J�
E�|y�v������c��?�ȵ���ӟ��V��
����6BL,Kr�/駽�uc	���k%����'$(��;Z*KJ�+�OuD��s��>X����pt���Q�U�^��K����C�k<��"���Y�ץG?�^K�9�:�xVb�O3��s<�Of5G��^�m ��B�H��Ԁ^��7m�nP���f2�D��N8��K���|R��% ��H�atyxPq2��JoJۜ�%m��)����=��V���0a���|O�n��x{��4�bD���N�]}mώB$�u:��7����;�y�d�Rw�0����6V  c=�h�L��b�ڐ���r@$�5КP���v��L���BJ�?~��C����-c�sMV���{)�����-s�AL��k�q���Yׁ	�`܊ �f�+���ZY�d)mz�u%	H� �7E;��:[���rds~K���h�h�l��[��A=�n�v�F�kx�U1XKcS�H�{;��
F`s2�`j{���=���w�Yvfw�Ӏ��	�!A���ҽc��,I%��i���>_}�cx�������Zg���}?!�b�	�i��iN~k�ln�**c�dDz�D�-(�ۍ��ڸtK��-�q�]������ၲ�}x�&��wD�9R1�f)�ꉘ;�����7>}~���L�7�f�|�a�a5�&������*�n��j��9/�/���?}��p�l�7��J
�bø���V�t,h�r���q[o�\�
��d����Ø�فt���ul
�`���9:�������3_�u�U���zv�V��w��#�=33��~��S�v��+��~���������Dw-a�g����D����%��x���[m<}zd�<������=UBP$��Q��e���k�T�=�-c�3u�~2([��	[��>�9�N\[����m=}߸$�0���d�"�Q}����\?"-�Hv�l�&�ʄ���ߐ�5�I�� �H�;��2�h���o6��S72V��,Q����輕�$$sr��0.n蝗�A����    IDAT��I"$��ǭGK#8��J�;�4j3�S#��Z��c϶��n�gf�%W�Sۛ�Q��X�/s�a�3������3���T;co��l�鬊�h����i~���V�A��(l��k�r�X�p�7�3.u%�dħާQ�4���e�C���8M���nZ-���&q'�Z7��u�3��8��!����0���`p�RZA�^F��'2���=#�4|�3oC���q���a'�^�ξ���v�^�z�;�&���`�a�Z�ҍ�-n���A�e'��%���f�(����`鼽�k:��]I��s̀�k�>V�W�l��RJ&��>?}�l�>�/�bk>Q�fȡ�E��sF�u�T�&�M�.�͛�Bp�/�Z��,S�\�|��1����.:���l��~�g;Z�)�ZXNg�e!'��
]I�H7�+I��p��s�)�,��f0!��6����`���Uc�t�G�	�Q�U��s��Y�]鵑�|�-����__x�<	����[��^��Ն�e�����;�$��|�����Q�-�qm3�2\�`�t�����wd���z�Мy|~��N�+��A"��?�3��]������gYz�� ����*g2I"/t�3eI"9�X�HA�{;D�|x_���3��<��ؐ�9�w���0�A�vG�4��ݟ���Mb����g�DF����Yk���i��.�@�τ�8~���+1'��4��g��bZ��L�`�Xrk��]]�{G$�/�n� �(2�َ�c�l���|]\ip	�5���������;̯�\�5b��Cj5Qmʲ,ܶ��Ҫi3�i����e��%��U��*A�_�_׈�FU�s��=���S�^��LUd�`�3�1४����$�V�\u�������n�h�����F�{3"���A!�*����9A�퇝ѵ���3����^�ׅS^�V�<8? �H]]�  @߿a<��^�*�L���:�r�GX~�hZ���}T��¾�K�k$�Y���׬���S�Mq>@�Η:Q��������^��2a���������^��k�q^N�[x����a��啯������LB<@��D�q������V����FP{	  �ħ�.���e��W���I.�����Ȯ�C���%��޹����Lk�׫�MF��^���>��l���/�Zk2Ѷ������o[�g�Z��<��YO��F:������(R_}�������E���F�B�HjX~���6\������UDx8?�^7~��|���6"|�O�D��T7�Zw�������t:APޮ］���Ͽr>�����d�`���-��V��p�Y�f���rZ��*���p"??qZ�z���/�/۾�F	a|^��Imc��Gtg������:��M�Z#��ǽ;���/���A�k��6�=:��[��5�����ĸ�����됗9io���+b7�{@ћ��6y���k8����b:����3ه���C����!֨VO<>�=(�A2���GC%b`K����R
1V����6�5�9�H��ƼJ'����v��&Fܳ1A�@U�Ho���BV6�p�������w��<b�l����INRӭ�e���?]��x˲��j���9*7���m ��l$�pª���X��`������h� %��
�p�vV/ըrzx�[�c���n?ND����|2����}��y���N�ϢO�I��0�p�Κ�0�f�0���U���T����`�n��;_1g�@o�{k׵��kCc2��d��O����f���A"v�B��y����b�$�T���D/��	Z|t�F49WB��aa�����u]A�eݭ{�݃"\�v��ɘ�>�z��6HRi���j�4�RU�KR�Կ�H��J��h3v������=Ϩ��㐢4��H2���F�]tv��S��ps!�#G����_~���g~����������������#�wX-D!�E�CY�Ғ�n�_��\�dI�r�Q����鬆�!�����;,Փ�m7�V���(��(*d}��Z�+��vPN�h��^>@:D`gzkP�j,�rY(�����_џ����¡�[}]j��gVÝ!<:�;"B�23$a;��߷�Hi���A��Z��ѻ�RӾ>���	Q�wNN���څ�;2�ӴڨIsZF,��GpG��+��uOC�3
�����['<�.��ZvV=:`����s*�����;��C&��)Z�2�q��3�y��47P��8#(����S�k%J��a�i�����y�~�*F
�.��
�L\�H)��I�i��v�b����B������w��?G��!��;7GQRJ��8P$�j^��hm�ᔧ���X_�۔o���q����s6�|��g��8��7k��F����)-���r8��n��"���D[� �Uֻ�0�a�析��6A3��2��F,�~�Xy.��c ��(B�*KL� 6�v��xpU�k��aذqԿ��7>ܨR���K����<�U �m�Sz���3�6�v;���c�ja��})6L�SI�>0����l���eA���M|ʥ�k�Ɏ3�H��/�%�M͡�à��1[�ڍ����Ҫ�Q)$Z�.kl���Y���QK!���E�� ��B�C���ԑ��LAМ����Q��xGֿ�3j�'r�JrSʶ�ӏ���~����o7�bSԬ>b3����4��Z���@��^���tJ,�رe�h݈6ֺ00����na�ť4B�콭�A� -/6H���Z����d��9�Ȟ千�"�t^���k�\�;�/_�[�tna�����89Aj�Uv�������Y�/Af���,}�u�kǫ�6K�{�g>��N��z�����5���p5kw\OW%�Ӥl�Z��0�"wJ^{f=�F'*`�;�`d���3�%���#u5����q�J"�41i���i��8���=�m('K{��[��l�AN�4�;5쥶��Fk#7�s�b<G.�<�ǅ�ܱ�T��>�ӷzSn��ֆH��/?S��0	b)(�tD;װ�e����R
�2嬏�mH���v��Ht���P��5c4SGi)�Uϰ�fS�؝��q�?��~l3;��"�69L۶�sO��&?S��Ύ�֨�fA�����@Wb���\�eڞ)��{�?h�����sj�'�h���j�Nc�`�O��έ}k�q��}��P�}F��⼗�*9��e�L�uz+N��D5R$X�BZ��_o�pqG_�������N����\�� ��]�= j��9���E|ts���9/3��i��1�r�i�k���-˞-�K���I�Ր�$$i�!d=@�hC�<h��W�SL�٣�{��V������il���![�zP:��|o{bw�^���!U�S>�믯�T�� >?��VL���J�3��c!�\cX%�-�[��ן�r>/<<�Y�b�\[��<�#�$b���Z{UJ#������t"/��W�Ĝ����\���}�}�t��L5s��)M��V7+Ah�QK�Xi��}fXx��g*b��J��Qug�Ў2���~9 �Q�7�]6�$DuE0'Z���&B��X�Bpy�N\N��n̋G-�4	ʽ�aY&�H�FC�9�4�&J������Yl0".ż��G�02����T� B��=Tw4�`5�#
��I�\������s98�Ee�o�޾�lzyd��ܣ��KqA�`�(�x����GT;����,��}��κ6ҡ5�9+�J54oIg���t�:v�z��B�2,��f.��l�J"Y�hO�:5�[��1O�����ԞY�W��FJYm�e��;�@ݶn#X3�Y����zQ��[��<g+MY��ȠBo��ֆRg@�u`��0�g�:kԣ�t��K+����!�q�TJ��:;DDLR{��;ik|Oș�d�����n$�^����"u�h�B�ɘ���5=��y^V�����4u^�)���n7N1Y_	Uk\oW�yr}"6V���^lVAU%���4���f�坓ٱx2M�L�ցa�Ķ��Q�ּ��B�󬝜")ڌ��6p�	\
؉��9'����R�)�FL�6@,�A:6�3��D����;����F�jD7=��.ku>�mL���&d#1�Z��ۭ�׿��?��|��?�O��O\�!���% ��@����.�%Qk�VV���E���J!��%&na3pq�z���y?������9/k{�B̰��(��}�����жAh2���G�@�t]	�衡��SK·0��L���Уպ��d����#z��^�;�U��d�0��!R�Ü~^>�jR��$Z�S�����աe���3�p�D(������j(e�Q��b�1�LQ�]M�p�66S=��y����u�C��w�߫��Z=���~#�0z��.���g�2?{8i�^�����OZ�ȪF���=^f�=qØƔ�v1e�R���ӗ'BR���ϰ^I!�$�4D��@�UM�3ҺO��H�M7�����<�P�ol/?C/���I��5�~eY��i�氆������׶��e5�Pk�t6������|��qi�;�Ү%�ĭW#�a��:	2��w'G�����>���Ge����9	37�큅H���a��wz980��!�e���U�-˂4�>�� �mx˲x7F��in�F��n�{H��Ό>i%��6r�7J�{��׽�6�Y�1��O�e�^ۼf���6r�lj6o����v���˅�9���t���#����%�l��8m�%�}�1@JP7z�R׫�L�	�]Ap:��Z�Փ���m#ˠwg��ɫ'5~�G���j�v{'�|X[3E�~N���ڶ�x�<��2ݕ�ɞҴ�j3����H�g>.�����]_����oj<��72MZ?x��,��x���2��x��o>�W~�翐_7�I��N["[P���x�βN3��PG�&����Q�jᶮ<������i�喻~�{�CD<
����5�mv���OG�;��k���9ϻϐ���1�5�߼?B�{����3Q��~��qݎ���>�&+����ƻ��l��q����>�����?=���T�ϻ�\�S>L���k<���=4���a�!��{�G�q�����b�!����ܴ�c"���J/I��pjgm7�ϴy}Y}ȐA�M�Z�ߞ����?��t��忠?��)�������˲p�^)�F&�Y�E)e������̈���gdJL� [��W�ca:�a���3ݏ�������<y��d`��}ODf?����g�[{��(�$C�B?��k0+��؃���ẏ{k�ϭ��ڏ\��a?�����"=���L~o-��ͣ��?�O;�x|�]{��?7��du��B��s�RʨD��>%1��"b×���7��I�#9z�NFDfuUW�����d�+���.��J�Ƥ���~eefIw@? �;�=˶�̌�8����"'�0��J�aC�U��:s���)��� C���:�C��j�prb���o��������?�#菲'(�Ɯ;lh۠Ù�Z�������ݰRN���l�۲`΄RuY1���~Ǒ��!�Q�.�q>]p:���� ju�юQ� d(&�����pfz#OP6�.��~�5��ѭc8��ѡ��y�܌c��Z��3������g�����Ľ��Q�B[����$Pk"�{B�Vp���?ˤ~4f��֡��x�ج���5r�V��� +����I���8�Z�c�}����Vm��p��lM�8����P�XS�m]�{��iB�Q��� �mi 3�|����O�p�rF��7���_W�p �S;�\���������%��(��L��3��qo�� �vʢ��g����wN�I@Tپ�ڪh�Kt����v��wF~�Ϩ���U���#��+���<^4|O⨣�&�O���V2MD��֐,����q~e(��@�igI{�GTk|t~�\cH&>���A��ӥTG���(q��z�sۃ���(�} ����gu<�R����mö� �*g]��)a�f0*���ƒ����`�6�0�nX{ޚZEMT5�L�Q�YJT�#h��`����{
x~NS��ЍZ�(Q�G&z� �!�!�B6����mx:}E�Nx�l�v{�*�i�0��V�#?��K_3`ki�������	e�P�Yy<�07h�	�%Z�00��ܺe�֛�n��U��ᐏ�
��F���;yd�RN�G�pc��b6�f�3�}�����zw���X�\�X�*o�
�}&���?HdM_�
�q=���a�MXb|{�PB ��6�w�{c OG��������#a��,�R[gcdj!7�@f�)-i��Z2���i��>�������~y���i:!M��VlLxN��V=�b  !��s�A�B�#�̲�?T"ɪb�Z�΅��ԅ�q����u���f�}����Q���~��#�Ѹ�������vE�Bx	��USj��Q�y�z'JS��,�֚[�eTЛA��V�9Z��h~��5���C�^�ň�l}|�]���Q�]\�����W��8D"r�垙M��`���*�i��0ό)SCYX��cĪ�Zdb�f��Y;��e5p"ū���N��y�L�S���g��9��5��>���k���@ͭ9n\��ѡtMQH�� ���u���oЧ.���~��|"��tƶ���<9x=�(��8�q��5�|Ze\��� �e��];�[���n!���X�i
Qk��AS$f<&�a�D���[獑��U<۲iվ������ck�>p���,��XU}�kZ�x�g��ܻ�,��<)�x�{�b0�v����C��w,o�F���]7�=���~��1�"�߭�jS8��ű3���R
��w(N������]�[uF� 'B�
-�x��b&��OO�*(�"M	\x��ȉ��{0��w)<<�<a�\�`/��: �^)?z�>��`;$]�at+�/-5���Ɵ��x�#-�C��ӣ�Q�F�~�b��d�G�K������VɕA�;����c��Q�
�6��g��t˚Ѝ��;h�A�M���P;_����z^Q����?�1Eu- !��L�[�,�wb<=Y�{���K0'@�P�1[�t���???�1U��P
��xE�������ڽűf�O&�:S"�B��p7|��p�S�_̢t ˌ4���%1��߰-+>�����j���7�`<_θ֡�]UϜ%��JwL��[�"�T��'��g�uEQ5Kap}�Dx���w�QC�{�b��-%�!��)��D�}�Hc���'���"���[7(<<�
�r���5j�v�C�-���������P&?b�9�HS^h7�dI�.��D�y|`T�ԟw�^��y�ix4�G�=*��gc�w�$���H&��Z"�.8[�O�~��@���%6�u������:�Q��A)�4e\J�֠�R�ǚ�h5�޾-�#c��HO��^���Θ9^��c,yh}|F��G4�>7�~��bT����$��>��b�S��7�T����of�K��a�hO��������l��o�`�I����3���J�u]�Ղ�oo�]6�N���>�c���)kOPb\�!�<g��YʆRW�ց��2eJ�sv�AZ���O��\�x_߰m7$�%��������% = �Z��L"m8���h��"_7�V��<��~�O�;����˿�?������̭��^ӳ�2yqKjM�D�R����P��B��$��:{�H�����Q�[�a~o�U**�t/���wV������ק2�|w�Ff��1�����|U� g������3B~�(G��{Vܨ >��8�#��4⑎c�c��~��>��b�4��u����h��Ý�Q���8�[�VJ�}��b`.O��8]���6����nn5�f��<Ns�<%�T�T|�<���Tf��-��9�K�����.R�����}�.��\�:�UN�G�n�c{!{�M#��އBx'�Z�H�`�P    IDAT�����h0~����E��8���F9�c��Mr>�u��c=���L��0�y��k<����h��d�������X��b�@7W����e�m�S��#)/�ܐ���6�&��X��h��2�t�P��z�Z�UT��bM�y�vFr��?lVv�DXo7��͠�a�Wɛp)��<�jy���v�y��B���1�Gl�h��0�']���v�g�ׂ��W��	?�����W�o�x�1[���3��|ѵI�� +qIԱ�Mc꙾�Кq�F���H�@ih4�@|�J*���"�>�/,�xf�n����a�q�ٺ�wн�?
��"z�.���edh#��H�=A�ޯ����m�E\�#e���	1٭ogZ�_C���vM���'���7�9&5������Q��W/�
]k֛���8�=#�JǺ�jhV��
ʊ�4!�Z!�u�Q<�	�Yv{>[[�e�!W湡y�������ʐ�(��9�|/��w;{���M��y��?�I��t�KW�43*q�w&޹ϙ:�����g�}`$4��0~v�4����>�g�E���ﶍ�����p�u��1$��G���xT�8]���T�� �j�)u)J8�����V�{|~�àX�)D�t¦��
~:���		d[�P+ѵ;��
�ac(PCtBk�c�HL��_`��i2�ݡ%uc����<�i�ؼ��\I��fdH��{�����o;�LU�����|����<cNg�}{������?�	_��,�7෥/<����
�[j�C��|�����s��y�|>a��!^�#r�Q�U��k�Z�ca뾤δ�������i�-����?Ҷc����,Gk�hmƾ�ew����h��?�ne�]��hA���g{����h���Y�q|�}&�� ���x���c|�ޜGk�h��ϸe%��E�A��u��E��,�������v�����V ��"�!�t���RV,�w��!1C��ۺ`�O)c���`k�<a+R��&�lbR���������-0���?h6����1��W���߯�sLtP�
Y�51$�F%��4������3���<�O���<�]�r(?m��0*������U��a8$�q0>�y�V;t�x��}k1�gr�V��f=rx�=OA��yϧ����������!"ޞ��<�m3\
?�O�_noXU���������Ox���9!gC�3�8��u�D�mYfW��H�%��PIk'�Ći\�bMb=[x@^�	��g3Ζ����\�ND&�l�X���d:.�}:��4���M:�}���/���?������������gLH��j�Rp��i�!UA��IQ���9[B�X���j�r>�����&�ю�,��R��`#p�)'�)l0�U��Ǔ���u��>�eV�xzz�z���3Ax�Vp����A�%��_�0���=O6�<k�w|F�K����"g=�-?0J���ZGAwdlq�b��H #˲�F0� u��a�����LR� o�6B��e杠�1F�'M{��;FPz�o���E	�y� ���iw���9��n�RBk
B��/A*��ͳ�m0%��*�u][&x[#�5u����
�UQn&�O���m{���}��i��n(�����Ԃ�vBUkg\��2������yB%�LV�^����e-x��=�Ɏ���S2/HRO��v�m�pK�#��
)�LJ�]kԑ��ڳf��xX)֟;���-G�^��l�2�\��Ͽ[l���Z���7�Y"˅X���+)�^�4Z[��6�b��0r�w�}��AT�ڀÌ-$nVx���(ۆm����5=��uHK)a�g+��C#���*O���D�ݶ2?!�˝��V��(�s��E��!>N�	˲���'�%���ն7A͖��Е�JV�;3���eG�ڤ�~����$���Ys�H��ॼB�����T����o�@�7�TLd�"��^�T<�����u[��f��)g,}���h��Fa/�n�O9AQA�pEǺoB_;�z�ﮝ�G ���M9�|>cY����p��ϟ� E�n�����f��a-g�\-O ���HQ<Y#x]7\��ۢ���u��BJ�H{W���{w�ҝ �����k�X���?���Ԅ���>G�8�7���b���ނ�4A��i[ND���M靠$��4aLC��zŽ/��X�#�8J��K��	�!Gdt�?���ŗ{��w��>�Y�6ڹ-G�M�rPF�kL����ya�6����5aW\E�b�����"��f�~�8�Zb����f��e(X�#�}��'�%��
)��EP��@V�>0J�Ԋ{yǧ/�AS����R^����b�Nx����\]Q�΄Uf$� ����ȧ�@�Ȝ Jr>8��5��	&䁞2'l��F�� VX$� �!�-,gۧL��	��!AÂ��k�L>NA%A�0'/x�%��e �h���ֵy��}p�u	���4Ё[�s��9#'�xS%��x[r��g`ʉ�᩵���E��J/	32R:{x��(��ɀ�R%�r�Faq�E0s�iNͫ,���mk�����C8���TՔ����u�����k�(J�`������^n�x,,���f�\_�lmKmH���������S>!c��DJۏ�S�������xH�C�=[�l� "1N�|����z@s�E<@a^�'}p=t����i�X���� �w��Y������c���7,�E+N�8M3n��t(�SS� I�,�LU�n�g�xK�X�❂�I��ԑ�
v����bN����b�z�v��Ȳ�K)X���>
�х�RO�0B�z*�`VH/�	?l	Wm^&C�u�F%��W�P[��0�IM+�^��Ƚ�4�[h(�|��/A���&ߗp�h�ԑիĻύ���zp��� RG�:
z"��废��8���NA��=4��
M�v�����$�?⟪YǵHc޵V��C��*����ļr9Y"����	uٰ-��"1�E5Y���6�	�R���/���O߰Vã��|�9M(ۆ�����;�Y��}�Ή�MO��nb�lu��Y����XTRQd���iF�7�!�4O����o�d�T�rr%���6He�`�]�{E[>��{6���A��m�ߟ�����^�X�򯯦��Ihʬ۩u�r�MF@Y���������p�K)E/��b�W���9�Qk�K�r���Y�Wj�@klD�[�3#�w���0�"1'i8�4e�4�{~5�~>�����ij�6N[1o�&k�j��B�6\�E�3�Ɇ"�IM�� ,���9JO�x��#e4тW���UVXٽ%�4͘g�v^|��b��(�{|� Ӓ�b_�}��8��+S"#��≞�����Vp}{��@>_���_��������S���
@;]���X�������3f�o(7���|�`�w¹[�V50�5M�tμcr����.^�Oi�Cv�>�!��C��	Y��{�D�z0��U�P��<!�u[��7s�eƩV\г��G�|���P�ink:��=�Հ�I_�P���S���`�P$�ܗ����1��Ϣ�����\��oއ �	���y�{���_b���y'�F���eF$����bJ�5)�䥜3ʺ�v�",GF����ܦ)1>�`�V�ui�yf��ҹ!�?����"^��������?�_�|A҂o?�����/�~mΞ\Kd����;F'�c�`�����#|�Z��ѭ,��ɘ��i&OXTq�C���3ji�22��Г�Hݣ'��U���D�5��V7��z`��֝��Tr4����c�g*���G��:0�z����EX,�\���c�B��˚�(˭�L5O�AªZ������c�wE����VC�'u��9`��%Vm�P�:}�g7��|N���g�P�6df�\�P�%o� Qv� 0o���`����˚�Z��U��eY1A[�<t�	�<��=�S�1�qDR����� 
������=����^?�d�*����pdq�\��nՁ ��vC�&�s�*���;��'Pf\>¶mx��7��yrT!�� ���o�j,Cۂ+.�>�������?)Y�`���o��"p׮
ΐ��
a�6O����#30�cE���m�,��;&�PE���œ[mJ�$ �����e �i2W�3i�m}��\��@*����Ŝ	�DH)#q�1Im��
��˚G��Iw�63�Xs���d��COw�5i�E�(�Lk�P=����Yo�	$���i����۠o���`��FL��3�N5��Udv�7fT!L';�y��3н� [W8Ƶ-�`>� �I����D�U-�9�R�IP�qb`�����1X*خW�X�Y����T�>'�P'լحVc����L��yƧ����ח߰�����NV����L�@��G����]n˨P��x�(�x�{KvEW2�-�t:�gh��]8G����.3�S��}M�RU��)SihDd X&<7�+/􀡏9�X���';�?�A��u �����ORO�K�J 7�^J�-���`��i�sac�gC��m��@�����A��B��p�!�2�X9M����njFv���<���"<��i���/ϗ	��	˺zn�y j
�+��\q(-_@T1qF:��nX�Z��l�s:M��`������"�M�%�)����¿{m����㪊�2D�2(�XI�m�jX������oĽ���V�;���ų4r`�wS��z�{���;n�H�쵺�_���9���g|���nx_�/}��0�8�j�H�Sǣ&2��!���]�/�u�^�Mh$�j~��r��h����~/�zŝ6mkʃٻ��D�6�v�wt�փ�e�P��(���!�����,��K�]�i�S�"I��UP��9 �ʌM���!�ld�m<"ؖ��Ƌ��.�12�+Ӑ�'^7.�����Q ĺMя��`�99�6�G��h���&ޟ�	�u�O@�R�׷7l���!��_� (��1#���Ko �D��B�Z�e��ar���n3۔&�T���\���lf���PϠ�%{��)
&�RŴ]���oo� �<B�����ځ2!���!B�h���V�ؘ��ܹR���2���k �h_�Aǔ��]wk���81EM���uxE*(BC������emkAq�$P��@u�0Xڑ��!Z!�=ᣄ�*�*��C��2O4#�����r�U���ĂD�`�3�Z�:1�����f" Gba�2�2�D pRL�;)%�zgv%���<�J�{(���w�uzL���~�Q7z�JK����ё[�)%�9��b�6ɺ*Z���z��<�[R�T��y81�0�&\.Դ�v��������4�p_�%ԫ���,G�]�Τ��<�O8��r��ʾ!���\@s�������9�MG&t��>�r�e1ANF�ۺ@����w�������oXD�7װ85�$C8U�O�g�{i�� Y{���)���~?8�N�/z7W�\;���D$W�$�Śk�?Ce/prT��`�r��b(���.��:"�_�:nڳ<����p�!�L�A�8��͘�GVғ��)T' �s?١��V���V�#o��S|�<(|O_`^�O�Ǔ���v�Sl-�}�ǜ뺵ܔ�e�w����ucm�,��SO��	Ĭ�/��v�,��� ��^i&o=9�a��="Q�܍k^���!$��)c��&.b��L	��@�*���^�9e�U���@���[�~@'c�|��0)��W�l�D�X�(;�F��*=��-3�4,���+��bw�I�n�@���Q�Y�F�^�Ϟ�K�aYq$Q1C6��@Gae	�Q��^�6���1D���F	��⥑���\4E���SS²����*�����)y�&�ߦ	e������Q�)SlB��#GB)�Z��	�}<& ��ɒ��R!>~��'�ӡ���I��F�:v+�Xk1m����mXw߷ZQ��JE]m�k̿8̒(�l��r/c�օN3!Ô�$ /�
>��kԔ>����L
�8�(�o6/�yS<��t���G<��G�O*A�La�f�߿zӐ�]��|g�J�8�NP���y�0M=�\�䄷�7�����H���+�B�Y)��QC����41��������-T�o0�����4�D�������Y� LH(��E5���Rs�޺�eu�>A�P��B�\cY���W=ɠD�H0~����.��ˀ�!���C�20�YU�P�ncd"'p�R�V�8h�n��t�՘2���` �Ѷ�m��h�ʁxOf��ehS�`��a �
h�u�>�;/�h��������u�Ҕ
���=��x4V�YԤ��&�[��%�A
ST7�>�jD�!n���E�sB����٬�)�ml[�	y�$����E?�J�L9K�Q(Œ��c��y�|��m�ۺ�}V�������|��dess����j� ��^x2��`��Z-���Y��!5E�x��B	��{Ќg�bU	
�PJdp�:���aoE�c�����2Z�$=�
UkD%�\��N���6E���@ ʖ'P+R��m$��)e�D���|�+�d�c%L��
���w�S����]�*�Tf�
)5# ��l����
FBN�4���o����!��&��RB���W/;~��qUKЌRC�!�2�C���y�����;� FN�ǵULjr�� �gLj�Jau�&�SJȓ��H��ٍ��j5��`�[����PC���nmq��:-АU	 qM3h:A�����
� /[Ŭ�R6�s��'"n1����O�H.ك��`���ϔR�?ew��k/9�i2"�������?�\>������?�����?�T����,�y�l��5;�����gs��% �[�L��eG�'���ws4�!���
��yR :�)�[ת:�<A��i�c.���R�JP0�j17�L	k�sxM��4
T��+9��!Զ�꜆29�ņZ�����豤����a�wU���`ϥ	U��*��%;��V�B(�������6GN#@���G�[��h h�֝�w��.!�=�,��� ��۴k��y.! �@4���W�Z�s������A	L�+�l)��u�����g��ī;0B�8�8�@m�����3H2Hk���)��;ݔ����.l�W��^+	�:�\*�zÏ�7���!�����Ni«�������Sμ?wN@�f�[\~�{�_��� 	U-DݲB6����Pyq�+�� ���a�Lp�p���~���r�%��	�c(��x�^AG <��s]�e��/c&Ʀ�	@�Y���<������Ah8y��w9�(c7��1��2&FW��#��Ϙ+K�	�2�*
��p��\[��E#i��M6�@W��[BS&��.��DZ�a!`�V�M��C����窊�2�1�UQ�"͌|�����P�(��ʧ��Q�TKf���3<�p\0V��0������>ˊ�ނ��N���x��������k:#3��l6	r���}`�j��=U��f? <T���>��F���VWj%)�
טZF��7�*>�(���׭bN3.!(��|q�:�ع~wl`��`�-�6�|�]�މh?K�=Ӳi���ۧi��8�iI.g�kq�)\	�^um��A����1|b��H���Yd�H���i������eI��j8�+H��F���&�Y�/��@��lZ�֧I�1x	�4�؜���c�Bڅd�MN{��W0�8� ��~	�L�BbMQ���EC���1��(þ:�*5�a�\�&`���<"��Oc��D�3F�Vcp�E�$ȉqr���N�%+���P�~]��x?��9�lm%<<�Y���4�8CH���1<Qt�;��Q��Ky\_�FK�N��xT��HKV�~W����x�z�^ۃ��v椏G�1�}���C��@a�ژ��L��Y����:9����3
�=�6�6$P�z,Dܚ\F��  �IDAT- �E({5�B�h���0��K�uf�wY%"��a �ʦ�	&�l���,����7K>��\T��@@�9C��3?�A��΂挚�5l[�) �\�e7P�
�'!h2�p����Qx���_ΓR��#�<6�J��-O�����u�pd܍��Dd��]�s�ܠN�6:0�n-v��Ta֯=�]c��}]��T�~�g<�E���WR\҄T��<>�c	�	{ws���@'l��+���R#'���� ��
j���dnF�1jB�q(Z��^y9��Q��jl�B͙8��XN8�Ćy��2�^i���wc˺+�(h3h���7K@1�>4�ZA ��u5��nN�>��7�X�f���n!k;�A8w�7���L�J�Ad9�:��DDK����v�Ib|�"�^51l�{�ks�z4L��p�P e�"��c�*$�x<OV�TE<.Z�<���B8	���i��ۊ����g�цӔ�]V��
|�zd<:%sG�C�4���c�1?�����)�q�}��b�Ċ9�/�p�#��U�;��Gz<��68���ϴm�\�=_�g(�Pt��iw��M�VA�<]�P���x�"�5��Ce����^�Q�Ru�k�p�>�"'\T��F�S�6�2a�d�DX6���ЧW*\��X{e���w���JQ(�ܕ��7g�Q���j��;���6�ו5g"��z�L�7Ο��:�;SF�'���n=��c�U7˛"Af���@V!(��$�����h��ᆌs�1���׾y{"r��ܭ(����Z��C\�dI�(*~���4czzƪ��톥n8��7l��	���Hz�E�\�Q��V�}��l.��0�\m�ĀE,��ȁ�T�QE�[�l�{co�����k|�6�Bu&�;暧=���9YC�wa2��Y:s�-'��?&-����Wv�ʐ�2�gk{)�0����� я=��`��X��hBޘ�P/M��`ަ֖��
D�)��.zDfL�{v�p��ؕ[���.�ݸU�i�hW�y�[~Gܓ��uM��f S6����LUI�q�m�U*�j^*���-�$�
Xo�ӄ���Qkqk���,A�֣�M,@(��y�Ϡ?ZS��0�χ}��l��fl[hw�P4��H�w��sC�+ ����~�tT��5d��P0R���Rx>Bq=��<y�Wc.K4=8?$��W�1o^/m�.(Z�,n��0��ڞ�#�A�+*NdȂ�<#V�&(Ȝ��䲊�2��z�0k�0,Y~A<[]ЗemF_���&T����H��0`r��`�9����F��ذ���4A��`��	R7H��L"ji(�-��5f�����!�9�z�߸I{"���Li �������� �+�9�Tv.t`1	*
�
4%|��>��=^^_��_�"XK�n�CJ"{H �}�QB��˔��1�>��=�M��*��%���Q"����6\����N��;�(������]3������3���@�[2Ҁ�&����rʸƑ�N�$���2�4���ܫ��R�
�q�C��~���qӏNׇ�$�u'�&�,I�JkH�b�.4[y�0�ȄQ�q��F"���9m��9�Tq���)��\��X3 ū�~���1%hN&�iF �YY����
���
-��A������5k0~�;��"ޯ�6X��G|'�gJ?R� ����v>�TuX�v�DH�cgG:���Y)�*������L��?��+ ��ǽr��ų�O�=��I�����a쨅q��=0�qf���ĵ���{�ΘXED��&��ھ��}�����-}� ����s�1ި>�u~��Y����(afF���	P6ܨ4���H�� �������z����c{�]�W���V��e�<��U�l�b�+V�Pd>�@�[ʘ"{�454�m�����[3�Ljw���[ܶ����'# QGs��+ޯ���໯����	x:�T�-k�4=����\E�Q+��Y��K V��ś노�.Vs��У�=���	A5�mt�vd$�����k�nws�\ss�&�C�-#<�=E���h �����9�&?���P�/"��� 3�i����.�s�
�4{͕*�q|T�0��j��;>C��cHH���}n?
́�f���IDݺn�����\�Z�*j9��{5�pO:g<}�����/Plxbë'b��L9NS�v��(K�d���9��{�.����u��b���u	��Ev�< ��OӾ���'v
ذ�ad�r�hWx���>���t����۹�n��(��d��GA_x��x_��ᑈ��M顴6�'��=q�!`��t��"����sl�Ͼ�١}k�(d�p�	��n��`��g�	x�\��c�F��$�i�M�*�g��qef��*��8L�  iI��� �����X>�������=2M .�(cN�@��3�����'��mJ��n90�A�v��dD�fY�J=>c�O�e� ���6�	_2��`����}k� ��N��/Ӫ��$�1�f�:���D��A]D����%^�<�(��ql@C�S���8\���������;�E�����VT�8DP���1 �R�al#S���Å��PWϦ�A-㨉vs��XYN0Y�\�1��c��s͏�zI�=�[jX�Q(Ž3��\��cc׿�ʎ[luPI-�����&��^�cډ�\���J��Yם3���	q�<��,���2_�������?�_ޯ������G��O�'�<Y5��DK�#�z��q�Ci�є�(3�<���r|�z�@�1���=�{�0�ȃFC�d�I�Ù�>wf�Ze7�ݝ��S��$����#�	 0�5�L�*X����}�����#�{�)����{�!��\X,=u%B��O;�����L/	�jJ���0O�5VU�K���^�j-ho7loW�Z�$��j8%x���`j%ù¿"��7��x�CV)Y�H1�B$�)�^=P6AEE�,��A�Į�L�������K0Q(D�3;ǣn�_�Fh�C�Ӟ��B(��YЊ:�4
Ҵs�Mq9�1C���Z�j�i�P���m�g���5z��Ǔ���!r�-`GJ�R@z��#3*n�gbP"Is�W)�A�	4~�@#s{E����%Jݟ��v����!֕��P9n��QA���ZV���F޾��X��S~ڽP"��#�8�9 �:����|ݕ��~���d�"j�T��=M��&�����:Fj�p+}�g9�����!
,rS0����ܔ���������:�6�P�򽗩t��wBr�gC>��'�$FD�d��[�XP=�GD��brl����z������[�?�	�|�kz����� oj-X�#��y�BЗ2x<�c�7A�����o���C3�{a+moƫg��9�%2��@8*Kap�WP�s��(v�a.q���b���ݹ� � x��p�Op�I�ץ��p��0�Ճ��	����k�
f���X��ⵧ�l��7)^���Ҽ:���Y4���t8gcg<���u��&<�Y7�{0^&PT�P�BL���@a�)f;k^��gD�.�Q�OɈU���31&N�(�����������4mr�&    IEND�B`�PK   T�(U��K� 	� /   images/cd1eebff-8d4c-4172-8358-6f93b12ef793.png V@���PNG

   IHDR  }  �   ���    IDATx��ߏ$�u&��s̬���_"��hDZn��� �o۲��4���/k���a�w~�_�I�a�G?�����&�ZY��"���RI\��a�L�Ȫʌ������U]]���=�3��}+3�Fܸy���q	l��l�����k�?,N;�|��8�l����R�:}쾺w���=Q��O�A+�{�p��ݍ������W�컗o���4�A���Ʊ66VE	3�3�1 ��L���|bwG�� ����E�Mk��`�c�T�fK�<k;���. ��p�<!�ݱ~3M��5�����6 $�� �Il-1��h4�a7��.��$��)�ԕ $����9A�:0� ���Ա�x�֭��#ߍ6X���`�VA�e\�v:���W��l����O��TCn��>�2r�������yf�/�i绺�G7n�:pف7�x��4�8����W��*� p㪝<���ת[��������1p]q�j��]����󋴽���X^G�S�G]�X�}wkw�
9�nW��n�k�/ �_�s��?����l��2� |0����h~{��v�Wf_��ӿtܸj��օ�D��Cuk���a�l�����f\���X�{�u��?�[;��/L;���_����z5`�Ez�ƴh���K�H'wk�����bq� �`w¹=��k���=%M-����|��&�k׭#b�iD `㎪v� x4�̈��e]s"	�睙���6hѨb֜Ț�4' m���d�*�Â�ĬaȊ(pqA�HJ*Mt�5���B�f��^�֑��X�Ξ�� �)�8�bĉ��OeѶ����,���[7o���y6���!}l��5��=�ғ�a�m�}���)��bw������-(�)]�-�i�`5O��#	�[�)�w R{��;"4<� �6Y�������wp/D ��˽�ד�t��v�Ȓ�R� f��(��Y\�JnJ�.@�EʒR�q��C �� �$Χ��� ���vN��Q2�7L�0ClG6�����	�g��{��>_Mp�s���1kZ����m�J��I���%�� P�HM�XP��5�&��BV�e���u�6k8f�ց_�T�u6��*�͕@]��
��4Kpk2@L�LFU��Ɠ����Z�"8 t�� ��YNۉ���'GSG�G�=O4����f��� ���i&sj<�mQ�q�g"��a�� i!\+tЃ��`�Ľ�`����j�W�ա�\ p6�yE(*1��2���0	@Y�j�q��gU<;H��nr �܌HX��p
�.��s���$vD�E���;XjZ���L��Kp�2A��T�X$����@�DN�Ⱦ �]u�ZR��f֌����o/��ݽ���p����|�!}l�cUm:������y�"���M�tA�BKVg �v��dm�Q�	 (Ufi�j$k��y���q�j�$!x�����.$�<�@��N��I�R�Y���C�:��Db����8J�kEu��"ޒ�*�N
��)~��-u0��F�+}. ��%q#� A
 -w�<">`UE�zb�j0��J �K�	�]�,��m� 0� ���8����$1֛�L#�*y)��Lr
�6��+ `/����� �������o3g*���K��4j���fdB,p1#6@�0Aۗ�3y&
�uq3�A������ȉ��!3w�35�fX�laf�1�HJ�89( D�D,�Np0*7�	�
^8�1S�1�_��Զ`6��#0܍�����O;�����[�Z(�`"8;� b��#r L��;�`�`q5��s7V�����sbe��`'r�	�N쀁�H]�D��0�3�3��RZ�؅@D�09��	�n��@p����F7��0� ܏���Cs��2��R7���_Q������_�o�����gkU�6xHlH��k�P������u\[�e�n ��#��l6��t��z��~�����eH���l|)H��/��t���\�[��Vs�q��W��v߸���׿Y���y��W�~�P����E1{e6��f^U��������鬻��� ���Oo������ʕo����On�� ���6�{�h�s�;�=':�;0 i�"�Q�u��ig�Uv�ˣ<ˉC�jO��խ�LRp���dZ��!�LZn�"�V)զd1RmYTr�,�� b䦤��X3s��������,,Ɉ �F�E�č��؜� 5�T�M��Ɉ؉p7B�.�Q`!� pa 7�Hԩ� R����ȸa�ƍ����Bd��I 8ca�#n��HU�*�km��NRiCw(��``("mXi˴���fi�Nn��d�7�12KHn�q<y[�@��n�R�9�<.�.�Z���ͣ�	1س�XXA�P��!����ȁTc�P@ b1��"Av�����Y�FB!!�`���6S7 �X21��3`�&8���� �r�@@V%*���ЇBDH�F �b�;�PJ��>��/ڗ��9/��{� ��X���D������%]~��%���BVEd9��&�����Y�DC@D`n���B������!�CX��>�Q����]��n�q@���~��27�aC��U\�����/�'��ݳ�싴XܦU_���6��>���C�����Rj�mƥb� �[e��>���{����lF7o~K�\�'r�������7?� ��Po �}���-��Ɏ5{����3�9�:z߫��l?���7��x�Σm ���6 pIw����kw�_�A�\�Ej_ݧ����+W~"7_�m�߄��7��ۣ���������ݶ�"\
5�٪�ȉ�N�|���G�Ż���&�CUo�t2��UK<χbR�w�I�B��#
 �/Q��(��S�J;��[ud ����/0Y�^Ea ��H͹jY�MI` �$�Y���)1��D�b�\A��8���ڲ����K��Y���q���q��Dn��T	lDfS׼��;3�AA� 2搌� �n@�n�pb���s�ى�����48,�A�M܉��9iMd�
n��V�1p�C�e^'"q��9P��R?/ܼb��j$��H8�~:P���{����rm� ة�O�;ء�B�@M���RO&�0d�I�	 ���ݝ�(lD���{S�9 �Q육؁�2�A��L`�
��s ��[���v���,�O�L0U���
���0@������(�
f'߫����0QO��i#��`�c� 1AXp8?@�����f�5"Z!�=��^i#�e�$h��| g�*��,�\U%x6dS1BX`pXV�	n��@� f�!<��렙A!�0xT��9�Ӻ��o�U���|�'����_�c�΁�&黶�\�t/��~�3����+s���6�?���72��?`�8ׯ��.��w��]��b ��4dO�J�/K�����ɓ�ҜbyJs��?��v�"K����2����fʾȦ�8�X��b䣼4���#�"�(Q�"S�r���X�`ɫ�7�,�w�u�h��� 8|���H���F�)%WH�!���� RU�P	{  TIn�¹�N# 	QɅrE*�kVQ3M̤s�A�j��HsD��IC4�6xb�3�A}T�`�fO"�N����F�n�U�p��斃��H&h0��;
��<G$���5;�23�č�7
�ɼ��kU��y��F������*3،YrΩ0��0��E@+&�Vۆ��ɂ	�ĴTZ��32wv�ѲW�]t'&עx��̉�b`w��C`�p&���d)	4�D�j�n8�9l�T&[e7���D��=��%'XN� ��hRf�^eY%Ǟ��{wGUU+�Q?�ے�/�wDhL ��u-��	 �p����#�yIrt*!q7XߦJx�"���T�( Y�����/$�
�1���?�c�"�9
YY�VK8�xpi�ɶT�B���)d�Q�-U�Ổ3��~�����BX���!猜�{Z�VT9���ѳ�~��po�^U��OwG��^�#�  �䅺y�_T��(��̑�r6�	B�Q!%�dk��f����u��W��s�YS��Y�3��[/6��Q��"}W���G#y�g?3ܼ�_��߿0r�w&�%�z�/���^����o{G��cכS�>�jJ�> LsG6I�yD�q"��J�} [  _tc�0w9�\']��9B�DHt�ف{�.k8O
�#�$�$�����] �ٲ���M�?� Ě�ݕ܌:�	�z�P�t�v1�aQL{F�ܤ��~���9S�W0�\U�8qq���. ��� n��+7ew'rnĮV;�ʈ�027�I�9� ��X��lv��~���f^���5��D���>H�>r/�WNNH�N`�5n֐#j�v���LD�w*�+rSm�Zkֱ�n��&���	d�bV-�h��Z/3���݋�X�HD�� D]���̹�W�݃����:w��9�����Lp��^�A�A���;�ɉظ /Vբi�kp�`���(ʒ�����'DH)���w�O��-KϚY�T{�a��B�{Ť`��7L�,+�:V@1��RiԠ�W��������3��$>"Z'�Ĳ�I\�X,���DTHM��b�0� �ݠ�@�7K�k DG߇nI�j�@D� �z̡��H!J�<'�d�)�Ua�����~�	q_�=�	N�����B���Z���C�ê9���K̣+fU@���'kǮG�1�x���`.���'���\�4f�۶(��yE��e�����N{I�<�������c���!Z�3\��3/`�U����b�:�(�Q���X�3���;��z&vx8�=�y�鄾w���<�l�A�O�#\�*����y ���$�b
 l1r�NA��F��Rm�L3yUQ��r�1��R��*5J�Q��:��SͰ�������H0{K\���8�{�F�L[IiˍX	yf��2���p##�A<� V��=O�hDN� �-�_��TGL��Da���;^�=3sΑ,o�c�=m�9���0� �+Sq'*N?%�s"	3�q6��W�:�[e�FnV�Y�Z݈X�qK���qf�� �������� g�VnV�i�����;@�O��DJLF��ff�e���4�p h����Ǡ�Tw6w�AV w_y�/e�����߯�R(�G���į�8jc��o�-��1FQ/jUOO�W�K:�
+��)P��#�  ���K��o�R�)�$a���$���8���ă԰�yL|��	���j�Q���ĝ~��k>�7VIV*��Cv:ξ�b�\=��,GJN_�J���Y�����R~��{�p?�z���'{�Ҥ=��} ��'="q'�8p��=���B9(���A�z;)=P�$����7O�8�p��u�]�����<����POƷ�i�|��v)��໢~7v#����?>W6�L�&}/~�7'�}�ߚ_��[�ίx��&u�'��nF#v4��0	��]�Φ���6f0�=��� 8��8$Np"U�"�)�m1s���%&f%|�@���u��P�fp�LN�`��Y��j}�J Nŗ�j��Ld)�F�1���C ����t0�N���U@�wJ�ٜ�H�wg7��������{/�2���SQ���c�Y�Y��ưB��Fn&�ΰ��Dȣ��+R?S���/�Xg��8��RQ�nK����v�� C�W�C�ɒ�D�_�ލ݀�����,e��� �z̄�z��������V
�Mv�o0	�lP3�X��٬�f>V���=���|�oR�9H�?^��ޠ�4v�p�$�H�2i�������K��c�ԣ���,�dk��_O�ζ���okHǺ�����{$0N'C[���ܩ�ޞ����>K���pd�]U������I?Y*���[8����pc8�5�F`éF�lc�X@I�!̺�EB���p�;c�� �8���[����o��)N�^�����jvv��o'��v8��g��1"�L���Cĩ۟o33�#S!x2*
���($�̂�I�/����
+��Ɉ( 'b#"��<�*͹���dfK���`��o�ۑBS���(RE��?���BÛ��3p.��y;��2�����j11X�L_�ļ<^�BsK	q���������K?U]�9�<�99�嚭?����Z��В��1I�8YS\����f2�Q1��Tw��k>S�2�/���p������P[�A#�\W��-o31�m_�>N�xP��I��0H��'f����VHn)Kލ�H�~ߓ״����u��	F<��~l��G��u���={�ZR��|vm@��i?�|���jWʓ�����Ǖ�ӈߙ��`���-�bZ?��wZ�����~;��BO�N)A	�!}�ZL����@4�*R�Xd�֣�k&�;K[/c{��!ϧʹ��ǿ����`m�m��a��ʕ+�W^�V���7*������~��`ވD mآ��lPYV��l��T[��ӑ��ia+�F�<$ ĸ$; V�8��t��V�&mf0�š��b��Ӿ'Ho#�S���IA. {o�Q��۝A'�*F��t">Rݖ�G�h���ݱS5`+oĞ�e �� ��0�2�9JTa��&ͶT�Ыi0�3 ��5��2�r/��i���i���v���
�^�0�ș��i
��Q�{�nu���W�_U��O�A�r�A������]�OW0_�n=Ni+�`�S2F�����x<�w������jI>9��k��s�YVR�<�yW=߷ߐb夯�i��)\�|Y���*J�����5J�Z���g]I�v�ώ�[�BBP�U��z�������Pwp3�����nF��ۉ�;�lr'�r��o����T6���T�^���t��֔��M�e����<G$�N��en��];C�4ݛ����+����+���g���:�)��8d�8�J	�2����8�s�����L, J�'�P��86�y?Xi�X��i�{�� �B��p�\��J�C��T�ݏ�5+��I_0 �37���6�,� (�w�lH�� �^a��|٧�  ʺt�&/�E�bf,zG����������~�tr���}߭:���!���'�=Y�>��`�Y-��C}*<���SQǎ���)���>?p����q-�u���>P�}�`�U��)��ʳ=��W�>j���B��o�����K�?�D����K^s~[�~ZS=��~@Ik�����71� ���e"��>�al���5Gj����9��(&{��F}��z�0Q4a�?G�b���b,:C��j���4�݄�37:fN�9�����t�
�9����߬_~�VuYh�}=x���E��!��!'CUai"*?|�#�����:KW|� (iQ,��x9^*C�������'/D0:!�����	� �!��2R��p_M����&gD�BV�$w)`}`�����܏���g�c��<~�t_�-���A�S��>q�w@� !�rF)iO�2  �s�{��4���<곤�Ẳ~���~G�vX�!��r2R@��>`���_�{N���QV�J"Z:嗈����X�����'�>��+���K�Ø���K�����$��9
�!��U\����W�e����8�(]k���9?�R���!�]��T�p�Rut���]�m^4�3��5�זkH咉= ���e�=Z�b���!N+�V��P꾟���r����~8�qQ���\y�`���
bU^|�6P�Te2�q����<n��ξ%�e��կ~o�{��]|��L<�x�̻����zwwk2鴍i˃��5����v0kǮ���y��C�Y�E(�Tn���1�ʭ�C�QCZ�..��X9oO�ZH�z.����|eK�B%����0Z��R�A�q����=v����Y�|r{�vi�<P@~���~?�C:�#��Z���)���{U];F�؏)pG�6x�o5�jJ �|�OӀ��o�߸f\!���������    IDAT�$��8�ϱ��ȼt���z����OS?W�'�z�����'�,��`�����a�~������B�\���lҴ��2K��Wa�H�٥�{<�E�.	��~���#z�=�����pߠ�Rڠ�?h;1���e�%Vp��� F@]�`N0� �1�@�����i��P�I�OM�Z������}n����ި~��3D���_���Nr;��h��^|���^�����k�qp��)c2ق�G���Ї�a�~q��Ѥ�:��䬧�� "䜗~|Gj-#�Vsku���;$��$�p�ĺ:���l5��0۲ݫy����$m'ɓ∤�cqL?-I��>,1���պ��|�uߵ���6�"�Q*N>�m���A�?|�S����m�R�c�5s���g��a��q닝��܁O���엎���|��%�{��u)O�<�8 ��9�C���}���x����֚�g?߶������� 60)�2� ����Pw�W�8��$0`��jBA�'u�C!����p0N���}p��� �!���o��k�(.���H�9����`q�+�Ҵm�'?EY�F"��{�=�p�nE�s��9c�"N
�`\J��}���&���������3��úIeݠ�I�yI�:���y���4Y�'�,>_]��u���دo���?����>z��mI�J�w�X�Dq{ƶ�?���K�i��*!Lq��tuK�?�P����0S��������n��o���ݟ�4��;� G�*���V_W_ކr1�0�DwS=��t��s����"��"h��߿{�֭�ǗO��3Y���ŗ�~���/�Qg��������TY��;Mڶ��8��3�w)Y�w?=���P	'�/M@�O��q��� �Xg"|�����>}R����<�5}��w���d?|�׷w�NN?~�Ԙ�(Ռ>�h��j�<<�'"!,-UU��k4M���QU1�Ǆ&61��
"		���7PI��N}��@(�KAd�H s!��~-�չ�� ������j���֎����*�q�ɖ������9���Έ���_Lo���F�����ة�EWј+{9R�1����·�;<��B�G� "ǖ@Zg�|�<c�ͭ��཯��D�2��F��A�^�}>��Ügu0y�y�{<;��Gy������q���8����X�2Ƈ���@eUA����������R��ޑoq��_�w<۝��
�s+I�ѡ��g���fF�]V���SXv$�% �J �$j��Q�FK׉�����Wz���3>�ן��HmB���l��E
���D��.��ю���9�7[\��\�ݴI���F�._���4[)3�_a���<����T�"�Ï[��V[��*���`K����zp�J�;�ez�#��u)�����I�����bR��O���?��u�����V����������ó�<:
�)k�:�O�>X|Č�nB@UU��
�
&,�8	;��KB}%"\�
�sԁʋ�;̙ �LMܝ��9�,-/s�dG�Nd�rMc��7��c���sAoI꯯���}��yI|sF���6��yֹucS��"�#�c�x�vƷ�`��	��,�'}׮	�_���[ �mH�F��ۃ�����ѭ�؇uC��R�;���;(��2������qz�+eyC%�r�9K�{R��*�|p2��4���a�ϯ��X!|�#ĒŬ�i!5��k���T�-H�8�D�2�1�q�T���"sr'"cH�E���%_1�G0�Y͂U���!��S]J<d'�`���,�D�S�/h�XFk��y�L���� kA!T�b*]�9������,�����`�{/�7���?X�U|�O5>R��+W��Wn�F����	o��z�s;��������l7�L�@���f�$|�
�O��9ͻ}:�eb���b��WV�~�C��*���M�q��I������I7�=m|܁�h�Q߯���x@�>�����r�֑�cfNT�B���	������������q����B�ma!̉E2�nj�Djf�UM-#e����]ۉjY�@�ܞL�D�����*檪�X���bfFo����^�t`u�l)���ݾ�Mj|>�g�,��U%x��@nI+&e��]���i-�+_����5k n�i�GD����_U����2���T[����?�n�w�޾��f��2X#�t�-|x�'a�%�F�jC�MF���� ��{q����sr����r�=��p���"~��?N��iWK���}�����G9�3��w��������n����W����Fy�>���c�d�`:ckk�QS�:ƅHh�� �j�9+���������fN9!���Y6�dj9gqgu3/Q�啟lC�Pa�����2sF���AU�,B�N}ri���,��,=]V"��Ւ?\��m����zOЬU�d�� u�!�6g��Q����^y�[���ؘy?�x���+W����V��ua2B�������t���������9	�W�_>��sFJ	A�N��t,��1��P��J2cC?8�01�oOg�|���'}ܳ�I�78����5|^X>
�>��ݫ}Gc�t�U"oG���4�$	�� �W735SS�;����)�T3g$r,�mx� c"���%rd��ȍ9���� �  �3S`��Zq��@U��s�4U誶3tI�@�'�a(�C�ə�劉}�V��� ��VҘe#�T�����dg���>4���D�ݽ[��gOqd�&_��_��\�_���1�zȵՠ��ٝ������c��R:��w0�����
�y/��.'8;�* \��J0����|�n��r.�idYY�#3��Z�+H�ݔ�PZλ}��yq5��<i'`}����~;���i�_���i���y�i�uJ��Nj�۾u.�O2�H�^R�ر��"��7l�jL&4�������%p���	��[#fN #��	� _U�7�5= ���vx+ �|DBu�p�1��Y����تCU[j_��4� �Ч���*
��qN9�9�)�kS<�/0o3�ڤ��� 3LE�vƎR�6f�ˎP��XCUP��Cr��A�x8j�w.=�'Jp%��o6�_6��N�C`o~������3��������"vQI�y�/՘����蕶;����V{0����)��� ���fĩC�������u�瞿�K�.a:�b6�������w�.�Z����~zr���,89��~^]x���6���bu��~�U���fAU���5B]�V71��SA�ٲiVPb�d$���C�]��D��s�w��]�n�����s�������� �v�����?���k�x�G�ɔȦ��9���5@� "����R6�='!"&�:�ZוrS��Lc'�!d��?9 �e�P��8�7�, ��5L�բ�	b�ȠI�"�L�*3`���܅�����)<i��_�����6�9F��ط���]��^�ŝ�Xg��1?����K��]Y�k�,=���Tu�[Q���f���~�~/�������������],�8Β4:֮U�)y4���rR���n��''�#�{i3- ,�QSa<��:��d���]���)�Y��V�_w)�����_(�w�!����Y��?���iFYj���Kӗ���3��a�ۉ~�7S�������}��H��=m�N��*[�:����/��9���McbrS07ĸ��dA���-;)H��'�]�$V�;�Go�-���(��()窊�0������bz݉G��ҿ:����'I��K_�&u�c;a1�)�4�2��^�D/���7ݻ��.u]/#tO��V�݃�y��䏙��(I�U=ťK���W�u���..=?��d
!�Çڡ]d�ԏ��A�;��s� ��i��6�pޜ�R9!@�4>]�=�ow��g>z�x֯o���#j�'O��a�op��� *)�����4�WU�	�"��H��J�� 㞃�5���?���)�Jh��q���X/|��<�ߞ�m��u���g:�N�ƍ�����ڵk����T���!u8�����O��>�į0���>�S�m�6����B�,�w&�ö����:�_hZ	�x�~_�	�}(L�M�$��PW�Uu%�źr�W]����ՐfѶ�	��≑�˗/ǪJ�h�O����\�ؾ���Wg�����/�j#��k�e Ūo��7�i�w	N@
�x�X&P�����jR��C�w�{��-��a� [��4����ն~�m>9	��g�7,�4�PUT̌�|��_�w�>�89�G�_y�+/s��59��s"����:'�@|/�����2�7�����\U�J����W! \U6��Ӆ� pJ[���<���oܸ�� �7�x�oݺE�/_�7�dŽ�_�v́��ۋ�sU�D���������_��k��M^��?�.χ�_c�_�L}������Ȗ���XJ2?,��@��F�����S�V�gAq�����8U�(ֱ�+a���+�w�t�]0���+���� �T�z�ˣ�횦��4����(��������ˇ��/T�
A"rJМ� �Ӄ4��qe�|�f�%|�N�!�1�z���Ӌ�nM����* �	)`1���|��v=�u ��x$��9�V��y�� ���OK�1(|��[[[����|9�e�σ��qj|܁Ow �:�W�{ځROkۿ���x�OWD"��H0OP�U�U�@�ݡ����3�����ڬ`����������ٍ~��^��R]�	���,�(�5��trX����4�F|�+_�����o����bs����{W._�������ƍ �/_0q]���_��=UM/���sq�"�����O�v5���:�QMG]ʵ�s���3sf"g@f
�$>��a �%�,$%P��!"�5ƓI[ג��S�uf�����J4����������-�%<�w�ʕ�4V��Ӧ��RK���-�����K9�q]���03��s03�FJ���3�z�7�)A���8ߠ˜a� � j"�"�d%<w�yT�B�D����A8!�C���T;ޣ���?���u���?����^�F�P���mۢm��ҏ*��Ӟ�?��i�_���9�����������=����5r���*�'%8+1w!63�|Й�:�/�eN򝪵?�������/��k4�ϫ�~������b�@�Q�9���Q��㺙T�d�ĉ��gf���Z4�{��s�����ޞ���/_��/��������������/��a�ʡ5�f�R7�@{ �CgPG����+�Bdf��vPSD$
��㣌�Ď�$]@VI ��q��*����HB ��kSp�Y��W^��t6��͛77��3�'B�&�I|^���V]�"��|v��pߩ뚘�Ѷ-��1��l6�0�L��\q��Wp^ҧp' �5�"����h�!����q�x$ :�3��[3��6<K���i���>�n5��d4���z����������=���=�'�t<����񒾓/t@I�B@�IH�,1	s���~� ���?0�n��>�����ʅш�����l63`��u-�k"��@3��0�ɸ�Z�!��
&NW"�$�:�h�9�d2�w�y��|�M�|�2-�L&��/����� �����o;���޾���Q]��� �Ax?V��l�97�5V�� b ��\-2-鼺sN�D� p��8�����V7�k���J�����[��ao{���×�Z,���9>cx��~��~����1}>��_U�WB75-�/�/��@�BN����7y�,9�;�fo�%��̬\j�D���dG��Ü�0#s ��SꯘO�r���#S�&��!d�[�=+��×�����y�gT�R�,�����#��m��}���jl�ꉦ�K���&�1W�8�ZTŐ�\~Y��Q)PM�u S]{����,"n����2&V#��6�r�%��.��]&�]��QTJ�Ή)PWC����nd$��"��su�6xR��c]���\93#Ɯ��,K�?[�EO�Yz�΅�w1I,Hߢ�岥�v;�:~�+�q�h����<Q~M���Y*ۋ^��B=��̞�}�=���X�w%
�v�����%�v�ųr�˞�����Ҿ����{��O>��%;��by {�����%���E�i�?��?��@K�����-O�QR���H��tx/�W+�+U¨+�ՙ��KE
���_�ݏ�[���t<�:쿴9���ɿ���_������+>��Ѝ|c�@k���S�2UfV�5X4$E!�h`S@C���A�3���,�=��g�{�=��?�g<x�@���x��!�o��?�) K �ө��_���W�������<)�� �w�ӥBLDER�O*t��#!�H�ǻ@̵{�#	o���pf�D�%,u�)\IJ
�����(���r6D��HrZݼ��&�ϤM?�X?��%����X����˕�~8�x���E廱�7ۮ'�.��B& �W���D��D����50-)�cN%S
��_@����ӆ�٬!�D2!%#�\�1Gg	}1ƥ������:�����UbA��[��[rGRۉ�}M��u���ܟ�F�ğu�g���'������/�ٺ�P?�{�>DdA#�iۯ/�^�1��<}�_�<��~��Χ)�2��倫�TQ���pYԃ*y�A(�>�r�D�؝t������D}X9;�"���r��Ϳiy/w��`௪��"U��R����
s��`f1�yT���ټ��ҹ��UA]��VA��Q5gÿ���2���{v��m>���Nj�ш۷o��۷�ʕ+:��h4���?o��"�,����R�w���'j&�L��BũvmG�h/���q��0lH_��l���)$�/�IA�W�F�4ճA]I=(�:_t��d�KH���\�t4��}��¢w0�Bw�B��l`!�E��2x�y���G~�H�耖���!-R��z�2R3���|�5�7�"ZҴ�vi��ug$b<w��J}s�Χ�Yv� �d�_��"Wy��4MKJ��)�|��_�Ó��Y��I�+/���� �.|��=ksu]RxD�s޷��M����[���ck?�+{����z$�f�SR������ӔJBU�eт�"&�m��Sl�R�M:��������������ߗ�÷������EU)�g�B�`�y�y�=tg�}=9�& ��]�����דɤ�'':�yY��ʪtq�EIm���w�N܉+$,qJ�̈́�KOȨbNI_|�RL��������*� �lg�}���}�/�B���:��0��"�(�T`H��,&qy���f�	y��b���8j�D��'�����{w?e0t�*��`c{D]�ܸ�&�yG�%��I��LL�I$�qX&{�Ƚ�ҩ����fvj�[�vAϓ�K\��F�k�?�\�������W������8_cvA�ʲ�����w"�9W�!Y0ѓ$|<����%~��do8�ι�?��4��I�O.�$e�K�Ue�4�YJqn1��Kݏ�ſ,����4����O�@x�w�w���n������M&p��������4�`�B��/��q��b[&�J��ŅXk3���tFJm��U�ˀ�����L=�o���}�YP�d���P%�����v�Νˇ��B���@uh�%+���>S��0�I�R�\����_�{WLs�Lb���`�i���wLg�|����XU��
W����u�̛�d�2o~�����
e1rZxmlp: �w��y�ނ�-��2��]`Q��-�2������l8��л�W�����$K��ئ��EMQID;�4$$$�6L�毛��/���;W�p6Ҵ2��h�r�i ݊�t��u�d��*T]���.���nA������� ����ߓ��=K>��]93��F�k�ʂ(�֩�#1)}�����fBe!�Z����D/�-�������ԏ���	d��B��묒��=    IDATj
�����%~o�"H�Tf� �@x���8������'��'w�G\~}/�mrܽh�E eل����!%v�fT�x���Y_��S�V
VV7�q3qp8�`�������]��Uw�#��	~� ,�<_t/[/.�Ó��M�|ON�l���}A���,}����x�{����eq߽�e��"��!."�d�����>�7�_:;�����:�IUuiY�~�e���(��Ƶ����n��E�я`��+{�'L���hu�b���9��]<��M�Mև�+���z=F��;�R]U�h4�)��e�Y��S�ŔT�,�ixt�\�Ϟ[13�>h�""`q^J<��[���x1�]�:D�h�>�-O��,}O�$�����D�.�jUI6�R
�����1�W���HUU�llq�֫<x𐽃�>RՈ]`y@�&R��ћ���� �ǉ������$8�:�����*�|����-}$�����,Q�9)�Fq>����ʹ���tP��u-�9��,'[U��%1��AV'���7:޹����v�������;X-�0����ae��}_���Ͻğ�����m�d+��j6�B5/g�]ȁݽw�=v�x��]H����0��RBP3K*�daݻ|��x��'`s睈8�d�X�3�>�����$!�"��\GY@�L�{��~�)��̍y����u��+����d82�#�M{�."|˯ǥ'9M)���ey�����%~��h.�b�u=�^3�)����R��y�m��]���ڞ����i~ûr�T���Ih���������	�N]�-��Ģ(���l��?���pؑ>��7�~��"�9�J�5x'V�SAI�"��;���v^���B���B����bT�G_I�\��/$e˛7w*_��\�uD^�m�>�M�'�$�47���I��`�9Y�x�;pa2?M9!��֧QE���"�*9�`��%���
�j�`8,&�M3crrL�-�tc])\AQ��m����nҋ�$����h/��-o�eqQ�/���c.�^��E�]��,iXvO^�%|Z_[>��sXN*������'eٲs�<����{s���y�e�ڦ_7����Г��Y������N�~�۩#�<���+��K�Խ����}R�vP��	�!bw$���l��]4x'�t큨�aR
W���b{o8l���w�?�����-�?��]�r%m\ۈι���w��^��~P��4�:�𾬮�q�bW�a*"&��oڎ�sڕ�
�����{"���
�AL�}E4�dB4c4�`XNU˪t&�"El�0��7ҹ�����r���ⅸw���
��c�0Srֻ���/�v[�&:���>tP(ԑĐZT<b��N9<إ���R�c��7�׹r�%f�#�r|�K��B>�CBw:q���m�8Q�yvY�.��N�[J�4�vY+vѤ��-_���C_��t_�-�c�"�:X�D�@41|մ)>��O��^Ǽ��8�bU%G�,��jw����oۯ����^ 1ѽ������y`S������λ�
����QxM�sVz��� G�Fy4��4M����)K�)�H��,��Kf��@;�L��%�h�b4}�w�ŋ��L�,��">�[�I�����J�)���)��=�D��S���L��y�����G�mlqu{���m,�f���N�ɹ���.�}�O"/�-���r$��g��2ֈ��w>P���w�|�c>+.J��~Z����/p�2��%ΐD��X���d�]A�Pj�k�4�s1��hP=����]�[Yv�FGP�JU%��`.��Kkc��������o	_ j� X
�6��G�?U�êPV�P͊b:oO=O�պC��9�>y{��yz���!D��d2�L����j�r�r��"X���P��h��1�S�p��]|��|�JD=Ε�#E!�4�f����'���������{|���?�'����ō7�y�:u]�
f����O%ςǹD/
t�Ȣ�8·��������$�����R�|U��ǹ���:^���%�E����Z�5N���T}0\4��G�(E��$wp�uM�s�jʔbi�v�4���_����H��B���h2(��{T��)�#�bJI��[Y��**�f�)W�z���AEL%��=+]�	X�	�������5���g����=qV��ʤ����d�u����a�ڳ��jf�tB��Z��C<%��, )�.��HsT$'�4GJs�'�����U�Xl�������k|��B;�0�6�F����N�9*��`�(=Ɠ4\O��=O��]Tw!����=.j�q�b��|��'E_��T�=g�����]�d�T����Lܤ�⯕�~�CZk��%on�������{��?��Ye�nؾ��_���o[�/�/�#W��;'���ʪ�(�<�R/7gɥ����ޣ3d��q*�T0�f����r���ݻ���e5,j�J�����f_b��~l��p���*�{BLfǄ��5�;�־�˱�F�"1u��M�
�D�3��y�{���}�\Y�� "�F#����z�*��Cf����J�mp�u�l�Zvc�6ھq~�͜��ҷ����/�z�h:���z�o/r__��t\�M^,����p.�iJ�rb�U-�|!)kG1�4�Y%���龰�?p���h���߯Zw�?����R]��
@<f�qP�n�L�!K����c&���z��㜊�Unv�N��a�I�k��0<7�[��TW�1&�����$���x<��_�֭[E�d2�������5=Yr9�X$u��라9� �, �9>�����GL&ڕ��,����ƍ<������,J~1��H�����:���"��eH�E�E�_&Z�����/Z۷x_�h|�=X��oï��^�(��C�ab9%HNπz�	�D��Ĕ,&u]w��/Z5_�pD�/
k6�7����i|ݸ>
+��mU���B����[)���,��e��v��4������=Yg��91��/�y��L���HU�n��;�\�o ���5]�E��5��1���ƾV�eI�u������ܾ}���888���K���%���:	�D�����J�ZrTՀ��rxx�����'��+���:����F#�s�S��d��e�ȹek߂�<k���n�/�'���i��ߕ��|���1O�fa�\��"��R�w�K,����ɢE_�����M'|>p铨j�-K�$�Ɖ�WW>�����VnnŮ���V��;gj&�E�s�[�
�h�o;�,*�8�w✊����RS*����ߗw�yǿ��;�Qx�?</��
ZO�f�%M�S�^L��Y���U!����^	�0H��#+M�� �Rp�"�W���8�5�l��}dJ�njC���ʛ���K�)7ߒ	Ww����������x�QY�U�æ#T�(Ig�2�Ѯ�3\���-���:��G||?�ze���IG7����u�+N�#�UX��CB�����(��$�|͋6YT�(��&8�)6��QB��9ae4 !�.��Ɣ�*�2��]G�W�$�	)���dXה*��Z�%|YR�
N)�m�41�LH� BhI��f��Afm0��7D�1��x�D�xQ]�]�=B��GB	(�(f���U5�@�em�fm͑bK�[�V`]��(E�h��pP���`�����ONh�Hj]H!2�$���%�0�Zʲ����|�&|m����nѻ{W|o�}=M;��ܻ�y�ߚ����Q�v���� G�bN����<��L�E�'��FD"��E^T��� uG��w�ύh��&��P�[�-d+jjs�V�9��l��ǜ�R����I�eH��hF�Pf��b�!֟B��GBBp�ߵ�v}PB����Ғ!��G�C��1E�A]��<��N��
�\�H\��b�1:�m�B𑤑 "������.�,�GI��Hj$I�CA۶e	>��Dт.��%j�R��@U1͙�N��k�x�b��༼a���J©�Ԑ�0u6�4���F�릙+�L�a��o����{��J��6�\�t?|�*J�K����_����˓�ͦ��n��5�BKW���T�y2T���H1��D�{�-Ɖlau���9�'�6��>tz�ʊI�Z�|��W�ջԑ�������Gw���:��_^Hʖ�$�r�y���V�%��$�rF۹��Ia���R캆v�B`8T�j��W^e}m1��>��#&�-P4E����B�����4���ܿw��W�P;�Kc0������&m�f�'yB{��X��-/�c��J�B�������Q�pP�:�4����l�t2�x:cg�hF	\]Ǥ4M��guu���5��֩
�w��}�����g�]���.$�]������L�)"1�$e�Or�*/ζwV���b��9�$W����v���u}����eX�z��8:�Ӷ0���!����9�`�>�~�!~�v�?@D�q����ҮO ngD]EP[��G���;l���rf�,�>#������qQ�_tϟ���CDR�$���b��0�$ 2q��dFgж-��E�c� ER��cR���dK��"��9M�[pYV�1&F�F�Gj(j$�#.�G �tr�^�!��������m���yҢ���_�����'�X(Y�H��9�-�B�RD5"^Q�UE�HRC\n�$	R��8<"�� �)R���S
W���fGQ�"���=J)1�:,����:O��̗5���Ec��gfQ̢z�$1o�pH�vʣ*s�L�=t?����}a'���!��M�lX�8�9y�R��=[s�%<�<�,�$b����s"�D�j�hf)��߿.�o��{��?������GL��������eaQF���=v�>U�r)3�'�$�+�	0��d2���{�ܿ��X_�Yٹ�p���gv�p|<e2��"u]0K1[eW�z�	�D� "�63�����2�W���*+�5�_����[L�S���l9Gz���T,��\UYor��67�X�\�\gme��.k 1��89:���]>��3�|�9�Ʉ�:,��Jԕ���1�p��k���k�z�ò�,�{ۗ�h��+�)���@�6��������������w�����w��	�,���O�(��V�^L��Kp����-����[ߺ�͗6Y]U,uЖ�d:�<��Ǭ���o����xX�K'�����9���h�"ބz�M����H�^�Ef�D���8=	����蟉�2AL=�9�0�����:�D�[E���\Љ��D/ƗɞWn	���l���?��	ƫ�|��
������&���J�D��t��p�Zb�������r*�̄����5������e�C�D4!�e�-9�f�)[��`���Y-%0��zo�|!����f*�rZ&�����4�u��Ήa* ��G��>�g/�W���p���DOz�]�L1��s��O���m�SB8ˉ��@"�U]`�ֻe߳����8�""�Du&��P��+dg>E�೎/���ƻ��������_�8�MD$���3U��~���X�N�I$��&̒8����Ԉ9�yդ�h2�����:�o�?z��O�n��Ē�9AΖ�_�b՜�(5�I�G���ߣ�;��"tDli��(|�O&G|��8_҄�nMp~���5��<b��>'�S&��m�fWMO��'}Q<N��f)[v��޿�gkk\���K;#�;W_��˯p��}��'��UD����b�]��k�����׾�[o���[��X��RQy�I�*
�ʓB�l�p���hQrr<a:��R���Q��Q�%W��������;�e{c�A�
ɒm���J�D��хDg�:������m�{�3>�U��;w�����s�e��E�w�U*��>U��A��p�[7_�;����z�����)6İJU�����.
?�iM���g<Nܺ�&��X[����s>��
'�m�	�*N ��}A�	�ق�-89�֩����I�)���]�w6񞒼Ǻ̗�\�*zRG�\m�@�X�/�u�ؿgbɤNL!H��M:{�Eu�t}�29���"!�P'x)p^Q�ݜ�v����]����M|?��߱�6_�إ����1g�i�3�xvOK�{9�5d]G" >���؞�W�!����Tɦ�6Sn�9��Ϸ�'��9���{�$/`�?�GWdKe"��ĮG#�@��|%�-��BL	'�� a��.y�5�O�ED��&��,!Qi���Hw�n��YbE��1�����:�Ǣ�vU�C�}pN������2@_����Bԩ�:ˉ���W�G���.�|�0�K�EM��>g3�#Q����$�ߥŔ�����8=���σ!�pb4�)w�|B�ɢ(����aUS�6ؾ�
/�v�|�§qxrHA�a[�i4��EOnP�	��|:a����L�W�յ-��t���)�=d�Ͳ�/٩��qH)���S��<U�,K���x�����w�ŭ��3('���$u���']���������](IB�y��5������׹v�5���Qj�e�DBgFH�������kEQ��oP���ؠ��/����R�k�Ǔ-��5����^ӂ�H�=�p��K��\���t�	�k�h�������6��P-UA:
/x�Yۺ�`4�HI���=�yC"���;�uH!���N?�O�-2�ҩ<�{.+٪y���Gc���v��[-��M�������!�d�����uvCg��ٓ,��P�:��@�ԏ1[�]�O�ʧ&QA{k�j&��소)[������W�=�_\vz�2Ձw�ښR"Z������T��-�Kz�Z"�EW��j-���RB,��e)e�j2�E�1eˍ�C]�J&X�Zx::��� �9!u${H2�Σa�A+h�Ę�EYP��y�h�/�+=E�yAd)�6�4�K�b��H�w2>��-0���߈�L͂!��ⱘ��W�Y-���o���i��&bD$?7jΝe]83�\���4]�Vg�R����{s��z/�S�n�0uw�|c\��x1e�4&�E fk��<��w�pI��+l!8�~�]ly���3I��C������b2f�������JO��-v6j�шՍk�|�!v��m�MNH*$K��\����(��YJ��b��落�����2�`<������5��'Nf�E�.,��E�Lr{g��pu�j��jM#Ncv�i��󖮝�4{w9>>f��h�&뵊Q��($E9b0�`P���D-�fmG;��t%X�F�o�h��y��0ZYa0,����2�]��|���!���]�/9\|��Mx0���b�e�/kB�bN�ݵ����>L�S��GH���56�����Wj�VG���
�+�ll�ě������O~�t:�=>A,�4�-N-����
��ɹ���'�D>�@��h�x�כ�Xv���]Om5���GJ�.�g��D9d8K�9uX�P�M�Z.����s�E�Qu�k˚y����8�p�'���2��|�!e͞�~��k?S�:����ړ��I2���B,I�X���%�1�]��%��^��\~&GÚ��eRo �Q�\ͧ���-s��U=��=U�y���L�9��	M�е-��u�)����*����>k�����*!VV�X[[��+��$��	M;gz��.[lEN�/�Ӭ}Y�����a�H�%K!�4 �˔$�nv�8�pxX��;u�b�*`�K�_�a�["~}�?5�EQJYV� a�N�N4�>��?|x�)N�K���H��۷=쓒&g��Ÿ���a<�l�[rS�Z��K�I�)�)i3��D�J��a�if�ܻ�	X Ԟ�^��+׮1v��q	��f�C����H@�1��h��I!`��"�9��c������\�2��W�X��a�����C��%�S�ڴ7H��d�G�ޣ��̚�q]��1`\WĶ�d:c���}~�{w�ppp������ߧm��Ρ�A���pEEQV��6U�5S��vyp�{�G4�zw�pr�G�Z�j0b��^�z���V�ͭ���C�2�n&�y�|��FL�l_��hD{7�"�	`JB� ���p��>�����    IDAT�����|�*eI=2����ڕm�]������!��*W���`��������1��N^Յ�,��Y6'8�42TD���)U�yr������%F��E�ʙ'HUz헜Z�R���αUQa���"��k�򂤯� �KS��Q�1s��(}EU8W�
Ż�d�')v�d���ު���j�Eژ�UU�����0��c ����5�vJhbꭔ�E�`KOZ�wc��Ĥ9��N��/D���^�[��VB����sTUE]E��8<4��	)�)�(r_Ԓ.u�%k�o�2���w����l����|�	��1 �0R�'�]��<�������+�5��ܽ��'�E�h8fc�7n������늢�E&�C����}��qpp�H"���/�%W�!j�,�!�R�
# �Q�>~&^�Ǉ� IUI4�L>�"`@]�Rץ��Z#!&	M(�s�{��B1��i[�Yx.�W׵��t�%"9�o������:��{g��lh_�J�'61��B�@�k"Ė���Ķ�XK,
��`m��z����:x���]<���fKR#Y�cy�.��L:,�ل��#hژ����5�zؓ�D�F��vq��u�#n^��:NNN���A�uL�'ܸ����q�����������_���l�rT�s�e���W�!�+�,�e�#�4͌�Ç|����/~�ǟ��d��FO2!t]H���V7���-fM�q�Ǭ�\y���s��O��ϘL���~���ˡ'B�~�(&S�	E&$�&����?�o�����ܶs���yO{��+�U�W�\�Wn����o����:�(hlll0��S5���XZL��w��&�����}x�4��ʗ��_�,t�
KZP�>PDZI�������G�ѣi�k�"!5���Ɩ�����ら�~�>��f���ˬ�����J=P�5E]�R�ifL&�̧��9�����v6��|]�Țؔ���pȵk7x������u�
];ez|���}��a��=��t˜�}!	E֪�Հ��-����rt����=fwwYT�[�Bz�bo&	⠨+VWW������:+�1�~����9��4�H����Sams���|���x��ׯ1��������)���D��'|��'�u�g�9xpb�R���Ң�%h�˯���o��������&�̻@UUl�o�g�����op���S���ݽǝ�?�����l����%s9���pj� Щ���If��c��I���������P\��E�W"-{���A~9�i`�eY�`P�JS�� A�%)���mu���7���e��o������ruSuE,�I2Ra�Y�{1�	�����V��}.D� �]?�)�T��Cb_%aq�G��	]B�H$�w$1b�'���=>��R�z�7^c}|���d��u^y�u������4�)�ù�^����;ʅ�.JW`��	��s%��p��ع������.,�G���<t���eA��u]����;�;����w�bu�fex��h:���G1�Lr����X�R4[L4".��������T>���~�7��_��g��bT4���E�1A�2k#�.��p���m��/��@�������6e�畓�%C�z��/�<a���E BE�T���b8K�4�l�U�"t�޷��<� �I@H���!U5�ƭ[4m��kTU}Z?x:� �SV�m�z�TՀ��b42��ٺ��;9��,�I1�5-��CN���6R����1u=d8Z���fY]]�I�C�����u���(KO]ק�O�L�\��V�ϧt�c�������9:�2�wT��s�S/��W7����3^Y����6k�EAQUT��tQb����{����������î��ҧ{	8�qEE�����o�������IUK��h���}����w�����#U`���D|r���Y�R�cF+�������}���u>��~�ӿ㓓�e���^K�������tμm�Z�d��	�x������笭���l�K&�����pER-!� _���ş���?���q��k+���ks��<m2�YIkc��dkm�O~3��_���kW��!�9�lmo�}�*߽�=��G��@�[7o��+o�֛�amm����ϧ$K�c���Nloƽ{�N����B��������kO4V��;��73�RR����peݚ;��O�#N��$���"2J$ĬO1d��sc�Rt�-��>P�(�Sw$VV%1F��EYX5���j!]�X��R�?wItu�&���[�_'���omŭ�s1r,$�&/�b�­)�q�.+�-m�xߧ49WbLU)ʬ�S���LC�!D�)�n���]�ݽ�����J�)c�\��ε�q���w������k��EB��}^��m98�P��A�+��U9���������a��:����	����f�>�ri� X�t��]/\��f'�A��d�1ϑ�d+'��&�Z2��f8'�pr2���8Ga�� ��8�ݯf����b�{�hh(���Y��3(+�Fe�ꜘ:��J������c2mh�H4��թ�T]q�7��M@�*����֭[\�v���uU}J@;�m|�O��g�?|�g���?c�y��!Z��$aD�V��4������6���:o��W�]cu<ƕIF��S�8��8�EQK̛Yւ����|���_�ɤ��<�/36Gk���k���M�������M����w�:e��x}���Y������ۇ�g�~�����LF�x���Y]]gck���+�olc�cPy��ʠbmu���;|���3�?�Pl�p�hA=�}�*W�^ge}L�"&�ٝ;4M�l�҂�(]�D��`D#�a.��������7YPU>����8�/*:�62�޹���w����׮]a4�4G)�FN=Ml��A<�H�x_CK��-��1{{{Lf-]�9Q��(����D5!�`gg��������_ccm��x��`p��s��Bb6k������=<x�l6���RP��=B���9<�=�>I�)Q3Įn�)�������D����%�8,X���{���B�^��x�$X����������Xx.����8��z3�s�d�l�=z�B�Xʶ�b�E�OK��s[�؄>|��L�'���w5����m6��E�0���]�T5�w�re{�c��Wo��ko�M��p���r`h�R�H�esz��R�tm�d2co����u����YY�dee��f�<�i�����?K�v�09f�	]�S�(r�F\��,��J��>��"@f�,fk\�!��9E��IR������0U���9�MV���˝	����>)j�OA���m$�
�E'BUЀ����� ���,P�!A9j���n��bEYgW�z\�H��h��ԣ1/]���[����os����1������)*_P�R��5�?����
��_����M�����,K�	]H�6ulllp�O�!���?���k�WWr MO2���hq'�z�Eb&{Zd�_j�>8��;�?�Q�
Qq����������z��ׯ�V��AY�Y��5�����@�P�UΏ�uY�N�'��1kZR��S�E���\I��J|5ė�a-lloQ���J�H��u�����mmg��pŀ���y��^��͟���>����R"'=�jf�[;W��wn��[o������~N�3�mnRWbA�r�:߾������W+����4��n��`�(|��y0�:���à�p���������w$s�j�p��xe_V����ޛ,Ir�{~�����1�\��YP @�H^ކ�Lm��`2�B�2Ӫ��3�7��� Z���nKj�� 1՜U��c����8�Y ,Ҭ/�VȪ�ʨH�����N@������p5�V�f:�q9>g>�3[L������S���9:<d>��&	�+N(�p�����^|���/�&(��@Q�����F�sA��������fK�UD��?�m�d�t%:{���xM�<M��tF��s���?O"�v>x�%D|�����*>L��cR�VN��hV1cK�)�=�,��V+�F%,���"6��!K���S�>{-M�;l�;����orvz���*;�#|3~v,��%(DB������t�x��zA�������3jy�?^m��Bo�$��Z΢%�j��뢁��W�|�3K��	��4��� TD���_�Q:�(
�}E���01�!"E�1�g9��+���sͺ��cV����ݨ�B��`��G�C�h�Ӡ�@3&N�,�hM%e]T�QXg��C������;��g��{����W�$x�AI�.��J�f]R�t�nT��NN��0��	(6Z�8�ع�������Oʭ[�h��qL��ZTW�e�"��*�����y�m���ҜCh�r666����w�{�t;�L'E9ie�d�@����0��&K���cgw������\�ˁjQp|z���S���n>���bI��	���k�7TQb�H]+F�9/�/xyrI�u�i������f|9����$1	N��l�D�w��sc��wﰾ��N.��x��K�|���d�B������~�.?�����Z#�R��1GϞr���ň�d�
�BJ�N��dlo�����v6�v��Zo"����fT�RV�����m����~v��z�Y��G����.·L���sF��XE��u��h⬢��O��6]>x-!hq.!H&>t�"7e9��*F?��]�e��e�Y+"b�^y��Kſ���8�Hh솔x	`*�&I^�ܿ��q|�굚�>@AD�	Nh8z�b�����"?��	��&x�m2��5n�챾��.�39=?c>�7#�f�1�V�4����G]MPi�+�<���`���M��6F��m�`��.k�,�b��"7M$��Jc���j泂�tJU
�Q^����������������;�5b�	H�����"c_Or�з�(^V�[E����AB�QT��]���a��G<7(�����a�U;*�s \5�A��A_wQ[5{+�«|��	�ST�F���o+TH1>ڸ�(�A!J�Zy�]���/�.D/�X_�tk�y�������O�m��tp�1��#+���<��ՖD<y�IT���]2��B�E���Ԉ(�����M�~�m~��coo�$m�<,���((˘kt�2:v.`m�s��� �=E9���)O�1�W�J�N����m~����p���<�[Ǽ�y����/�/Jfe�d:��6������:[k=�ַ��V֎���E��
���C|������s��m޸u��A�4Mpa�kT�:��ʯ���WY�$�*���������F> Q���7�����gO(�K��x�#-��������oqcg�V�x...��g_���Cfe�$)e��������wٺ�K�Ip����#>��#?���b�eP��E�v�s{A7ﰵ> ��d-���-�V�Ӌ�_L�$E'm���JR�����ذ-�~������x����,��]��ua��F�%\����~���+|P��H�}Ȕ�\�M�����^zý����s�1~s�ר�\PF<�;'�YQ>i��פ<
(�F7�R���9�	���^_��TP�뵚�?$��/!(V)�MW�'�RE��d���$��u����޽�9ؿ�5�lcΚ,ϥ���J�"�6�F�z�I4�\^����s�n��9�y��.�7vٽ��d6���"*� �K��=7��F�9�x�f��|��)K��G�}fV��W�=V��`S|��-1.N9נs��)�N^N��h��􂁠�C�i�+4����o!�����S�h�5`b�%����EX]^"�P��B�Oy�Z2
\G����H�!&�xoѾ��̅U��M�A��R�G�ΗjL"�VT����=���n߹�;����?a{g�f�(8?�����dBQU�pɀDJ-%��Zl���S:���5(ɘL+T��%�"ow�qc���Gܻw�[wn�j�(���s�<y³g�h�q�S���c�FJ���0"ת�*g\^�svvJQ�h��TB��r��]�}�]���0F���>~ʃGOx��)�Y��(~Q�!�s>�����ҷ�e}='5�4'��D��z���r6gV��rR��]ƣ)�6t;��[x7����ٯp������QB*��$����鈧O�s��.���5�7n�`gs��ጲ��������g��-�N��Y�1Ϗ^���3Ƴ)"-L�Q����6���(C�e�ł�|�pt�x<��/�֓jSq��͠$E�%	"qj��t�����$AJ�$ }v\U�责���9Ϟ<�7��/��8?��\�DE�e���_	/�(�ҳO�`��Q�r�$@)&���BK���y�4|���������g�uxSB���T���[׫�;����%oP%���]Mx��y��������՟��o�X�U&��"�mފ���ky�};�@�]
I${�6��=�֝7IjO+����9NN���8�]fs�k\�
� �����.�y������t�~+es{���999�r4k"IT�͸48$�h�؆=���WYYL&��666�ی�l5Z��(B@y�8�wq̫��#K%t�E$o9b��d(�QhІ�5�ML%E�+t�1LC�F�(�p��Z�H���c��X>D���x���T���W��Wk�<{oc�l��iE�j44���Mu#U1��	E����}��N��`ݜ�Ι/�+��N��������7�bgg�0Ox��9�>���!�јEY`��J6i���@;��{ܻ{���8������9��r�r�hz���͍=~�����~���&y�CUU���~�'���/�#?N����^�ٲn-A�E�ź"�D(Eb4i�����ݻw�qc�ԤX[2�y��1���o9?��|8�v�J[�$A����rD��T6���(���;��+vw�9::��!�@e�x�,j�(n�9�n���D|��Y�_���vH��S��-J�>;"o���;wnq�(v�6������sܼ���0�����}�.7n�@)�t:����|��!�ć�R�� �£Y�Y�{T�o����u�EE(�.M��J���.��798�.����k��D�Ơ���^���΋�>��3~�O����e�yZk�jb݂��]D�}�R�%�k���Z�|[�_w�^{���/���������^6�E�w]e�%H��36ت���X�&K�5��^�h��"���weY�,�V糿�_a�V���tU�:���!z25{�׭���"r��-���`+��Ds~~Ni����Ռ3�`�k�3��(899���)7�{��B��g}s�v;�����j���EH�kޛ֚n�e0�n�ɲ
V�󧨝�|�����B�DH3���z帮>Ռ�B]⛍xxu-��T�Z�(�5X,�ɳ�,K�=�wx�_�����4�n���:_�[>���+�}�k4�$IP!E� ���eFŪ��"tZѤygg���I�YLLg��`��veZnܸ��FDe�G#NNN��ˇ|�駼<:�(
M㥄D�[T��7�����I�#������ޣ�������u�oq�����s���!_|����o9>>FI�l6��Dl���k�)� ����(M��F���^o����v�I���(T���;��Jst�"���9\dI��������&Y#ִJH�k�.F�h���T��J�e�0�/��x��$�#׎�/� �C�L����#=z�����ۨ��	,��^�h��H I2n޼������Q�G�<?<�ɓ'�F#�fZ�(W!:'5i<�"d�6���vsnݺ�Z��%T;��THL�H����kl�]P��H��,Kʲ�A�a�>�G������?棏>�W��Z�h�$*6˸FTuu�,�����]nb���J]�}��u��\KgfM�j������?���~���l�,���[�[7��eL�s�y��^[k��R1Z��t����c�EI\�B��q��R������_|o����z���������tT��G��d    IDAT@�I|���U}�y<�D(M��d�+$�A�����{�TSy�A���Kϋa�f�v�O��ؿ݂`p��#&�)B Q.�?��P�p��ʕx*��0ڒ�0yn8��2�z�<퓦��1;���'�Fl��Ȥ�� m@��.���8&P1] Ҧ.=n1`~vJ���*����7�7�}��W�4�8yV�! ��X�9�c��5�h敥P�"i3��VL�/E�	5$���zM A����$x3��'̫�m��.yk�v��1��$9b��9���.�g]t�&iwy��>?xs�SB&T��8�dt�sbk��Z}���]�-y�|�� ���)Y_vY�gԕèA2D���y}�!z��,���1��8���}�;�w�ug@^ըI�0�����?>���(�i�&�A޿C�o3�Πq�����f ��{9�BSzK��RL`kA��|���޾s��~�j���x�%-��Zz���_�	�������cfG��я��Q��U�����W�@�v !���s�Jpd��&twY�%-�T����������wz�䴶Zm�4�5&�X[[�;H�zG�JQ�9N��.u�#oH�-.��O���EB�:�qA�w0e����N�Q!�,>�H�ٿR;��P8�(��C�R-9E�K�82���n�c��/����_�O��O�͵�}�m�j��=Ϟ>�w�����o�霾�(U�I�p
�n�kn�z�����,ׄv�{Xզv��VD�Eb���yYF��Ω�0�O)JC�Y=��s��>�!e��nVq���|��#g���}����3pe�$!*�E"��-��K���ٔ)UƽbPT.�i�`�ޢʂ��V�٤���R���myO��>�M6�zk4�%�0J����x����$�������� !�R_-P�N���D7ݸ`�f2�V��I�N�T��i����4�*����� U��{��T�uJ�%(�q�k߿��������^W���$+h����9��e��O���t�pt�h|�V�&1	��W3���G�e�t6n��$�¶���D��2�]`�������s���m�ӡ���v�S��q�k
~����*&�	��^n�TV����Q��^�}W���6O!�t��F�h��"o�ź&p]��,gms��7�*��P������Y	*�;�`��>o������Z	�.�8;�уǜ��,\�����ӝ���r��E���������{�E�t2a:�b��V����N��Fb2��n�fkg���-�<��/>��,�9���DY��Zk>��i���W�]�VƬ��,� hu2���mm���esm�^/��G��GF�	T�bQ-�\����ǰ����������y����B'h�%x��ټij��ڤ�A$���N�,	�vމ\HJL3FLp��IIL���Q%"c��Xg��1q&X��K�窕�,ƀ�
������چR�w��MC|��m�}�Ngc���8�ء�f�6�޽���g'����޽��۷����9���<�����,3D��K���@�V*���	�3�qd49�$��qA���yJ��Z�V�6B��|��%'''��q)�h�]���0�8::����1���V*+����{��4Z�$�։�i���A1��c��p�>��? >\������'y]�����n���@��R]�	ޛW����4��5;�oqz�#z�d��6P"�9+���?��?������������z�����3���6!��	���Ңoy �dCp� �<�W�'�����숃�,���2�Q�)����%��S-ב��E�ƍW)�
,�.	v�h4�����l�n7#�r��y��HL����(_�����������׻��j"ˢ9��5}���w��B|��k�RB�bk"�|=.*,sa�HX5�}�E��e(T��������`0��>�$�h�|^0��=�[�tY�3N�^������׿��0�s-�$y��t��W�p����4N��K�B`<q||L9_0�ssw��`��"{�>y���pȳg_������?���xF�b�%(�,���'�s�v�fk�O���LB��1��'hI1�Kj$�Ҿd^�Iۊ�{�p$1^,$i	�|���QQv�iuԊ?i��:��<ĦPC��$���h�)Y��q�uAK�vY`�����Zu�u��^�H�;��c��Z.�%''_<cVN����j�Ij���I�ZX7���ԾB%�nhiH&1�f�p.�DΝw5"	���
.��8|򄃭���5�z=v�n���?"Ks�o޻���-��.�ل�O����CF�<Y�!1�9*a%f��`�!���5\ښ��S,&T�ʥX��ϑ���xo�
噌/9:~��'O8|�yQ�t�h)-��4���j�q�"�R�R�D�\������%�����u�*��	^��D�J�ȮJÖ��y�ˤ����{z���/~��W����?���h<>Ͳl]'��^!��#ڈ��Z�e�Ue)W}KaLs���t���M�r��~��1A+%Ai��!�F��y"a������TR��u͙������IxM�
�L��S���b@y�R��huKUL�O9?;b:�E�B+�HҢ��dk{���\�_4Q4�@�W�I�o0~�1pVJ!A��QU%�٘�x��fT>.5��.�:�+b��9�@Y����7�����Ѷ�Ղ��A}Q�xƇ_��ӫfԣ�Ҝ:D�x��(E����(e�Q:�3X�~���]�I	�Py!1-*;DDa�6MB�縺b:�ɯ������3f��		����_v��I�1QMmd*D�V�E��A)E�=�E���;;[�Y4^���(�Ŕ'�>��ɣ�py�t/��/:`�x(}�����,�2	)�)tPh��i�D�_'�x^N��iQ2��)�%$����c�b�Qe�!(�.T��:�o�77����`Xb@�53�f�Dى�%&r�$P�|(�PTT�)ò��:z����U�s��ZB������ٳ'�������!H�&�A)A)�ҁ@���2~t�6��B䲪&�'���ޡ�4"�D�S#xWq9<�<}��v�[Z�6��?��w��更RE����b��/x��g�'8_�[,:�x/,=���F録X0:�����O�YR��-XrjU������+�j����t���H�I�ީ�z��cV�E]a�IB]�WԐk�kR�^����υ Uei�rc�$A$/-A��}���L�<TU!�^O��n����A���T��dY'�z��ӿ�ȏ�u��%�:S�eVV���9|Ղ���WH�7Mv�
lcB�""��
<����+k��V\��9��#>D�Y\c�-#iUK�7�݈`�EU$�;�lz���s��ȩm�h�!o����e}�����$����z����2���_�o=x�r�p8d:��� cZY�~-�"B�jJ^ݑ}��s�f��`���L��n��x3/�?p̖���j�7:�t���л�T� �HZ5i\�y�j��q$�$	:i��Qdy�v�M���jaV�(�Ap$IF���:PU5*8�/Ny��3~������)�t�Q	�����I�&��x���hcل(Qe"�Iw)��bX�ɑ��W�`H�൥���Gǃ�e<<"O*
���:��FH�xm�����<Ƥey�Ea)m�V��m��*�(�0Z#�B�cr9���/N^2�Ϩ�8*&Մ��2:4�Fŉ!����
���� <4~E�6�RsM�(��@��D�T@+��btq���Ng#��Z���sM+���|�t:���X׎����.�gq�e""�Q�DB�Fi�I&�
:U�<���m�����I@�L�J�&<�q�W�gCN���O;dY4��Z9k[�l-��������/���Ǐ2��"(�ƈ�#^����
���E��<!K�Mk����G����C&�&ic���lؠe	Ҩ��5����(�bm I�>>Ьe��kJ^��*'4������Z��U�A�އ�u��e�
��
��V�8��7?�:yxy�8__�닋Too�rx����;Q�����!�j�8rJ����[�B?�1ʹ�Tu�TUi����s��2h��
��jσ��}���B*Jk��VB�j�oz����^��Õ[� ދ���-[�W�9ML�pED�DS,.99~�'�0��x7�t����8�h��u��J��l���q�4&����i���l��Y�,[tL M���}�,g6/vD�b�ثuݪ�V�D��׵t�ո:6�ZA�#��}�`�J�-V#��AGT��f�7F�e9�Ic"��h>�tT�zE�^%�i�Uѧn��c�(�1:?�����GϢ��GR!z6�i�1�n���5Ƭ·J���ʢ����GO����$o�u7��v�R�Ep5�ٔ��3F���bM�C�9�I��k�$(�N���삗����<!�:EEQV�N(B75>AH��_I��H�x����_~���h�i8<�S|0(�V�N�G��f:)�6�/�ll��1㎈���(Y��b���hţ���|��ƀ��aK��hƳ�S>z�%�ш�l�B˽�C�A\U�r�{�L&��c:u�%��(<u��h�:�IS�iP~H[1%o{��x[�G�(ݼ���K�; ʡ�`�soy���wYT���$�:�
X�N��t���S��O�m��$��x����@�%�ɬ�U[�<#1m���*t+mI�
	<8���_c&�u�B�����l�٘]�VYnڜ�]կ.�W��oF����~��)x��DEDi�m0�����|��ϊb2�v����)��]z
���� ����4�x<֭��ot�_b+%::ŖE��L��^�#�-���"�z�[���h���XV�l�F�Ң�(Z���������^��+ct��]�Ba��-�4I�}�%M<��-0J�U��&��{F8Y��JS��M�6�������./��!�$��ɑƻ,6A��Ҟ�.���C��Nא�ڬ�Ek��0�̿
��~�k�f_�����ﵓ�G�xdV{s���+�/���j�_q��o�b�4#����)�ݖjN�5&��Яb-�ق�dĢ���5��k������������UE1��'��Z��ʤ�������fιՃX)MՂ�d���3�=����q9��]ۤ�
k���HM 5B�
�!k����`�ńZ"oL�mZ������
cbsrt���G̋���'B��D�^C#
%��L8*.�#�ʣ��Y���xhe	��wnߣ\�9>z���|5&�bJP0���L���a\�XB��傋�S��Oh�����o�L�V{�2�sqq��:��@ek���.P���
-�o�˫H���1'8�b�b�=`k{���]���i��Q����7�X,JNG�J�5�]�������z�x�s�P3��<;z���ǤiJ���h�jŕ����%�|F���q{�F8��F�6F�b��b����t�$�ps���t}.//լ&���;�6�t<f2�dQ�i���-���=K�]fl+uM��$�HC�_�ZYZ.5�_���⻖������	��|���S�|��I��Å�^�?6J��'������f#�pz�~���?��������1���E9wO�q�*+ŢJ�"��f�?���V����^9Y_�u7�Ʒ�9PJ��*4���('���̿���^/��T$	�DB��κ?jIY����Z�W$H��ؼ)#TuE1��=�����z��\#��m�����B�eE$�/я@l�L"�V#���Y�I�����A��g|6�[�v_�.���\��;-2�F�\�7�^V�+���b���D�E�Z,V��Չ�ʸ+�4&�:o�����(�'g'<{���'���1I���6n����{�9I kKL�$&gmm���5���UAY.�E� 6�������r�~}��\�x4���!���>���#�<IQy��;�c�bVVܹu�!K2Zy���Lo����EM�
�3L�ct�w��t�W�,�X__����z���K\ KeI��rV���x����.��%Y�C�d*!x(��ɘb:a1_���Nw���w)���Ֆ�\D�OPH0� ѓ0�wK�P�ӨA�;|1'(�r���/��i�LF������~�ڠ�˗9���6 UUD��tJY,"�aqδ���B+R�!h�7qC����&a���`�?���w�����bm}��o���t(?{@�X0����b��2"�w�v兠^�<�����no���Gy��f��<}�gϞqzz�W+iL��xo���q5*Tԕ0�sv|D'KI�gm�����n��[��ՆO�Q	Jiʲ���'O�����OYT��}�Fk� ��gt�ED_�&����B��Y2z_��yK�Jϑ�D�jU�E)��4�`���Y��cv,�0׋4mϒ3��(Z�V�_tC��{�%�On'm��u���d���Jkkq��lj�Z�(^�̷��~�K�~NW�h_�zq)Q!���Q*�J�|��߿/�����>��C�I](iϕR����ת�-�j!J"�D�х�
ثrt������j���>�B������^��;o��BQY��6��������S�D���$11!�l�Ѝ���c]�u���
7&��h�������6�OO(��t5޽�9Tl,E�>ٲ���ż&�ID�p�nB]�e�FQ7�Ө��RW.B�ί�4�4���\g�'-kG߾łn�����[c2�EkMh�8�[!r�.U`y;糇���������i4���<~��gsn�Ϩ����M�Y���N��O~�3����#·�r��Rʪ��KT�"�߾��![�&f��g�����j���)UU�����������W�LQ:�פY�|1���2^�xy�_Wܺy�V�!o��w~��`���]l��	E�qV��Z^�8���%7����	���m����4>��cF���b<�ɵCD�%Q!�g>�1�Ϩ���ʨm���ʒIF��|��G�����"�Ak���]�Ii�Z�L��s�kOYG��[$IF�g-�
WVL�#./ǔ��	�����c:t;�l��i%}���u�w眃��eI1�9�g5u]3���8���ϟqyYPۈ�4A����
��߿�_������{j��1�� ��ǻ��=�{���7�կ~�d2i���,��6E���,퉪x�7�[G�Փ'O��w�~7��2�jA����?��������@�c��JҨ�vok���G_|�txNU��[?�����N�v7G�h���Z%X�wn����V���c �G���ʹ�Y[�S�\m)˒�dL&��ycU��i9Y5����7ڱ\kJD�r�p8H҄�*�i��I˪hk�Z���5�����>�&�����Lc��A-���i��m�~�ӟw������mv���o���m�H-BR,����$�$"�����<ֹ�O�r��r�B4�.�Y�IL��:��H�D��!��K�����A��������㏿w�(��z��������T.B�^��JI���?�u��fÑ�*�X��=k|�[TH��cU���/�NRҴ�Z��HCr��6�*ߠ�}�_I�Ccyʲ1�C�q_�7�k-��R�S�Yކ�xl�ڴ�4o�e-"v��[]Z�i�am�1M$MS�xW��BՃ�B�f��|�d:b23�M(�cQ�S&�F�3��9�op��>�kk�SC��S�9�]0�g\��P�|�Jd��e�z�*5�?G�j<:���R[����{��6F<�d�~+gmm�v�cm@K�����zLU9jU1�8=>�r�&��6F)��6*l��[���	'g'���,���"�2�&�b2����K����F�}7v;J���3��x���G_0�[���u�t6i�Z�:]n޼I]͗S���#ht-w*q�y(�)Ǉ��򋇼8���<�W�e���×t�5�Ulml��{��ݽRH���*`m��5E1g6��P��Fc�HL	���J`�����wx덷�ٹ� I ��*xt����l@Q�x�����1�$|��M�5/����?3C�    IDAT|Nϼ,�ᐧO���ssg�b>���Grޠ|W��cL��Fm⫨.����kz����~/GT�(A��zO�bڈ�)�^�;N���H���+[��<*(���Ղ�t�h8$	�Ʉ�(V����=4��_�{�[}�9ޞ�m�(z�H�E�:WՠL��R�?-�������ԡ���N�]�>F���_\Cr���W�ͺ��I�2���j�V�.�^��)�t>����|Y�}=��g�sN���!��c��ޙN�-����Q�V�7�L$s�
�t$!.N7��*s�ܽ:�kIĂ�Z��o�# ����j]W3��V��@i�E�м�u�Ĳ�[�dF���I�������[��{Z5�ߡ\"��g.���G����vz��t:=�2XOK�u�.��-0]p92�Wxp!�s���F���h�2��m��(3\]���Qc뀳0�O(&c��PԴ����f���O���NY�������PB���},����$^�Sj��[��hmQ8_���Y�!��;�yA�:X�F�w�X����[@r��X�̊9��/.y��1k�d�a{��w3L����6;��<9|F���5���V��D4x6���S~�ϖ��W�	*$�ה��U��&��D��cs�M;���ln�@�a�\|�/G�"8-�U��P-x<�3�L8�Q5�ʨl��r�cP�������Q{{�dgR7�  8D*���m��6�8����J�A��"��i]�L��)�����;�i����zl7mJI�C�Ao�v��{�#%(cb���jWOh�J������|N��{����?��'0	�c����L"��9�&x��������g|�EME�7����u�t�,n]���b��H���999c8���
.
��5���������+馚Ǐs9R�q�-J}M+4^�&�Z!P�:ˀs%!h���u%J%�uκP�Y�1E�MI����i˟�I=i-.��M��+���?��%�������� -R�VR�O*�[��&I0FW�z]����t��u܈E:�%Ѳ)�_˧��oЬx���9P[+�7����%"�ޫ���߿>��ÿ���[��W���E!�Vˇ��b��I{���X��~�<���k-�%��ɞA��h�8tX����$�J0є��W��#������o���1�
)�}u�DZ7���t^7On�Zln�q��>w�q�{��khӂԢ�܂��\pt��O�����c���]��ǋF���$�	��5�h���e�b4$ʠ�`E�XB5c|�ç�v�`n�ڦ�O�m�r�U��x����!����.OrdYz���{�="2	$�B�����j>�j(3Y%�43iQZHF3��h-�?@f�ϖ�^i%�dM�E�#gĚ~Uw=�F&����p����u�G"�LTݨ�<f�gDFzxx�����|�;8'�Z��y��:�+:���@Dh����.��k"�8�()5�Fxx�KJQ�F��-n�{��[(F��o]��u< �Y��Φܻw���h@�{k.R9a0\gta��I��̳u�*o]����y�i.)K���+b�kc:K�-�R
���p�.E��2k��oq���
�A�\p$.WxӷcK��V\�T%��P�%B64vE�,m��'O1�[��1��1���[����1���ѣ) 8�S�x��)�qC�b��� ii���*�f;����vΚ��T�6�͘��5����_��3��w>�l(�X4�o�\K�r�d�	 N"F[�i���	�4���G����翡��	��5�!�c���QV{�RX	4��wwB�3&�k�qy��!%�@�az8�����i޿˝�>��'�ۨ�
Vrߑf�!���/�~|��Qvw�u~�)W�΋7�n��@]f���y�����2x/�HmLM(lBJo��?j��vY5>5F+�ݵ����O�d�>�� >�����O���G:�����b���+�;�Ժ�lTIM3[�����d��nE��ub!ʏ�Ʌ��҅1�X�R��K�����U����fę@߭���(�h�h��4�XPe���x_�j�[��v	����:hD�JT$!��p.d]�vI�>��ٿ*3�9��e��-�MSVD�$��������2�_ЍkG�
���tU�!d�6�r�*7?��?���~��K��k����^�����m��u��K�؟Ly�7f'9M���p���:��m�>��|;����fF�5��A�jIi��<݆_H��#޻u��Kk�oq��m.]��<��g���K��|��[�M�Svww���c<x���>I��o�BR�U�%�{;�'f��{4�6��������}b�`�$ib|���/͔0�0���֥.\X�	��X���amT��ŷ-�ㆺ�D1�u8[`m�e���0Fi��w�&�;�Ƿ��w�z�2��̩z'�2�qX!j������u���N�o����SNժ�t̠OS<!Lr���{̏��b�!�������*�������|��`>*>v��C��Aei�	�}�k'�lm] Ě�3��g�lS0*���'��<�������,")֮��F�O�9/A�$�~q����}�t����Z�!�-P�`M�B,��<%E4`D�.���1�����1���s�chĄzU��[bPJ��g:�#�Y��I$��ɴ��G�-�l���s������b�S8���Ң�������=Lw��1�oo��n(Ӭ�O�̧G%b�!�j�8Ve]Y#�u5�����4|�-��?�O?���~?����Xo�������9��5��4�se��PO&��'O6�ww�tC�EI����en�u.��E�6`�qh����%�
"b:џ��T�L�1���/������k:5��ƙ@_Bw��H�B��=]~�E����Ӹ�J1�!�V��Iٜ؂+��&EUs�*LgP,���с=Y������������X�SY}��M�:�[����h4����|��G|����z��%$�Qm�M�ea�8b:�Y�ؤ�z���p0�&�U�������Y]���O��6��^��2@�1��#M��$0�3����8�Nx��7ih�7��i�u�8k�i���Jz��m[f�>�W��'������石��Z �^S��)O܉�H�	��=�ٲ�����C�Z&��G�~�d�MJ�%I�D-��{�l:�`o��G��y�W�^Ŕ�<`�����ȓ�S.]�`4rԓ=?���_���~y[s�-�C�%�W�t��<3��9��������;��F%X����Z+m}H���N����.��?$�DU��5��
�;<ԓ�GgL�O�N']Ex���͔�B�ޙDY8o��`o'�EM�F��)����������{��x���6�g�4�Y�+^�Au�?�X�f:�Bw~����Ε,*��\5�ӻ�.c ��ͨ�MTeA�a�k3[ �n�h1��jn��'h�H�"m8Z��s0> ��ԶB4g&��ۯ��x�YM���qHS7<Y�I����b����|��|̅��
/�=+z�X7�	��x��g^�+��j��j��N�)B�FA���$�B�	�������8Wa� }��'|��O_A��W|�O������'�Z;M��ǅ�ֶ�ș�Z[��¬��{{����Ҷ-�ᐶ^tԀ�E2��dڏu���L)�jV�cz.Ѫ�aT.����򓟸�
�oO��FkL/������Ǒ�2a��K�U�K~~�ӑ�ib��e��{�M�����E�tMy�:��X��I˞ږ���o��	>}9@QW� tm���Cd\O�I����0EC��)���eg�)��Ɏ�H��~�ij?~̯~�+�<���o���ϙ�p�|���"b�1B
D��:�������<�~cZv������LC�s�ٳ�,9���f�����p������MӐb���t�Q�&�B�S�*�����=�pv�W�Q&��_��S��Tw]�[���L����s��}.l^"Y�`<e<��g}�2kÒ����gw�.O��gz�K�BU�C!�x(�l;�}�8RPB���f��?�*�)�1������|����~���� _?%�O�O���Q�@�DA\�X!Ɩz6CS��䰻�)6� :E�DDsG�f8c(J�T�^hSM2UK݌��W��!�m���o)6�EI]7�Pж��aN���C��RN���C��b��ռ�p��f#]�UL!��8����:5�K�gP�XbP�5X1(	M>��IH*X7@����b�Q$Ke�0����̅����-޷�~9g�j����]�[�����O���c����is1/��: 5�b�y�W���fw����[�1ѵ6�V�vXɪ��Ŀ[8[��u2����a8����G?����_���'vs�q��?Y�5����?qI�'�A1����4m9>8ܘL&.�,�D@��<�I��Y���`�8�f�����#�N��T%�:��lc*���*$����3���s�U	A��$Uc�(�|��E'�~��S����C6t�Wg.����8�V)�k(V�#���2�޿��8�qٖ��U���~���k��o<��_���t��*�k���f�	|M�cB}H�v�<��d<g�g988 FK1(1����;��1���~������|����6t�-��Ɩ'O�p0>���#O[�3���-W`��6�:�_7��V����>١r�������JLk:��k#�@��hB�p�ϸ�	dm`)�!Ea�}"�-e�!J[�����c\�&ԖH��!Q�1��Q�QڀȄ䧐��I!���1Xk��@���)`�Hg:]O�k���r�)�Hf�А��Y���2�m��bPr��JT!h�$���qW!D�`�v�#崣��H��F���lJHu��i�mZ�R�1B�&Q�HDf��WLYfB�<�u�o�o�{q���,@U�o���b����͆�JW@�L�����lC��l�}�I��M1`�ҕG*�mC@	����{9�|>F��F�9��YK���/:0I�d޶-V���H1��L�;|\��*^���>�;vrn�[D��Q/�$Ĵ�
{�IBJ~�!�XSUv�&L��OJ�X����~b~�㟙���gG�1������V:w�R�ܞ��c���z�Q U���Q�g͠���Y��#y1*2\��qQ�x�X�Or����j�uSծ�KlLq���`/�n���x��,�O�����L�V�q�&��5	�N�-�XTɓ�Ƣ�U$w��<,�Эf��)�m����Z�F��lfk
<-�Xc+�t<�Z�����%�P��w	�RT�v���e���>`K
r�1M>8�*�4�1�3p��{�7f�ʈd*� 53��Sf������}�n����1J���8��!�<��~���se�*1���ȣf�)I)�6?15����ȕ�
�1ⳬ����;�[��bp��J�9Mn�RPtm':i�j��-.�rv>y^U���sʪB"[uV�i�c��l>/H!Rh��~�ՙD$c��su\�P���s�6B؁�C�����>R~}вh��#��0L'm78J�Ďc�1� ��@Y�m�����'H.͏_ �ݙ���EJ����`�J����:��^��t�-�o�!Q0���S����k�':�N׵/1�<g�.���UC*����I�4�'����˔U�82��{D��k�Gl($�^#��WgX�Ou��EP
F4��巏�Pu��q.%%H�R�5�[�H����I6W E�y���\���������7)X�)�|DT�K�f�W�RJk�&R��f���؋&��0���J[��+��O�n�?�ѧf��j�w�����S4w���n���'���R��*�K�1�}%�������U����d�1�r������A�ˆ�>t��������?�Ʈ~iI=Vk1)��)ϯ��Q��L��11)��@���Jj�0Ŗ�%v������gc��U:F�0&%!�u1�d����u�?Z��7�JB��}CU�y���(�������EvN�/?�wqH)Q75�{{f��q�����n�V�����
!t��ɼ[ċb�ZK+������r�끗�*(�"��B�٪Fcw� gW����i�$���V��G���O��8�~��U��*Q�:H�Y�;c�F�����Kg�.�5��O�wf���p��7>�[Ě�K׸������>������I���6�E��m��(T��!������]Cz�0v�XhQUuRu�Y[M7�f6�!�)��d.��^/Y�u������t���y��������^}ߢ8[!�z�=
'�ݚD��d���_�+8�]��Z�I	��]X�8�w�����S�5M�d� ̭WV,Z,I�-W�j��X��+2@��<~����]BH81E�1j��@����!/^dss�A���0�����$3Σ`����O�ǐ-d�h:��B3k��$�:*5��XYM���2�8
0^%�8�����*��i:���y�&��͓�����1W8ۈ��v���%�d�q��GEQ�����ч����_�6������U����pq:������z�O,l<']��'��>dk�謽��dR��ު�쟪�7+����!��)�Z�j�4�l4�N7Ƈ�E�4Y*�V���ŽesW,��E$��I�(DT�ALix���'v^��-�3rlI�HL;/�:s,"9����]��RM�QJY���֗���A��>�X�*@c-�a�h4��+���kvvv8<<̀�Ȃ���t��]ڼ��o��[W/�6Ќ's�O��B_|.�Vy�� ��++)!��*�3�v��\�����A�eA�:(8��������5����?����o��=��~˯;��N0�����4�+��ê*�Y�F�U�O�[8�/[�M�?+Fͧi���TվrՌ~��?��ʁ���w����?���>*q���?�,������U�+_i�FwyjL3S����b+�?J��7��w<�[냑Sgdm0l�1ƇP6���Y]�O��y�^�ڟ�Si�_Ac3Ţi^@�C$��%q8+��ί6���<^y�Iӷ���$�I&�K"&i�����`��;͕&b�nA��� ��a}m@QX��Q9�og��<a{{�}���x)2UE����K��" (Y���>�r���'�������VX �$Yk��9�|ik��׮r�������Ã��2O�+����N��F�����lQ#�pe��>-���E!ar��ף�>�W˓�d�NJ/����4�uX>!�k�$�F�Q��j0��?��sM�j ��i�Q.���p�P����Ц;X�����׳bˇR�n����z�%���vZb\�&4��8w����}W�vW�ߨ��ٌ4���������
6S9*�5�~���v�b�Δ�rMqV\ҤҴͰ���tR�,S�[u���h���~��@5%$t ��@Hڦ�T��^��|����:rxo�Pp	�6%HJ�uH�9ӷ�^~*ɵ�BF0�!"�͌���\���/_b8(�~��Ç�~��z4����6j}��%�b�K������ds�kX'�f-��v��E��5��iU��$B����pĥU��qx����cU�'��42��v���i裐��T����x��_�3�|���q����*Nf�~w��� �o&�������災��qϩ*Ei��i"EQu�z�m�Uj�Z_ۜj�֕E+FRR5)�.!}��	�}��~
��Y��^/�֤Cm�P��G�!<����ڎ��ҍ�{ab�nĢ�k6��B5ҡ	0�n��6v͖���?֔>H�ه�UAGU5�UY�\TM�o�Q;�mx�}�ڦi�v\���(���&^������R�c�6DB�F�[��y�o_�	�ŵ$d+�؈:U5"G�ď퍗{���;��#����"]C��K|��;���[\��"����Gܿw����K��}ȕq1k�b��(��P5(��Xc}4��'���=e�`/[6��y{�{*ٹ�ϻ ��    IDATH��Z�%���鄃�]���2�N�L�T�����Aa��i�Y�TL6}�k��1��'ѐ�0Y�>\���4}��e:���E �U|���y�5^���_�G�"��Ѣ��N�X��DFeYVj��� )�PT�ںn�1�^5����$�=I�`�Rnc���ZQ�E����jU�q:L��D�Vn�GFt+Z�D��tr	�+Q규wkɷ�c���n8W���Z] �@<���:F?�L��I����t:z��|�nKO����{��.lI���FB�4��U�I��1\��~��� �-��i��(`�}�$�dR�6�/T8Q�Ē<��1	���)Pcx��5޻}�wo\g4������#�>}�o)��ި�8�̲)����F��P��������YSO���:#Y��-��N0I��b%kg(��Id��4������H52'}+i�#^ F�bD���J�W�e3ꤽ�����w��v_���y�&��b�{�%215�Y@U(܀�pHJ	��_��E��u���5]S����R�B1�)�!�Ԋ�Z7j̄H� �u4^ ���v]�#����)m�&�a��� �c5O.���cw��/��2��\��-��\���E�����B!M�b�{�F�|��?8g��MqЗ�>.�X^�d6E�PD�pe]W N_��wOP�ڳ��FM�2\[����*�!�W�)x��w������7x��U���޽�l?~ȓ�;��I$�eF,���	[qEE�F4m�(,�{�ׯ18,���|��_�gUU1�L(\E�b!��RG�+��	�ʕ+8������W0�1�\~�׃,�
  ���������r��Q�ٓ�2 㤮"�������<�D�wg�A�	���q����}6�s{���,Kʮ7o۶�I�vZ���/�����糂ھ���kW�ɯ4��L심YN)冚��Wg���.8"٨:!�h�����{ՠ2h�j*�"8gP�2�Xi�/$R���V�zM�Ψ �
�*;�ͫ�%O�����P8�jJ���0�8��l4kf.���s���ׇ������;�eM{	UW���}v�(�K�l&�>��\>)�}0���ӟ&�����[gb�Jk5U���%f	��Iz�>�~�㪪HbH�-iC.�غ|���y�;�x��UF�����}u�P�5�]�_�N��j�blژH�FL�ŋ�q�m޽q�A阌�9�ߧm�DB��ш+���u�(�BdPX��u6FCJ� �L'�L�����1Z��	�t���fiۅ,�Wo��t�LC߲k828<<<����8�}.sx�at1$r�a5��<��E�)x�Z�h��(E�*I��S����El0֥���8��AEDEcD�dj��q��)]D-�4u�&��!�!�*xoC�4�r�Ƌ�u�S�����Q�1j�Qb�x�cw�)��MN^���`�ٲ��ֺR���}A���XN�������!t�Ƹ\�Q�z�&|�޹q���!m[s��W|��_���}f���a�D���*�������n��wo��kW0ֳ�󘇏�3����1FhB^iI���GX_��z�*�/_f}mH�3&��1��H)��p��/��=8�Mq�r��z�
����8~9zV�(���k:�3�Fͼ���~ Ů7�t�|�ShE0�řO��[�5bR�)*�@JEU4�I�Ģ�k�.�;n?+��EPє��dU�A0�{������p�{s��߿��Y?rQe�;���\��N�<ޘ8�{\�+���M!/uu'����5Ε`
\5��[7���l]y��2LǇܻ�_���ܹ�%��!)eX���	\��� SW�+��pĻ�����=�~������{<����l�%kQ��I�jD�ź���$�j�ƥ�Wٺt�����a:�g6��O����g�!���P2�v�v�V�|��Y��x��h5e�c	�'�E�ӋS���X>7G��]�����}�CU�G�f�y�Ҩq��������+FZ�5	�$�FAS���hcD-�I��,7�l2(J��������rG�|���ӂ�ש��x���`�1�<C���!�կ����gf����RKnM�]A�Iz���j��h�(�؂ \X����~�ÿɥ�ˠOy�����_����<y�M���j:���C����9�5��ܾ͋�����ryk��-���<|����'���]���U@=V�`�)sJ��`\6v����>�Oi�Iw#�\XqV���g��i]l�	����c�oE,�{��ih�����ى�П�k��+�����-ֆ���;Q)�B94�1�5�1-��`:�*kr_�Ō�<�Dke��]���5�B�V{����^���sm���?�J�"��:1�
�&����˷4���5��j"�eT2(S<]�]P�P)%bR\Yq��M��}��Zcw��|��o��/Ν;w2���PK7X/��ՕZ
g��իW�y�&W�^�,�z����~�ٴ��˒f1|���N1�`��Rĕ��FC������d�����b<U��G��J�JZOڞ��{�}ľ��w��}�D�D���g.����)�+ˍ?��`��YW~�Z�1�3,)ET��Z;�Є�[P��<.�`qe,�Cմ� ����~r��<�e��ke�Ln�YΔeiLW�e�I"�ꕽ�y|��L9�*
ߚ^4yU#�X�dR����EE��X���L&5o��ۿ�����Ν/i��c�
��v���T��\�����n�s��tL&���=�7��>�i
k�{h�%F%���Մ�܈��%�]�εk�p�Ѷ-�Ovx�����pn�g}	Ë�Az��㟷�J*I����������W���X��	�������%D�Y���[��3K�v���8A4�l.߿��x_�C π���U�a�x���}Z�3���{��&vټ�M����9 ��+\��a��j�M����� �㍎3��Y�)C���J�b$:�Ϟ�c�cK(˒<@�d2k�������9�?`4d����5�Ic�����[ܺu��W�������Gܹs��;Oh��Ҭe[c(�2�#�V��x�"��~�o_�(
�Y��M�Ǵ~�R!� A^A�9���j�3}ov8����=��nguss,����e�y�=�Nd?�U�K_%{�u���=���m����Z���.���4����z�ε�0Z�I�}ǹ�,�g>��8F���8W`l�ֈ�5�	��@��_�}�'���8��#$I�Ĩ��Q�ѨI��6a)vb��� u�>��B_i+ �S���&�<^��?=���m��wvA�J*¬��D�x������O̚@U��쀠`�a�q��[ܺ�[�(�I�<����|�)���S���`��QC�<X�X���Q)����*�X_�k�����/�՝<�W�]E�Y���t���a՟�ϼͫa��������S+��x8I3 s�`ur6s.u�������wr��<.��f���7�_s���v��'E�w�y��O!=+������7�#�d��ǴB_���cN2��O��%F�U���ZO�~������IX�-tL�v�M���Ο��Y��;�,�Wڑc=p�}��N<[��2>q'�I H�\?��7��z�K��)��x�^�[#��-6�礟S�T}V���f�g�2���Y�>�E�j��"�=�G�`>/�Zͯ����[f,!�ު�tm}��f��pΥ)����v�j��ε
ߢ����'PL���|���*�����}>|ȝ;w�]��SU�gQ+F��p=�L�ommq������u�666�L&|��W���?�w[!���tt� 1yF�7o���ߦ�*���r��]?~L]��f�\�����߆X�p�N���~�-H��y��=��޾�����ZyrtBx,�|F%���O��߅.^��~���=��n�>���Ua����[|�c��҆E�/��U����M��,�_g^�Ǖ��� �ˎ_�;�qΉsN�u��uZ�����������[_����O��G�7-F�VEE� ��r	�Y�}JJX^]�̩�+����}�n��'hBU��!e9�m2X[[���?�>|�ׯ_�ãG������/x��q���ɫ��Bm�^�o0�aL�h��͛7y��ﰹ��d2a{{��>������4�{�@U��6�"s�on���e���Y�d����X�L~�3kF{;������߱[��a�Dt��Iz��d����㣽��n҂e�N�!��g[�*�}��l���&A@���nU㉠�E�A���Y>Þ/�c�AO���~�o�?�	�y��q�Ӥb��eP'K��J�w��V����cL""�\a��1Xg���f�{.���;��g��ŵ<�%��Ր�GE����VTU5_i�1���
�f�F��v����8\�(�� ����&����G��7or��E��}>��s~��_�t{c�����$h�%З'����Wʲ��[����y��m6/l�t���`�����Oa��sߞ3}G��ۣ�^g9r���:�*�B��(_o������:H�Dn�t\ ��|�G�:"$zI�2"�������j&e��벤g��N���.tvϜ�%����2sܛY��+ow��'�Ó~}�ذ��>I>Б���2��S�����e_G,�w1;h�􄉱��9S:�ֈ�^ӌ���'�g?��Y���7(��������kn�E?�b"V���?���aޝ�B�Az��:?I�H�m�1�N�!�u�oB���o������;����ŋ�D?~ȧ�����/�~�F�*���ӗ�ж3���ck�"7n�`mm�m۲���xrH-�r�u��r츕ٷ-���8��g�o��W��93��m�Ukw,_kk^��<y�Ư׳��������g{����ѕ���u/<�f̋�N��%3��9�*��%��J���LO��=��;���<����q,�i�(���Eq��x����z��獛}���U+�Vމ�Κ5��5�����1gouߠ8[�ݢH	lJ�`,�d��|c)g�5�{�s8W�W�ٳσ�&3��^}���dp8��p.�ԂZ�p��%nݺŇ~ȕ+[���y��W_|ɝ/����!�� �ퟮs��|��������?��}�֥M���p�����rZ��x���m��M���c������� �\����X���z��"�x��BT>?h��$w�:��L�gX�W�<���3�)�F3S*Bf�̢�d���*�3�ǧ�O�J>(DMWh����J�m5�������~��p�5�Gu\���ī`�����^��ιcu½��/ɋN�2~��3}=��3} )%��.2�IuՕ�!�J_���/�E�g�g��
<�oz�	���|�.�n]c�4��5������@�����v,�8.���F�2/�7�t���\��1��Xm����p8dww��0�����f|����E~����e4z����~��U�i;cP�q��{\ڼ��H�6̚)��!�������]�dQ��%z֖ q\��i�h!�|��&n��8��K�z���>ޕ8���h�:�x��ǂ�[-�XT�0��^?�>��`�?~!(Q��,���*^���4��o�xn�����vL�1�9��@&溾�LW���@/<���7��5͋Ɏ�� p�ƋX��|?�}��3��2�{��nk��lB��Ĉ1QL(4�ʵ�����y��ę@�A�ɉU�D��"�d^�:)y�������u����z�*�������s�c]�]��bTK"֔T�u�p8��W��x�ob��`Pq��%޺z��]�^7��)�lK)�A��U��>�����_��_��w��`�x����';s��=�r���f?��f��:)��0b���q���Y��*qV& =�͸�N�xFW��
0����XT0ϋ����Ed�0'k��V6јȋ
5�=��~�Ȍkϼ��~��ǅ��9��90[a:�/�u;�wʉ�(����۷E�`0�,K'���Vq�)��y|�����q�����q��Ό�`�w7�ɈD1N[�$C`��r���{�3��ٺVZ��aJi�.���b4�{����2��_��'�bLs˓����yY�x��������ܾ}�����r��=�nr�)��*��[J4	Q!E!%�A�d˖6,,)$��|N�>W�Un�|(s5�&8����o�q�-�~���i3f����Y�|��OO�SwmI��~��
,L�v,*b�-r{&���������q����o�3��ߥ���TP�2�ޓ�Q̯�����:4�4E���}�]Q�l�_N8=/b5D�6ʲ�G)�:k��Y_��o[�FՀ�t�`�(
�4�(*Tc>>���!$R
�k��q����٬�mg��e*Wa
�GЀE���!N�X"�f�w�p8�mj��2�͘M'�豦�үB҅!oǀ�����%y��My��!׮]����?����u=/2��)%B�\K/g�?N�������|G�r�`+��:NwgN�W�uW��>�s���x߫�a�x�[. 9��{�Ngh�c�e�|!�е��DD�X+)E�օpoc��9%�-��i�fE�d���f)�&�Z�^D�r��Z���d�����۷y��	?����������"�7BϞ�Ч�\'@�H�!��	I��l�Rpue��?�ՔMl$�ّdH�`PJC���q��gO�9��#Ƙ���G��ٌ�F��⌥��X�4&�&R���!	�*�2�̍�B@K��A%a�+[QC�<p
T�+�d�`l�MCUX���/Ė���p��0&���P�:B:�.6_��A�#�,_(܀�j���W.1(]�ڰ����A�A�.P*)�"��#	V�,q�0k[|��x����d����F����t�C��p�2><d��C=~�ݯ�dg{�Է�R!�|��m|���{�_�N&=z4����<�GZ��k��}��܆�cY��鋗^^.k{����}�_�g
U�I�y���)�0)xx��b�ř@_;D��+*��;�a^b��%-m�.tƂu­���C�Ww�`{�EQ�������Kz�QG���&�������RV�M��W�^��$_Z�,n�UJߚRW������ɘ��`I+=<�������>m,�����6`lg���5�ѐ���J:�)�Õ�XT@c"��E�G�쀌���8ہD7}$�u1�� ���	!q��8�`I�����pPRV����䐃�]��'��|2�F�g�k��$��Z�ZT#I-��z�mnݾ��k7ؼ����pP�֕���iIE��4�.��*)F��Ě�l�C �@���T�ӥEQ ���T�m���Y=�+L�Ϧ�v�{�����d�`�z��2�t���O�}o_�������m�+,q?n�)��q�8
��_)��#����8fO櫲���{��y��V阽��E�ͳSG?��N1%IIŘ�ˈ��%�ŤP�&��s��-��߆�Od�׿;
�fC�j�>���8z#/?�t���{�q��E�������]����={�c��j5PUU�t���3�58�0z=N��L���oy�fm.�*������{�r]�4j�V��|ٳ~�q��I7hb0�@�E�ePٺ|�w�y�˗/�\���81����`'S8J�8�N��� &#*W`
Ga,�C��R�v�
+�Pƹ�bĊ �RXK+Î�2�W��1=ܣ�M��_�����3�ݽK�	c!)�W2鉭>������r��������K[����&
+�X'x���dM砪OU/�[[�����l>ى0�-X����Sȩ�r�ƈ��d��c���K&�CrEr���ު/�s㸔~ߝ'��q�ެ}����.zP�0��;��X�[8��yR�g��C�`(�b�Y�:����~	��Ԉ"��1u���Ι��<�aq&���j�J2h���Y���S�g���C�����6k������K���� �� �o�DoΜ+��Nu�    IDAT�~b�t��-ȀO��u�EG�gW뫃Mh b���ƐR�Z?C̳��E����:�~�cy5�� Y# �5�߼�����������¹��Y��0�m��ӿL�SЅ�����K;k�5�����93h�d=!BH�	p�r����e!(-)��+���3(+�z����������}m�C�؁"A�d0����[|������w�JH��{8��$c;p'���c{V=����wk��T!%Hm���&��,WR^�AE]�L��y�����$i�$�C�D9�����f����n�Xb�z x2pXf񀕖��鷾S�r���o~�����х²Fo����Ξ����>�{��)�Ŭ��󽐀F���ak��oz�q&��xo̚؂�u����E���X˫�eEJ���ڵklooc���*��)�锭�-��X�#�1��~�%!�Y0��������7e.� �~G!���I��D�8︐o�g�=]��9��2�e�Rg�c$a�8Z�;�}��?��ܼ�n7��-��&�0����w��$���~k���|Uf��ɶ�vђ@�#��2<7m5�� �QNhX ������dXMK�\�$�Q�U���s�#{������dVeuߪY�d�s�9'N���X�[���8KflB�C���`|~��?�c`D�T��1h��D��=](BU�)(	�u�%t*΂�w��!?��S�%�m�	�)�yۥګ��H�J�Đ�3�pr�>�l���ږu۰Y]��\a����)gGt];�],}uCUUx�ǂ��9�v�ۢ>�FXT3�K�,��ߴ�]~�fu���
���r�{��sr�.��,�Ec�Z?��9;A�D�u�İo�>j7E�4}��4# ���_�M��LGz���ϟ��y��@��T�=�g���@	U�mۑF0 ��V�?_��-h.3c7WWw����V����f٭z������3�EU�AS�2H�w���)��r��M��?���DY����/�3�2��j��A�&T���ВĚ�B?p�y�ܸD�0ҧ��$���B��Z��ڍ�����Ik,V�3]�wb4U6��ng��{c<<�*j���ܽ�wN��\A"���-�͆�=.�(�|��E�DM��.Z��'��ɳb�(xLヨg隖���eg�m�����ق��i�5!�d.2�g,Y�ʲ�,K�ީq81D��V�k�t<���6�e��X� i~Eeuu�'?�	?��_��ZQ��|�l��ݎ�n����iƍ�9��n���u��U��m�^������Ȭ��v�_^�ێ�m *�|ƃ{�y��#���������yA�X��HBL�(ߐ�t��~}�����4U6�߾����noo���2ӻS�~�y�c��(�1��nԑ�78���c�}�ѽŶ֎Ǹ�M��a-�1Fڪ�1�M|��wX��"�ҧm�g��ɒ����cdou��m�VUE�e4MCUU��.(˒�(���O�{�xæ�{���E��l0i;���'nR�7'�(�L��5�C&tB7��!!�q��Ǩʻ}ᛲkW��*�O�Ӭ��eYZP#�UΫ/y��%O�>e�^�c�\2����}H�գm{�lY����� �����v;b�cZ��:��I�SeWoi�5yn������?�Xi|U�!&�k���"�6�>R����(m�u���:ʲ�w��}��������3�2�*s\~��n7��*�2�����2qз��Ib��뢌,yq��8kH�����sN~�GGG\�ڂ��W��w> ���/��/~jbS�g�T�s(0�w����c���&�L	y�����l6c6���y�!�}�@fzb��X?$|� �Z�EQppp���"���%��_�6Қ�y����V�������l��e��l	a�FC�T25Q1� VL�$�F�l�/`��-�G�)��]��0��-�ŌˋWj2�db��M为��u�!�	��O�tp*�Hw}9�n���L�J�l�ح5�e�Պ�jQ	]�fĘ�֊�%=��a�!xBƔ��"D��;����m}�)&:����Q0�Md�k���#\�!MS�n9\츸�S������_��/{��"��Ξ�}�����ꞣ���@`l>0q��آm��)�G�T���l6�N
\~���.}tD��8>��3���M���"˩��3���9��T��Ѭb�
��c;f�3*>%^�	���Liw�t9���)���eH�t���D�03<�4#ֽ~�D�JG��iS��P���q��`�6��yEYΨ�/Y�~L\,���[�q��_=�i���-���R�O�D�Z��a$ �� _�ٚ�l��k�ը�ٗi޺%o΀|�N��e���Ƿ����so�o���ӣ#%`���"��c6��X,F	��븼��*��?ZyVrx�����NNNn|��޳�J����w��%����9�l���]N�RP�Y,c����^�FJ��������wI�<~��jQI[�.}ݬ"y��k�B�M��g����r)�ٷ�n��8o��jL��AEzd얛�@��G�T�s[�
��~������&�@��B��zE��HfY����nǫW�X.��y�l6c�^��hQ�F���cS�\G�M�pvvƿ�w?���ǜ���L�=�����{P%���C��I�)B47
5RAG��>��&3��:T��A#V�lh;���6^�z�j�����+�&vTT%�_C/^���v}���c�5j��	�?�,�ą��"��}e{��9���1�Rц���3d����?��l>�mClH�ж5�F��L�k.�/�;�[Q4M3r��|�]
-`�皻�K?�u�z������r9��<y2�?�٢k;88�v W+ EQpxxH�D�躖���1�$�4�ۮ�3G�ٔq(���2�q!Fc��1Ħ���:Z��ڭ�^��a���(��g�F�og �j��5F	�O�e9�U��O�Q����URu]ߨ��3l����T���1��u�͆�,_C ~{���m�
���c��gϞ��9�g/�!�����0�`��`"Q+�S����I�����91��V.z�`%K��%����h�c h���l�k:�`L�EQ7��5�5L:��b68}�MDd�V��7u����U����:ɹ��z$���d��63dY���1��y��[C^��yI���w��c7:|o�K}�����wk��g����T|xn�i����'�s�{�= qT_�z5�iV���@~ѿ�$u�!�%���,�'��!z�vsE�����bD�{�k3�&�6�=m���4eI�ACZo�Z�ױi�X҅���,{�Ӗ�Dxxg����wYU��tƒ��T���״&ݻwoD��-���!b���$�O�~�������n���n�b����HJ���M���iޯ��?�E��g�=�vOhۖ��3�;2�rK���x��W�&IC"���\z1�yyC[��܌�3�#��[�!���,�r��$�#�8g�rK���}�j�BO`z��a7���C~*=-f��,�XT)-�.!�m��5�> ���b�YƤkS�{����ϖ,���������3N_��nT�� Lc�o��eY�/{��%��1�Hc��4h��x��c:��N�8���j��}ey�>�I_�m��)]�m?�R�u�޽���GD1�gC�)5dYJ/�!��������� d����%��:x���	�W�{�5��j).
���������;��[o�r�N�68c��g���*1�[�H�~�P�sb�cg����־#���AlBp}M�ZK�&h}�\���V+b��e9:�������Y}gߜ����AJ��u�j��$��#f�� &B�l�:IKB��Dl/�# mDTq��ӴhD��p�<�)
�ҡ}1I�4|v�&�@�j|��f�Q�@mWՃ����yۊ���;������]�α\���}�sBӱ^�i뚮kGt�,Kf�YB�eH�����Pۓ�]�s���#�=zD�~��r~�v�����g-7Rh���;{�y�o
{LQc%���v���?��?#��f��
�<����ؓyz��ƨ���\B�CHE^�md��b���{�r�d>���l��j��wt�����	t���JK�F|װ�l��ի�^���jeڶ�U�1�"���ߴ�s��|�~�w7\]�����H�zo��ŝqR>>~��<~���7�?~<��?��c�裏n��<~������e�gv��a�QA�(j��w;ޑs.q�4N�p�T4L�餚���Ӷ�f<M�0\�N߳\.������|�ޚ��#Qގ�M�9Mͼs��y�"���b��w-�'�*��Q�ۤYB���GQ�HJ��Mڐy��?y~�PcZ�1��ƪ����rpp���)�|��NO	�ë%F����!t�\��؃[����::����\ڷa�{c��n����,���p��14�=��9UUqpp���!��h������5l�[�O��y���;w���rvv����&��%�J�e@�Ҽq߬S�M۔�2�wH�W�/�N��S�n�������l���Ÿ~ܤ8��=}(�@��8��n�_Z�25cb$�@�<p}?lgm�������W�5��2c9_pz�k3|�QgK���n|������y��v>�}�C�1���U]7��fS���Yu���V�������ݝ�鳏?���9|��G�������g������Ţ��=~�<~�8�'�m���u�e�������Ν;���ivQ��|����޽��������#��n��_�f�7���Ǯ[�_��?��r=�1�g���V�7��3�ϯ���.OO�Ν;������?��G������ӷ[�c�\z��0�p��(��Sq�����S��w���$N�3gpʦQ��Ѿ��n��e��'��T�,#�k=-#Bf�3�Y��2�K���]AL�!����	��Ȋg,wf��CUU l�k6�Mӌ�l6�ZKUU|�;����1��?�)?��QB�/m$�X��M\f!f�eNQdI�y�0i��.������9g�HS
9fdƎ�5�Z��1�W.c��sxx���]�,��
1���eM۶l6..V\^^��/�dl6>������y�=e1c�7c �x}f�Q�o�������`{�k���A�|>�9w#m;Eꦭ�Pձ�p<�1]ō�6#�eΠ}�zP'X����u�n�����ݎYYrtr¼�(r�s�*X.�{�=�+	��{���Xجa�3�����m�H�F��2�vm;8n��X�t�ģ��Є�;u�y��k��(�J��y/��$���h�����;��]8(�͂�My8߬����Y�i��E�m�����D���_�W�a��޺��f;��J8V;�{U����q	pڿn>��O���v'�[���Ƥ)�F����ٳ5����QY�f������w�Т�,�F �ЃI�]��֫PF]Gs$&�F#b�.�5�|�
�nr5}�J�h�0qI�,�vW����m��*)v;�c�U�pJ���C�u����#��>����sk��ιxvv�
�z�O:�R��h4�)�u�:��ؠw�����N^�IL��i�����������,˘�f8�n�o�F��}�q�\������kS�}P��T�������(����w��x��W�%˃��,�ˤ���|NUU��\�s~~�f�D�w�y��}�s��~�{��s>�O���3��Qr��V�^Ƈ4S�%���0:g_E��m68}��5���!��Jz�\Qi[�v[���Rf�jVb���9稪*��B��[�&İ$#xO�D�6�B�Gc���.��!�?�O��ǜ�]�HUUt݊B���f����&��w�E6� E1��5M3�]��ƈ���m[��-����|>MӼ6��E#���=X�4]�y�(�����G���{������#>|HY�����](�G�wPv��H�O�I4��Ū+=�_Ί��6Կ=��e�Uӡ�klB�ľ7�ZQ5ǉL�ƴ�Ĉq�U���(�5;1�V�.��F3+f'��,l4���D$X$8�A��UT�ݖ���HMl���hT5A4�5�v���fp�ҸZb�]yﵫ�0""b�����I�D]�z�g��%���:2o�ع�Bv���D�Js�p�!*�TH�M���K�F��f����fM�	Ar

�QP0N�yI�1I���9�s��U9���LͽJ�.S��Nb���Zڶ�9��J����=[����a������M��VN��ё�"��,DAMT�FUׇ݃ߵG��S?"y�KS$�3?�|��fLqu�'�_��5��?o�*+��kz��?��M��(�N�(o� d?�<=����FUӁo��E�ݝ�7���s~[��mc��ɞ�����3�#|	�-�kgJ(X_]1�9��9!��6\]mȲb��ʲ��|���]NNN��"��("4!�-(燨ɩ�m�qx�./_>��/���w����٫Wx�R��m��&�,�y�j�Z�?}�_1lR	Ŋ�3�!@����ޝy�Swqԥ�+����|�٤Pe�������]ץ���yY�u���"��(�˄��,G�py�e�kX�.���e�Г��o���Ֆ���@3Ќ��gcZm�b����.r$�<U�����%v���u�r?/g���̩��N�����N�������~�/׎H�n�%[��Z��x�#�y����� ��M��#%$�4���f@���������~����srr�Ç9::��@w:{y��t����Z�+�]�|���a��h�]�_^#���
11���FL��J��0b�11m���9uY�5Q�!Hf]$�Iʈ��� ���!�����3E�r�X���8��:&ؠѢ*�˽�]�dY^;��!�1b��ykmK:�`�M�mTTՅ]�cn6������	��jUc����D��ֹ����NUQQ�>�����i%5� jhDE�u��X[���:5]1�N���}�e;��Řh1�d�S���Ҫ��l��Ζ&���Wͮ�;;<�7�9�!�+3��u�e6k�j���������~�O�������5�o�@*Q��bT@}*ݠ@�I���.^ב���i����y�/B���T�'nH�"���Q�e��iï7u���OӖ"B��d8[�1�O#�%x� �A�\ˮlYg;|��
�g��W��@W̉\9Ǹ�g�Ny��W���6qآoA������1Ό±�9�.	['_������&��S�N�I��E$z��M�qxxȼ�06m�����n����kܮN�]V���'-Mo�\*r���W�����9����?����S�#��+���!�v����e�t*{P`��o�1Ӵ�4 ����o��:�y���c�n���!������ܽw��?>����|�ᇦm��ߋ/x��)/^�`�ZѶ-�k	a�:ٔ�*�$���ը��V�\�;s�Q�80*��x�J&J@�1�Vq QP��W�8���b��F���	^�rk�WBhQ��q	Ռ��n2K-֥�c�P�N�O��K���Y��5	~�C׷�T���}x}���m���Ö��*
EC$X�(�^�k0�͊�	A����2'�K���D4�BX7Ω�A�s�Q%FED""Qc4.˼F1�]�fm����La��f��k��<8yZh�c�w��3��umϲ,<���{�����������_��g"��r���rG�d�"�D���5Q}��N�0=�yD��?V}��u��7'ؾ�"���h�n*��6$e�#����۾Y���ĩ���O�����"_�l���X��"6-� �q��vӢq��6-�GK�,�f��>v��nP"B9�Q7���1����?pvz�v�P��w���� ��*(�GJ���ucRAI�:d�^$i����$ۍZZ�a���޽�F�e��f�P�%�K�'b�46k�@���X��Ҷ����s�뚑�:�?;�ɧ��{v|t��W�\^\�Q�?A����_���w����3��uh�o�L���4�3�7E�޴���!�5�J�4���;�-��?�GG�ѹL���cUU�m}V�Q��    IDATo��V+�?�ӧO9==e��"Q)\��D������Ԣ���Q;���+T��!*ɿC1Fz=M��Bc����з����j�9q�I�� ��	>`Ħn;�K뗵L�HU���1�nHE�&����±�w�J��1zBPp���*j�WY � E��@�j��XL�R�V��=�c��>!�"XcG�NH���HL���t����� �Gt����::�l�n��� b�GI7
C�X�GU$�2(�f�2���B���lV!F3�nU�s���ф��E�$�>{�������)����ݭ:r���uf�UjF�"����D��V�.���}K�µ0�t�o���C���������L�!��&���^�����42��T[K���,*P��E �@e��l������A#����@���#n1#���y�:�Ѿ3�Ř��9�S^�x���Wt��g�o8��̐;��\oi6M�v[|r�l����ٵ!�lL����}�o��9�s||�G?�pQQ�9���ټ�	�7+�%	}A�DM�I��ƞ�\Q�I��NB�EQ��S��� �H`����=��v[z�� �n�՛�~���?�toJ����Lm��,"c����>��C�����w��l��IloBTӶ����l����'=�a�z�S�����;���l"�b��R1�1���1!
1$�I�������1d�%�=�!ɤ%~VD�`\r$UQ�e�z�'��R�y�6��x]U%�y��\U�_�3Ϡ��0��u)#��<;�����۶��U�����`��%.'�]ZK��I��7�6�X,��QK�$�.l/�o��q�#���)H�#�Y�3 bDpVȲM�o��\���.#�G�;��NRp��Q�U���,���{Z�Z#�m���A�U��E�a��hu���+˟֮�������ӧ�[:}���j)")�TS�a��`H�nzw���+��_r��|����x����}�E��@D�O�����ЫwHߛ9��ocS����׶m����kG'�<z�}��>�Ō���2�ȋ
QC|�ֲ���5D�����8�XɈ�ӵ����W/h}ǃ{w��J���\UE�#�~_ץ��r��pq~I]��e�s��"�or�n8Q!@�c���~�*����C���!�������O?O)h���;��T9]w[ʲ�����y�3����w?`u���┋�s�֗d�cy0g�I���t��;{g_bӖk��=;Ӟ�S�ox̀N����5d���b>���������k��k�����t�3޷�Xʲd���牎�bS�D�P��mi�Ժ�w͘�v�Z4ڸyTET1�H�;�H�{G��A��W��(�'��[*����c�b��J:N�-�mI-!&D��_�D�5t����~t�Āok����it&�Q��?ט�®k'1F�bUN�<!v�TK�54J�:U�ś���8:"VA=�D�+0N� #DA%�XR����)�� X�I�u$��78k��tmHWbr��]K�Y֑4�u�6uhR�wl-bL:�oO��ɜ��Ǯ�|��I�y!�*bT����w�l�\)aU��s��r+�om�:@��,�����)G=���kT�!�����GNÄ3��k��-������<��S6���/�h�vTr��6]0~�׿������q�&Du���E�&�����8>L���ܻ�٬�{��1�.ru����n���1� ��$+`�`l���F�6Pf����.M�c^��+��^^D�4��l`躖�z�sx<EiF��� ��oZ�n��z����b�����<x���lF]�\\\pyy�u2rc$(h ��������'M��b�ɝ��*��O?��?������uMYe,����e�o䝳�m������q��=�{�f!���k��s��y2���s�ݻ�ݻw��Ί�ԫ�+��ù$�rqq������zX���Eǖ�0r�� �wF�	����9푿069� ����8�O��Ǻ����9@��e�	!v�~�!�{��:���@�u����@Q��5�O�FDL�H�9Bp=Zx���'�SJYBķ���x�1gm��r+1�H��!���&�`�D� ���1��D18��N!`A#���TH� "�9m����}.K��	tɡU�RA��)���c
:�4u��E���֊��k%7^M���/L���Q�u�uB�l[U���?��?2�J��_FUU,���TS����熿���q����.�}��#��Y$��$�v�t{��	��y�o����z��u�:1s���brH��~���y�	�w���T��\�k74�������@���=����X�E�`1�ٻι\����3�N_a�b�z�d�Źl,�0���dGׅ~&�/��u���c����}��Im	����n���+v�K|h0ɲ�5}Sy��Al��+˄V��Md����%WW�\\�%�2"w��a6/��¤#���;�~g�m�Uy�c6��Z��9���,�>}�ڸ��}�ћ~k�(�N���u�f��x�����L4�>C!�o78�]�h!/��~D�i4�E���2K)M��b{dӆ�'�T�Oȓ:))c!��	�A=��	�2V1�@��X0=�-e"ҹB��H܀��y�-�әQ=F!�*�IB �"!^#i`ȝE5��U�I�T$�J������Q^��Ū>C�������t�1H���}��ͮ{���5�K�֌���ǙaL��#y��|O�a_Je��з���H��ش��kE�����Jg��$D/Y���mp�ʖ!/Y�����:��<���5�}OU4�$���]#}İ����_w��& �O�������ސ�"���*��_��6ٴ
z��~]�0��ZF���@��lVr||ܣUk�f�fs�z����ݶy^bm�t�&E�=�Y�!:��i��*�(E&, v����ӗϙ�f=R��;c��'�f.Oܕ��ӵ1��L�;֙����q���+�>U�����������2�I��Jfe����w��O�h��̲Z�X.�TU�ԑe�횧Ϟpyy�'�|�j���'�����(R�|6+�w���:}?�9���X���~��Mg:�c�Z�l6��ݻ<z��}��k��ӷ>Ӡ�,˱��v�5+<x@��R������ *�H�ԗ� U%�^���`�s%#CA��%�D�����ñ�Z))%���(�Ӎ�؀s}#��WC���Dm����������'��W���i�����G�ff�Q ����%R�Qz~�D�I{p������{��m�
Ltt�?ǌ]� �$���\WYw��Y���E<��8��~��)�Z3:s��er�D`�X }�i�����?�8��EY�g�o�.���&��eծ(�:������ό��Y?�����ٟ�ٟ�.���J�ʕ�]�ԵA]Gɦ�r"��Ut1pqq��ppp����3��,�����7#�c����!�?��2�h�%�6�T�c:B�ݘ�S"���5�]�I�_�1=���M%ZTu�쫪��t� :�~��qkR���Q�9�W+�(����%.�8>>�Y5�C�����wPu�OgO�c�h�1Ĥ>ف.M~c0�al�n� �:�EL�䁮k�tI�uc:��̲↰��F��K�Ǜ��B=���BE1Z�S�i�bT8樷��`��eX�"��C���6,fs�Y���9�����k./ϰ�p�H���}�v[lY�-mӄ?<ZR��M����sv�WW���윧/�\�J��|A{��/W4u��Q�a;�qii�qBQt�c(ˊ]�b߀$O�����_{H�"��T�)�2U�)�Iʹ�'�4`5"�������5��N����]���ã9���E�'F!XG;���?��c|�l�5E�H᫳s��/ħ?��������n��a��k2�:�.8t;d�
�{�*�n:Z�Ĭ�n���G�*@�$D�د�W��:O3o�m���_.���Ͽ]�T�U��w��?����:Y;��h8;����o�#%��-&z�A�T2:brB�W[	X"&v=��}�,K���m��|��/^��,��ΑYG�8C�
�،�_����U��bA����1<z��|N�u���s������%���ylϰk����(�T�d�X���Z���+}���T��y�5[�U��!
��d����wԈo"�$U��H�q"i�	�����z7�A�92w���t��9�~����+f�*Q2d�&��@�Ћ��y��ډ)Ö�*� �'t�=��������_ЈnS�u�	�"�Nh��8�n�g�q��0M��7,Ĩ��WW����t7)*!]{Rv�ZK�K��&b5�������|kC��4�3b�X�����U�y��*ۧ�=��;���=�����r+���͑9�sng�e��7�?4ָ���bq������ܫr||�n��'?�	>('''��?��Ç|�;�[��ЦJ����f��>8'�A%r-r�����O�"���(�V+f����5a̶mS˜/5C��uUUq|rw��l��5�1de��b4�yvcQ��&UI6)�����4"�FޚI�J}z��K	��!��}&�]��6p=��sT���O�<��'ed�&n��Ʊ�D�e4�TM�׹a���cK2#��>����3^�xE�4x�l�B��������w�4���PM��Wu�SN����N��i����yV�>��qyy�RB:�$F�r>C$����~AA7�o;DW��PsN�v�<u�i�@��fGizD3"�6�a~��:���s���v|g�1%����D*�jO��:ƧGTԠ�;���Ħ=�m�)��(s��Q�A�y�ٰ�6��f��?E����}$i���ck�A��իWq��=���z̦
�r,�����M��6���qy�bWo��u�����9�>*1�^��5�RV�Y�o�njb���Y�(1�� kՈ�h�k��"j�ب�ֈ�tm�����.�� &b�11F%��Qɫ�'�1VĊ��%&�;l/�"Q�=�$�b�%&R,�ԀŰk�t�%�kɭ%K���m�c��#�!�M�PDERn]DDQcDȋ�!�:��V�h�ѐ�� ����$I���DMH�pbF���(z�F|[L����<ύB�#UQ�n6��ƽ:�l�3���Xt��^��f�uu�Ύ�Pxa�絬Vw�����>4��#w�]��Z,we�>]mοqy1__m���#r�.�͖O>���G~�_�:��[��~�������w����z�n�A�������c�!����u�{|ұy휦��s�7����c888������a���8�
�?R�;�IE>F�(�E���`$�/gE_u1.E$�7�dLS�)e.JP����װ6�C.+�6�kS
q$`kPZ���_��NSb7y	�>��zр�I2���'O>���Ã%��"��K<���#���c�ݎ���� J�yֻ���J"�����iȳ�!Jd�l�ϒ�rQlv�XU�/*��6�!�(��Sn�v���oB��3�����QV�jFQ$��#��A�+m͚t]c��a��u��imC�4dE��{��]��A^���Y{6��*q�G*�TO]�~�_�x�u��&�� �o�}�:1�����}u���LE{�A�����{1��!D%(X�1�r�9�����;	���ϟ��:!���z�}��^r#��0�^��NM�ӛ��m[��i��w�����GwX,c����fKV�D�]s�WWk�THB��qآ����A��^�Q5Zkk���ͮ �!Q�Zc%`�F#.�P�J�(i�S�F�� �ص�c0BT�h�E�ɜD��x�,��Q5	8%WL�Iu&����h��|L� �C�EoQE���C�ƣbS����'jp��bTo���Mu&����D5Q�(*&`Ԩ���^�DT����A%�:qV%D4L�����de~EP�ZŪQk�$�K^[P0Q��D�"����Z�}�pyV�l�n�?���ؼ��mk/W]4��ZSΗ/c>mB7��;5���ms�`S>}��r�f��ɬ)K[:g�u}L��ϖ������<���'���<����������~���<�麎��'�>�����z���:���uz��N�x����nJo��m�ޘ��}����X,������v��7:H{�Q�+�-�_�xfՒ�,8>>����fC�J拜��M��(g乣���,+0&�cL�Ve(�W�}$���e��-ƪ����[���q�y�˗�	[;�\��'H��p�wbBHZR���4u��O��η��-֤��(�4�6�����Ǯ�����$�@S�l�[ !�yVpxxؿޓg���<{���nGY���'�P䡿�~AE�1-L�˷�o߯!�r��}�/ƈW?��%)�Sf�;ܻw��|�^I{y�Q��a�|��{]��g4�ѣ1`p�����C�1�Vk�.׈���)���>�W��x���_�o�&"��篻��M��N���J����zA���j̐�����$g/�ɆÚ��ڶc)ˊ�G����|�;����=�����m9??�B��m^s��Nݾ�K����hc��Q�%�Yjƺ^�YoJ\Vp��{#��g�~���Ϲ�����紭��k|�gs�>�2#sE��U��,�X۱\΂�U\�bи���^Y�M����T7�1DDB�k'-5�0FZ�N{�R�bD��a��B�@�E�5�5�1#�%CU����Pi���AU� q�gD�H�C0�#ј$ *�l>����(��b�H!ΡN�LP�1�^@}J��֤�a4J��	"*B��Q�`� N�1"bzb���+`D,j��DL�1F��g8��N,N}aqI�P%KM݂�(Ɗ:�PE��'bTd���fWKS7��U��Qe���(��b��˳�6��6N�%&����]G��p���s�x������ӟ}2����Kg������~���{�71��gO������}�v�e�M�^�I����h�D�b5L~��Z�q��d������ hŵlF{�s粛|���A����������ײ�J����s��E��Lf��UE�%�n $j`�p0���x$�dO�T4�&6jJ���p�$��b���.����ͽ�t��`�}�7^4� �ɬ\���⶧�ͷ��ַn0M��@)�T->b��������.ZB�hm�T��+}�) A��(���ֈ�dD1ZU
4Zg,�e,��-m;�,�<xt��>��O�;Z�9��mFw~�2�G�a�m��Dƌ�(�x\���Ÿu�![Qr�y�eͣ����{�wSd1J�6��~���8����+{W�&��O�N��2V꬧!(|!����>x:��u��ǆ�A�0�%� xK�v�g̦�NC0jz!P"�$G*�	��{0���+��'�8<�zL�^ 2�E��2�H���4�?�'�'p�B�X,z��k�������Z��{~�q/<���v@��٘[�������+/�ҍk�l�@5�'�Gg.���m�6ı�8E"=?�u%��r���w�]i��<�gP�Q|����G�q����Ѡ�!u��>����k����1� ��D+��4@�_�&�"w&�m[;em3v��V���^�_B�6�(�\���>�Wo��V�g���Yk��+Wx�߿_ ܾ}[������Z��U�:(YԕX�ЎGE8���s�oo/���$(��tz �U5Q(
?j�6.di��ɲ�g��"`!4!�U"���ZP�NL�MJ��B�.Z' M�S*(+$�SBy��RBz/�tN� B�
1�/�`��2�XQ���B�P�F���gI0��R���)8�C0ʃBH!\�W�hB�Z��,=ai�.�M����BdƁ�o}pn[y�-�HJ���/��?F΅�y��;����_�B(u�>n��_�u��ڰ�f����2�����)^=?<���ի�x���������ʫׯ�����{�QU����5��M��Y,�H\�|�B�8�Z5U���J�I&� ��K���F�ןdu�P;-)D�o����J�_�.��9�~�u^}� �و�i��ڢ�sF����Ƶ����m��^"�    IDAT� *�B$8�d�s1��\ܬk��1�B�ՆJ�h]P/�@�#���ݽFg����c)�M�W��HV7"�
8p�&GQd���5��ªRQ5��%�t����X�4zW�Z+�Zi,	�zpF)�(��Ҷ�Q&��<�E{~&�1L�'N��1O�6@w���Ma���ה�EN%B�vL!X�*^�Qn��,�~�C}��(F�gG�h�����
�c��,/O'�����i�,�9���g)W��{��	����OJy������Y���_�����$?X�V�����X����]<FE�	R��d��ǝW�ɛ��;ܼv����іs�Y�q�ڵ�/n��|�����K�,˲��:ڄ��f\�������S/k���9|t�|�$7��tʍ�n�IE��`c�U��ٔ�h«�ޡm]�&����> Bt�t1>��/*����k�e+�:w���xY��g�TgR7�1b�_+���?�hƍ�r����]k�r~|,D��HQ��9���^-��΋�B�\V2m��cW�4���u�T"����)��-N1*8畲2H��W6x)�t��ޏ��FFI�*��J
�#��ҝ�,BK��I�U7¤V��A��R���U\�Q¨�DV�m��C��؂���5%����F{-D� ����+�Xu�C���<���uP�U��B@�&_��̜��if'�X��ű��+j�r��F�Vu�װƸ�mE���kN�3�PB0��6-c����@cãr��>��A�X,�G#����{�'2����2�̨�^��7�1�����?�?�z��M������X�i������,�������'Ҷm ̲��֯G9��'��l�N�?�#ȡد�'R1*��)�.�g�c4s����]��|>g<�!��F�1�;�ؖ���oq��mv�v{Ep�c�"���f��%8h��
�k-���UJe��q!2B"���{WnrkQ������}C��U���K��1[�X����ȁ�9�q�t�WcGJ	JS�%mk�.���A�<� (�̠���-��($BE��YI��
���Oi�$��e�/�VI�j��l^�x\��ƛ�� b͐�Q;�6���5�[�R��_i%vV�(YAH�X���ɶ!+[[[�y��������5��3�v<YW f�f�R�8E!E�۶e>��|ޯ-Ҝ�m��o�6�Vr�خSB��I���u�D��	�0���d��yԾl,m3����5����������F�&h�|���	����h�����b:����#|�}���)�{�"�3E1��O�� �m9:=c2��d@*���q1fk:cgo��x���uՀִHB�≕�A(���U�B��Y��A��Ω��_����:�3�te�e5,��$xӜ��4AklfDH)d�/��Zj���Ef����J���@��"ӍkE�&���a<��E��)R/3��v��j��Y�V���@.sh��Ω��ZZ�h\���-弆�	x��m0~�۶�ң��^kC�
�@�(*x�ڊ�P�IW*�t-���!����I�*���RZ��.SN���{�H���VZ�s�\ȫ��:hmCM.�R�;���0˰�b������ ȂZ[8�E봒N�����a��c�\:)�h�H��U���L_׳Ҷ���I���K��;�^{|�Xܽ{��J��G?�Q>�N3�n�\���rY���ٱ?��l�_�1j*W��_��)u����X.z~C�XQ�2M�E;;;��k^~�����<��h��4��HD��r	��y=O^��}�(Ek��ҥQ�aX#�h�h4ekk�K	[��QV�%�Ķ2EV d�m%M6�s,DId~;�]k,��Ź��ֱ-�{6u���"���qaPz���
�٬O5A_�f��ջ�HY��6�d:�!�+c:�,��ei0&��Ľ���n)�U��K��B�|�]4Yu��-&K�K�Sb	���*�?3�S��9pP�L�	����Ǉs#�>���n��,��0�8�r���n�x����Ŀ�d�w�L�� e���-n߾�1�b�c�X�����x�J� �{�(@/d)힎x���_Ş���W���"�08M�(놲�T����P�e���y�[,��|�f��b�7��f$=�yyv���H)���fgg�=�1>�ivv�z��ml��-�A�0�c<˘Lf��cw���-������z�eEU5̗͠i���ŕ���|o�ʃb�5���ն�vP�� ��(U���i�?��?�������cl�?��?6;wv�ݻ��ܽ{W�+�<�n������ �O���uM.��\	������t��6���ݻ]�6'�����׹�=���x�Aw�#���Wu��c����R�E&��t\�Z��w�����?.r9j��s����3ᔒ8ȥ�Rz�XN�B��.ŸiJi�N6۪�B�|ڢʕ��m_��p�p2/r�Î��K9�b\
�j4
EY�J� ��U= ��)�쁗R�u�hfM>�TB7e��,ggJim�k������'����ޘ�F����\iSN5��,F�O����������m;���G//���GcJ�+H�ܽ{W�����d0�a���r^~����'ׯ�����>0����-�,ʒ�|�U���M�s�jٮyI)
�@댋�9R(��":aܺ�{04䞥��1�:���0z5|]zm���E%���W1���Sc)�u��L%�Uu��/*&�	{{{��N�\�}/Ҷ-{y��,;���`�i���S��PJvi�mO;;�loo��k�`kg�E9G����ׯ_痿��ZK����o������X���mۧL��y��F�NJ�X�1������$:�$���R��D>����,K�g�ϳL�#B�8_��5e:����`��6F�mF��W=؊Q�؆-I!%�d=�������4ϴ����*Z����I��4Q�l8��s��z�F1.2Dp|���<|������_�¨JȾ��t�s�\L��0�IU-���f:�0�a>?gR�}1E����%���B�P&R���ӚϺ~�⡽��l����阓cz�t�P�uEX�������G9]������ �4���.:��PUι^�nx^J���";U��c�ұ��k0�B)�K����4���E�W%R����svr�������7پ��:fY�F�ؼ��>����`r4�a�����O�1,�U_����˪{�h\�ل��bL�:>��I�����ߋ� BD�����j:۲U]����Z�N-����]�����O�n�S�4h{�O��O�B�w���@�v/ ��Y�ON3�d��u����������~��B�&=��m��+���������w�>����+ ~�_��O�I,����],�)�O~�Ez�}��������L:�&*��O��Z�{>�������&��𘦶\,TU��m�;⻖Q�$6�o��|�����kO�mگ�n����Sۜ��	C��&l�� V��H�nBNN����ϱ6�����9:�(��l���6�ٌ�h��2�R,�K�m�P�5��ؑAJ�Σ��ry�w-R�.*�N"�lo]�ڵk(ex3�,�"���׫v������o$��1%�V��R��r�����Bj�#:N��zK]5ض霅�P;nd�g�e<)�(���K׹ru�,����d���y�8���
NRt,�x��k��;<ݵ�a��%i�]8R����cGGG�����7��|��(-E?߅ E�dq.���>(|�B���_�E>��
]�Pֹ��]�>ϲ�R����v��5�N��Y����&��4PI�V���Ǯ
�E�s��+_�KW@V)��CXkeY�<���ixmdX�nױ��#�Jc1���,��w6��9#��"���T�1|>}��a�.!��j���%:�v����\\,8?��kAz]��Z�������y�|hl0:ڹ ���8/���_�n�W�~@�W�$!�B����֜R���-F���%�V���1.+���B5ֲ\V]��AL�@�GLR4 .�q�{��;�Х�:5!e�_�S ��FA��{��D�u2�����_l��%1�+�)���,�Ƈ�׋q���R6Q|��M��Fi��He]!����a���=�HK�u�tE�E�G)cd*h���J��/�~��n���x�=ί���s�]��@��$>�F	���qH�2����<x�����s� :��ὥi,�q�2B!�Qp��0N��0��(2ʺ�:��b�G/,� ��qL�&�(��]�$��b�/����>��s`�s!m:m�2?�`~~A]V�F�ј�Hk�u՝k�c�Z�4-��<Q�5˺BJ:0+x�]����Ż�������_w��߄םM������5m��@��C��/�����#|��E)Z���!��Tb6F�2��z:~���] 9 p��o�RA�R��i�
! ���T��s4�C�6ri۶����~s�F��OT����'���:3��BPwm���$�_�٬�gi[��%U�62��U:����J��"�`�Rʠ��� ��r#+����}/g/�͸�A�*쎔z�;ޮ.�j�[��L+#�m+�Hmc����������lş��DN�[�l����I�䋤��퐿�*��b��~���փ�T��-;u]����5��x��A�Q�͒�ىo��ki����L_���x!�"D�hO��-	�&��E����c��l_٢�� VU�_�H<�L���bY ��u�x}%��9QH�-����Z"�Ƈ��A'�#�z�T���-R	��<2�6EⳮsN���{R��E->(�Δn��v��0ґ����&�֚<���۷oRU�pzzJ�ƴ���IN�2nܸ�h4�������DG��� ���N�`�S�C:F����Ն@-X�C���k���4��}l}:�����f�Kkݧ8S����UJQ5yV :�<:F���YA��H�P]z�B�tp��^?��2��>��-���N�B�H-�
�����n.|X�9���t,�
�aT3=��J�h��&�7=��)%]���|�|�<�i�lL\o�~J�a#0M=uE,8�b����� �B�B �]�7��_�	��F�Aߏ~����VB���k�Dx�\��M��=��r_�QMc�VBi���	��������,k�]!GU�4sXq�I�O���G�@�u���@_��z�=/�K��fD#mr)�eQ~"�z�`a�֚z (�x۠��f~qF]��#9wTh�rk�t���"dL��`l�-K�����N��Y����ՂE9�n+���X-�k8���_F�R�\�0W�ù(vj�AI�:���}l�����،<�jg��w9*ʾ��Z�����=v�jI���`��ԇX�m��M;���"I�Em �}#���j���#¡K��o ������tʝ[���%�lo��3�Q#D�f��7n�e�>���������n��R�i^��|���xM�9̗��Cp�����ۜ�B�\nC��#
<��k�ް7y_������ZO�bb�4�d�QD�*��*���يk����f�A/���E��#GXE�D !Bt���*��!F�Et&����ԋ<��t�����Ɇ�z��4�ctUB,KiݢXU�6�W�~Ew��ή�����>:G���7"/�pa�r��Ʌ_�WԞ����?V��Z�L�Z_�PI�}�loX/F���!h��Bʖ�jp6V<�e�b�`�\R՝j�`���gll��GEV�6A��ؐ��;������nO�����i#}����HBFmom��=��~d�8P�Kc����bR�T� c�B�ض�#��n,ZOb@Į�6�M`Q-�M��W�%ی��Q���۟됬�eYWuk�wR+��նu(�P�'ޢ�D�碦_��v�z�.��c�g�/5tH6������ �����(� 6\�s���d?�g����lm��ٙ"$�&S�� XJ�u[��LF�Q��� o-Ai:l�G�DQ��:ܠsI�δQ��˾�%�>R�v��xX���@k�^d��=+z��J`��[�	!8??,0��%�p;	��<��{�W^����N�^k&�(g"%k�����A���`�\������w���i�}���k���/t�͡�v��m*lS�J��º��u�2'{�;j��s3���M��a�_j����>��|�9�v�AV?��c��N1B���]1�s�{'D����E&�pA��?Uw��w����ϔ���i���K/�d\��ڦ�i�ۡ�oi����1�MdB(B`�����CU�,�Kʲ�i�ޫ��L<y<��|��RR$.ti�4!C���K��~ÈFz���5ӂ7��t7��K3D�	�u�5Z!B����M�S��6ѳ�]�^A���m� d�<�9��6t���bU�`p�%�g(=[Z���]����^>�^k����09L������%�R ��?�w��9�[���g��l�z���k+����Jhvw�0�ls~�����z�!���b��m�@a�jx�C`ӟS�u�����'�c�|So�����
@�llϩ���{7�1���w��Z�CL��h����G�M���	e��;��u�����Zں�>?g2ʘ��\\��qqq�����8��iKU̻��ܹs��7o2�N{�����J�����G�qxx�GĆ��i6��Y�q��-^�u���h۶�qxx�9L�OgyT�t!T�'&�-��*�����ʕ+loψ}������dru�9��!��߿߯ǩ:XJ�Gע|�YbZ4�@�,MS�45F\���՘N���4�W�<U�.պN�H�~e�������}�C)���	K��&�)rYe�g7�v��<���  ����',�K)�T!��)������e���!{&����Ea��B�.��M����ŭ��!d.�Y�ڶM�P5�Wl�4\\\pvv�"��{z<���a�b�e�͎+/h)�>L�$]�M�aU`\��?p��TBpx�ҴqS2]�!.Tݿ������RH���xD�F����Wd��Z���ֶ����9εa�F��Ǐ���REj:ס7/���d����{\��G9��]�"���=����X�� ���Ǳ�(&�|�\�r�G���s||�Ėa�'�6��#+_�ml�������z����*��}��� EH2u�I��X�y��}�1����y5M#[ư\�,�
�$����(u^r�:����=><�(88�k�"�D���d���-i����|�����7�d{{���^$�/�ܿ�w�}�>����}���Z���lM�N������?����e���>�������=g3����&r�V�h�x<�ڵkloﲻ{��l�U[�uG*��6!B�Fݤ��L�yN�\a�!�/Yn4-�֦}�Ź����=�6#�J���x=7��%o���=���E�}��5]���22����{��%�u��g�Dk[��D�TȂ�)�wNxB�k�����X��'?�r{H_ۯ͞�*���ۚ��Bη��(������C�~{g�:[�mB�z�y�E����t���#����JM��Y�e����u֥Z��fк���NF�U�}3B2�`]����)�#P*0�Bȼ����2��N@+R{-O� H�!r�\@���Œ�j�"�;�"�׫���=��#�ж+1X����N��B#��X�AZpb��;hs��\ń	�Y�-1£q=A^"A��;!��b��"����Ł�ӿ��T�W@ ױSIE�5����,>�m^�l^st���6�RKPc��tdN2��A��l���.g瞳������;�!M�rxx�T�(�4
)A����Z�l�2�Rh$���8�dΣZK)v���b
�G��GT�#\3c>o�׊2LX�#=N7�� L�h�/tu���ʣĂ�{���������	/����#>�茪�bUMۖ]1��i���S�F���A�!	,|p�#>��N��ͮI�1ʵ0Q�i�αl�����Z�Lf����    IDAT�r=XQ�l�����a[a/.x��}�|��5|��G=�mK\��"$�o�^�oα����(�>�����!o����(]����t�W9e�
��h��#�2
�y�o3����_��w�-����_B�d�s�&к@���AP7'y6��+���0�����{�G���y��QL����¤�c����O��ã{d��)Y��i�[��	�;Zo1�m|0\�im9)+�|IiA�]\�chj�4[ܣ�-�y�#���-M�E�����O??���9���x K���K�+32���~YU���HtW���Q���Zl� dF��ف�ʠZZ	��u�[]�%��p_J�Q�d2YE���W��L�3�`�$؊Q����Z���m��]�gu�PE+����'~���5��v���O~�g���F���e�������m4��mS�m���qV�\ۚ�r1�"!hk�H�ZY������t��S}2��i���<~��'m:�M��I\�gِ?L$sί���+%k �@7��--"��I��e�����ަ���8Kq\���pzz���9��"�r�_�o�w�R�[[[L&ڶ���,VC�RA�-u]�eLM��]pzz
�����t� �F�u9�1)
����0jZ���c�2X�%��R�bDEM[u�4��9??���ggg�(t@
�)�e>,UU�ӟ����^��������^A$���\�� �Eɣ�c�j%>�9�6��Y��_�6]���1J����*I)�N�YN]�#���>���G9���|�"�D�n[�f������(i�9�~x�G�c�Y$��UJ!t�����9;;�W_����=�����ƭ[�\����"�
�����ߡiJ��k���=���lW*�aEt����޵\�ٍ�����&�=�;WؙL�'/���n8<<���}���p���b�������et��O�~}�1��dC�4����&��2��g�&�h���v~}�4������<?�=��lD�N!��cc@�	)����Tq�w�{�m[?Q�|��ھR�D��o��y�P���������>����y�|欕)%�8��2��I�uC�Y�n��?ib=m�]69�mN���0��<�g|��6�7\��0!�m�I�V����1i��X�f�{��sH��z�*����P'��x�ˈ$!�?����}�������I�t�fdQ�,�cggg�����>GG'�Ŝb�Q6U�Df��޺��JF��8M�s0�C+�4�}C�<��P�������9:9������R��ô/ҵ�ƴ�!����Q/K�}��-B���� ��K�p�tk2��o}�;�nvU����s��d{{�k׮E���'g�<x���t!�����4K �����~CmMc�n�m�_ҡ,�`6�f<���t8�y�`������cL�۶�J1.F\ݺ��{�Ř��өb�&�)gg�|Y#��
.��he@)������|�{�����s��U�Q1c
�� I11�~U#��(m����()P�T� ��,�|��'����f3�2(�3ݽwx�o�Z��Ԓ�(�m�g�~�/~��}�q}.ж5�iim���E	I��]˦S�i��� ��5�`����mF�6�线4X9KB���)�����Cǉ}���?�������f1x!;�2!@�y��|�h۶m�.���eO���y�PJ��u���������U�^�u%�i���n�z���3�c�/��I���?)�&�����z�M�˵�ަ'�����=�t�B�����$�O�(wQu'j��V��<�#}�i�=�}�-��C���^�@���0��w����"�z�m�`%��$�?����i��T�����:23��.��f�j���"��j�Nx���6�4��9�E.��0�B�0�I-τ�Zj�.]�,U=_E<dlٖ��>D����j��E9?���u���3<x�Ғ�r���)�����C�b��7�z�:��'a�)�Z+��7\��4�֪`���,�x��Ke�{�TdZ�n������W��/x��88���&G�8}kɌbR����~HӾʕ+c�f��x�W��u��ѽO8�#@�LNn��X/OGl�v���m^z�6W�^�+�r���m\g�D
M�%���w�޴-6x~��_�����xo�ʐ	�ف�����T�9!������l^���j�NNN��_�����?e����;/R,�����p�F�n�t��)�r�7#zC����a�m���y���ק��/�qY�am����sx���ވ.
!�A�����|�*���w��]N�|m_�.}?��G�,)G�r��<7�}k�"ǅ<X[�U�ؾ��m���n5���+B?	����`6'³#}���gġm
i�k�T���&hn�����3-v�h�"�i��7�҂��qn7���'�����)�KH�ٞL���6̛�
��TfB�{���I�%�E��/��<�p��������)Zo���KKY��pq���I<�'�g�<Rx$�Jx�z�s-UY"���Ѻ�T���G����nh��E=%#J�����cQ�?:��.b��!k���2s�_֑̿����������Q*� ]��1�!p��M�wv����{N��D]6�i�g��xo���Z�@��-e���K-�����Dmȶn�R�<��9?��ˇ�>�v���@l��#׆"74����|�U��aRL1f��Uv��"��X+^�4��A*�����[������Ɉl�̜����G�89����n��׸ze�"����o��Q���S>�A�Hap>�Enȵ��Nb�*99:`<���������-���}�O�	�Qt�5�9��E=���#x�Qp�Y%����˂CG/9C'p3�;�5x�|��eA�V�Li�Rq�w\�ZO�򑻙���� �y�k2!��!��}�i/..��/���E��I�>U���fu!��.>��=��R8�2k]�"y�A�tΒw�Ti,�G�6A�����'�U/� ���'�Uz���n�06m<��u6\L�����M��t��ӳi�s��9���@��@����0��#i�)J�e#cG�t�����soC�{��(��>V޸q�o������IPU�Vv������#���� �7�.(��3��F
��l@k�eTu��);�>�(f��k�LJ2[
��)�@����)���T��ց�vR���˷��-B���lmm1G�7�N�������D�.wP�|2f�6l��MkЗݒ�L]V�4�b�����hIP� =���P�������2����Lg�Qڠ�F�����G\�q�7��m�����;c���9����+�������!3���)o~�[ 3�v�dň�_�;�1ϸ��<��n�Jl"���r*DY�kj+�]KSW�u	�#e�ZVZ�L�ZK�mc�8HB����ȠR���:��63J	lmfAV�T�&ْ��Pӵi�����w��a���;��瓢|�<BH����(*� ���]q` ��T��/���9B_�W�}o��vѶ���#��*����Rd��s�;'���d˪�5��R Ն��:�2�7�'EF�'z��ϻ�Ƕy<���_Ԟ�"H^�Uc��_������{~<GÁ7�?6��.Z����>k[��b�m�l'�b[��}J$�U7����k�x2����h���Oxh[�/N��BjW��˯F}�N,7����CzK[/pv̸�L'�MC�ZH�-}A��(+ٽ}qԧd�

.~^��l_A/�,D'D��\�޴iꔢ+�G��ҭ[\�~�����6lmm��=������C>��s>��3���d��R�9PisY�����:g�!1�&�b�O?/|_к�-�Z��#��<S4�pX�"���.�������}˻��:Y�ڠ��z�:CX����;�����?�6W�_�0����'���|��y����G|��4U���n��c<�p���L�S��#ڟ����#��drL$�E���6Ff�%3D'��%���K�H|yD�*�S�&�s�ZE����/��G�9��^�o0��Q�˲O_��n�����@��>����JC:A��د7�!RI%ʵNz��!���l�/tB_�W�}Y�����N��`~h��V��Xj�#B|P���\\�b������ڶ�ҽr����j��\О����_�'�Ӣ|O����MI�.W `��6mC�Q1�.=��=�mr�.��<��y�n�U%o�e���]B`�D��޵έ]��jrP�g�EH0&c:����KU׼���\0�M�_q��+\�v���=��������R�������'L��'��e�s��N�?BG1��zįA�nu\2F���ƬG�AU!�`�V��D�SO��0�DG��U�����:�m�N�r||�2v����ˊ�j(�&�d�b>_P�j��������zd��q����i�T��� |C���%A*>�
���e	�cr���	�~~���9�o]#�69٨��k�|L�O�fʝW��|����=����:��䀏?|�w��w��3*&h3bY9��'ܫlӐ��ֈQ1�(
2}��ͽ�?���1AI��8��5��:���#eҿ��a��a{�T��[,bˌ�}�m)�k׶4my���;�w��	\]f鵛���Vlϲ��!)36�	�9�.=�'�כ�/t��Y�"���
�۶�vޣ��(��J[�6~���EQ!�L��[���·+�h!����9+ j=���Ӯ����p�X�QC	V��4d����~�EC`�xp J�~�%��m��S
�o�tC�LmZz,�K�RvZ������g%��������A|�^j�7Y#D�3��z~IU-㢗�]�2��\�w��	��A�:��$���J�`mۢ�^S�-��@�����W=#��燭�ڶ[ػ��m�RQ��...PJQ��r�7t�x.�%�~�m	��V��ӽI"�1��y�.p�����Y���"j��lw�t�ŽO>�O>A�N�΅���P=??G�t:f�5鮅Z��q�	��xa"N��x��8,�HU�����Ti�e87攎�R3M��ܼy�s��atN���%�~�9�Ucx��7�&����,%�ɬ�F�e�d4��D�X��|K�$�eS�yF��(�춉�i��j�B0Oh��O�E�G�G�@�#�K���$�P�5����!(�b��3&�)��S׎�7n�ƛ�ag�!X�Q�x�d��?x��G��#S#�o�1�L�8?��'q��o�v�I�G 0o*�]��믿�{}���D�ڶ��]d`-!8��h�=�}w���"G"��e�
i����MS�ܬҠ1z[\>+/i���Ul��/��D�e����f�Wi]��Eֆ�9Yz<��9}�����&�iHQH�6�M)�Z��dY���jq���G!��#2���Z�P���t~t�:�����dk�oZ�Fk-�.r���͵{�ry� ʇ@�C|6+�`5���L�o剈u�1�w����O�e��
�o�f�ox�c�*웑���!��;'�I�����t���]��\��7a�]�a�Lj����5Z�l=��&�����w5nW�b� �Ĳc����)3��lo���͛�<ċ�h�sx���~�s�O�;����3�A�B�9 ���)걊\���}!���9o�c�2�qcy���|�7n��g��͛�w���	�n޼ɭ[/���e�zf��8L�{�c�E�%s��n1Ҵrpc$�XI- \��'b�G�G��cB
�A�h�L��B�T��#
d"V�m�x��u�'̗%J��b���t̍�7�y���%! e�ֵ?!�'bJ�!E�:e�+� +P4�Ц5<i�^���q6�6���(CN�e���|2��S��c��K��9��|:.�c$4�5�S}p��,)�����5���F�CX�Z�f&��[o�~�<������������n<��&�����Jd�û�!a�����ZOUU}��չ��5�N�%���$�#V�ڢ�eY/߰\./%s@�	�6%W��>zR�q�zuB���wi߫W���&ppp�sm����s�{�1�F�~[�oӫ^'���6E)ʴj����m܊���;�N��൑��X�9Ej�dy���yUrpp@Ӷ��#~�o�u,l0
k�Rj�2��������+��L&���7�:����<v�H}WS�7i"<{ %෪��w�v/�T�l�M���C...��f\�~���6U���_���l6coo����_�����-�n_����'8��m���XW�����.8l��@J���:"j�I�q��k �Z#�J�,� �֝p�H�Q2�輏�`	�fgg��~�����1_�� i��m$�h��h�k׮��K�����-��(�8օҤH1D �틄�,�c  �߀��W�MD���k_�Ս��_��۳��X~���\]�gR6�POs�7���a��y�e��!(�cr
c���Z��8F��b�M�I!*˼Tm^
{��6��N�Aߵk�dQUҵm!
�mx	P�����&?�%W���ٝ�{>FD�SD&3IV�J]��%Ah@���� �hh)�J�6h!h���$�����Ph4��"����$YIfdL>��fv��{���##��,�ٴ����xG��|�;�q V�ng!�Ty:���V�N�q��"lӃW7f��.rڽ��`a�:)���ӿE�J�Q��?W�����
�?L*C��:\-����͛7{q�rqqA]����_���~���?�n�d|�M�}
���c�o=S7�j���-���s
�v'�!��u�,�8::��F���E�ц���s�3���py��~�9M�k�&�US�i������_��_SE^Q�K��of,����k ���/q*~0��������y��	�����w�]�x�.W��]Ĺ���d�ܦ4UU�u}��1-�َ����c��U��� @�F�"%�^���_�d>M�l��1Ɓz���FR@5����X�'-x�iRpt|���w��Z�� � %vr�|FQ8#����Vc7�`�Ez��S���i=�Ȁ�+=�A�b�%����1FT�L�!����^sJ@<��!�X�D�jp>���N?g��+�p�Z6|��w?wwN���S�]��]���e�����bY�V�1"��k!�x�
���8F���Gu���_��?*l��������hT��2�!�6u��M3�<��@�Ո=���y㺛lhV=M+�P�e�NlW��:-�ˀ��Ŵ@�Ĥ��tLA�"��f���i�X��B_��w۟籧��1�ئ�v [y��Z���)��P�+�v��x!�~�>7};�=���+l���4-��~��|�;X���ϸl\f(\IY��tng�o��&�~�9��4MC���0����t����4�����U����.1�7`��϶��}�����l�S9�T���Y��uC���s~�ӟ1+g�G��b�prr£G���@2f��WdW�]�}zs*ȏ=K6ݗ�N��-�q��&*��v+���5�w�}�b�%���fB*�Qk32���ɞ�e��4g��rA] $�؂���Ѕҹ��_�X�f�%�!�%�;��3 *1.Ukƹ�uC��|����8�y/��@��n ��j���_���]��)�����Q`���l6)/�q[@�2�AMU��i,��u�@|�_{#?~'���=�������;+�2^\�1bct!҃�8.�S[��؀i��*����ލ�v���D�RNۮ C��f��`L?{��/�������_��]a� (�����o�Y,���^�S5d�
��θ.��c��
���������<Ϲ�����t|�(�Y��X@x'��ٕ>�4���3��!}2�]�e��ߧ���}��o����_���ڶe�ڑqN�m
��4?��OY,<=9�k#m�	!�����;�|�q�M���/*�~`ڧL���~:ޏ��r��g    IDAT���x��	�}����T����_>�����9�����o�W�B�qxlH��뒗�`uc�h���'
�k\@�C	
��z���s�L2ж>z�lBǦ��1DI�W1�z�e0)�,��jr6lښB3�v�A�jE���_Ij?*x]NZ���a;g��w�Ok?����1����Ϝ��o��F4��]�igN��]V�y�^���]���_zc�G"PU{�<������Vk��?��˲*���
	�*�JQ	Ƙ׸n��������,�[�.����m+H$�Du�*���T�0�`�Y@w�5��l\���2r�:�D�����rd�՝�q��M�_|���a�ڶM��5�H���m0Nd�
Y�.h�0j_�~�/�x���]�ї���������_'��y���i��, �l^H�W^6~�v�@������[�U��{�ɓ'H/#���O��|����٬��2���&����#BE��%������O?;�Ó�G���/.iZ߳'��נI�f�+�(ڂ����\0�&'��j���10��|�Ij���P�%1��"'ONyzr�r���|NPX�j��dY*�I��  s��$ ����!JL���d�w�o�AVfUNV䈳h��+}��՟!���OQ��,[�B�e�QSg��1�N���^9?_�\%V��cFr��i��3�.3�J��,Q�.D2 uߵ��M@�v-�}fZ@,�f�,I�����B ���#2^������Cfh7�m?�i��1ﶰ���u߱�ױ�S"c�=�}q�����o�믿����׿�m�"BQ��Z�AИGW��ߏ�j��裏����Z��bv�W�q���B����a��M|�Dc u�<v�������U�o�u���N-[�y����:�su[_��&�aBiۖ���T�>{��������l�����|���ݞ���}�睛��Ƙd��4�8���W�s؍��k���|>�/�O�>e6��;w��?�c*�|��gt�S�9���*�M������/	�_ �Յ�m[...x�p���%u�����5�>�]�]������:��-QO[��.`]�Q��(�h�~��d������A��k3ʪ��o���]@>0.۟�4���k�P�=HR�e
�F�����d����([����&�Xr�&�&���_���<x���kpE�s9�1-U^2�U�U���1�_;bo/��9�+0���gR������Y��X��m[�������h�2}�=����̐)��i����o����>,^����#9U�c�Z��\�8<���o����w����m�K�~���\o�!�<�؈1?}�C���;8�����r���zï����j_W���<c�*�͆.���p�f��&���!G�`����7H�%K�A׶�8�������G�tL7XY�}9}���%ٗ8���� ��{x]Zvxn�����kw+la��4(��g��:i�h:Ď;�����1��Q��#6st"C�E��!�}�%���������L�b�f[��������%fk��4eq԰�g��ĎE��9��=!�(��?�I{�؝�v�� ����m[�>}:�F�g�`�1�F�:1�"�` ���H9[`l�f��X3�-�B��d�h�1l0����,^-j0J�5��ir��oY>=�,�4���~����}�EG�C����f�SBlh|�j�A�/����J&�e�/@
px�k��ڂ<? R�v�ɖ/u��7�^b\A�AME�w����,Ѯ�v-�2��A������f��g���~9ccN��9�+�l�D����%ưI��,�ܤ�0�1�brCk4Z�1ڦ���nr����bFפ GE��s�_���:�񂱞M��5�r���KU?@��<_|�>o�(6�>�l@�
��p��&Ȝ�7XSp�v�0�Ő�!(��D����φr�2+�v	�ѵ3j_�X��7��	��%F#y�g�>������'?ͪn�\�
(Lj�+�d�x�6o�s��|�����#��32W��!M$�>uGQO�"��
��hP��2a�˜�)MS��[�IZ���s8OC�Q�C�?C�>O�r�}%�
�:�d�b���IZ���d��to�|��>���|�,�z��<�ɭ#DM�(>��A�1�4M�E}��za�WEE��mOz}�z�K�fgq6I��2���uڶ�j����߼���|�?�����>{�����&s�����ͦ�+3��6t"񍯾z?~W�8la/�ce�|�FD�#�aA"���X�׉i�!�Eۚ��x핅R�EU�,3��JQ���Ij���O���اo����=�}�ݸñxј��#�m��دM#�ADݶ�4����G������u����E�/ұL����x�v�M ܾ6U�]}�0���W\_	=��k��9����Y�H}?SjS�퀚�ӅK��=� 2���y*�@���^�7��5j_��} 40��u��Q��,P���oB���P1� E�%��j�P٫22"��s|S��Yb�B�A'��5=���[Ӹ�=S5���c! A12�=���� b88ا����4vm��eܸ�*��������=��v�%ӂ��|�D�F%�U�K�K�["�.Y�Q��])Y8Ǭ,	]�z��,*Y��S�k�CQ� X�vM�58gp���}J ����M[?����b��n��;�?�=��&Fx������֍~��ۥ��eb�h�I��]��ד6\7�O������A�\S���\2 �ymZ�7�[_5�:����[���g5b1��ɡ9���Q�����7o�^{�����tE��˽�m�\_,�e6_/�U3�F��S#�]��߷}��oZ�����<�YQ�m��ں ����""��L�5��z��TkS�5�B�P�Fa6�spp���UUa����d��7��h�	;U��1[�U��&�]��U���tz��ƴ���s�D �l���=�Z�(��dw{���դI|��@z`���Ƌ�PI�{췟5�tL�8��ɳ�Ƨ��Ŝyf!�t�s�ӄ��D��	��:���*1�����CKQmϑ�#���Lc� &��o��Mz%VU�7c�����7߸����g�Y-ϒ�N,m���\�+'/��DC�$��{8�����oq��c��%��s�^�xM���.Ϙ-�S��$��yU�g�^�k�T���&}ڬ�ǿ��0�z}�����,�)���r���������#n�~��܁n�я��:��A�a�����7��Fb��	��J& ���4�b��%�EA����A4���;�dF��5��5upq�����`��uZ��"���Dv��a]�������$���+�͒��CL0Wҟ��cj��1q	p:�(�kDl���+��WOJ_o>�.��ʀ��D�����(} p��iX�ZxMר�m���AS;df�4n�2�޳W�Q�mӐK�yꮥ(
n�r��w���l��?��}���;˪�m��z��iV����xs1�F,D�R�ks��k�ߏ�⇻w����՘�T"�2WU��E����>-X��U��#"�,���V�#I�s�֭�a��a��i7����{fS�����Xh+��YFj�c�����/N߼<+�U�q�v�9Gx�04�쓼ܶC$qZ����4�t��)=���K���d:��}h%C��D��"}�Z�jV�����7g�<������әQ20eەί�>M�
27Ø��S�Q�d�lm�e	��{�Ǟ�S�ٜW_M�x�&U�&͕P-��!v�1��������'��G��O~��ݴ`,1
"I�Ӽ����v�dICi&�W^{���y��-�3r����ˋ�h&��U���;������<�.s4$�E�6��V$38��&,;H�-;���nY�qx��W����c*m�6V�Cn������َ��3~��_p~v�_o[f/��R����7��3�ԛ�f�D�C�;2��0b2��Q��!Y��� 6ptpȭ��̪��Wl6��I0b��XWR�,c"b<�j�!�b��eP��@Ҧ
C��T�#F�Ce$i+H,_���OÒ��jp�R�͘Aʰ6���6�S���ϧ��H���UZ�an�(����,i����ޭ��}�Âl��]H����9��1�M���s��}�3WV?��j]o]���~�)�g��wc�e�4*1�h�1��3k�ۨwZ��{��_�p�gf�����hL��Sj����^�MӠ>��ʲd�~��>�p6go��|���zk�x��#�:U����,�ެp�1�͈1�^��҃�ݔ\�BׯО��>㺆��k^�<wטy�V�<�����B�X�9�DljJ�2�y,�L}Ù�od�{ʪN#ik"\��DIiЈ����#��y��_9���#�ք����xd� 2�,2�5��%�cR��*���
4Kj[��� F|���[U!z�{�n�<���)~IYVW�EU�����w�Ƿ?�.�=���!?��O؄��ށ1U`�ʣw�1Ơ��YVp||��߾�뷎�Y^����?�A���31���f�7�88�KQkh�5{{{��-`0����O_	���`��㙼6-]<�����Yl����T`209yQ1�/8:�A����K)C1�9NZ[�1�2�~��F�f����g�c��g��,K�WԤ�cR��G�:^{�6��6�2G}@���K��ϓ$A��`�l$�8ź��<#/�5b�S�p�!���8���.
�ce��@�T�g�3�I�D�m�_�}�����W�����9�з̆������p.v37]wu�we?/Z�D�f.B?[I�碑е��,pրFnݼ��w���?;�</b�7���<+.���y>�WD1)�u�*6��uB��j>�z����~��G�_����S�}��_Z�;��9��yL���*2e�B�EA���w>��g%Gܺ�*��=���'�z�`j�P��{2��f��ގ���)=�|[�iD��1q���a��z� �E��)�ڦ@�x�=U%hD4�5�c�!�b^�bi�@���S{~�����Ę������׵!�������H�޸��������|�Wy�W�厧�����SX�3c뼘ͩf�"��e���2�8��r!�����im�y��_��[oP�
�6E�#H�>�׾hj_�GVV��TA<�ރ�ϷI4.�����⌣A>4�`]�S�%CUU,��KU1�3c�;��#J�6	��	�L� ���n6��c@���i6}���N�Pb��,m�+��;`V-�=m�4��u�Czw�L���8���F ���;䭷�Ҭ7|��4�ŇTt���8KQ��y�M���c���w��tmMY��Oy���V!.�J��,��&O����� ���#����QM�Z2l�0���P{�1p�����'�!�[�J[w�.��ldq��	�b	l��u`����|���5���W3�sS��i��U�Q|��/$�ug�hL�O5��O��{����(J�>9����N"q�}���Rڶ+˂�m��*xpV��hEPcqA� z;�����޽{'������~?�^�;==��i��<�L>#��W���1B�v���WF�$Z��#F�,fs||��|k3���X��\��|۷�I��C4U�%����*��]�]�qE,<a��c�^��{��o�
1�?ϓ�~(��7=Cd9���c��4�k��{���zI��&��F}[0��l^���&�9v?{�}���u� m�P�2I2v6��+\��Bf�TH$��9��R���$��,�c��;;�Ȅ�}�I�4-}FDȜŕe�X^\�֎�y2c���׷vm �P7�:��i���^�l6�(g�9#Ĉ5��o$��R��c:�^�8�,-�A���l:V�����-j��.x��"Y��Kתźl�oEl���4]ϔJ�K�~��1X1��IŚQ��|>6Mͦ	�Ͱ�@q��s7�����X���a�v��2��u����6
Yf�Ǽ��?���&�����%�M�k���Y-*���'|p�ۼr��1p��)���'����E��Nט�U��������v~���-��AŌڻ��h���m�R!��AcD#��Ohj75��B8�����j*n�IB�y�Wc���p���|
��ސ�麧����;D綝�ɑ�|�"�?;�Pb�Ȝasy�_���G�7o�8C[��O��������N��������w�<#s.�E�v!h�]�{�������㏟��~��ٟ��E#iܻw� ��?�?�P>��c�������R���q��I>:?��~���� �/��\������E���B��������ƍ�_{�;?ߗ��;NN��ƍ�z��}�}�������_�p��R88�{ĠbrUo��S���~t��òX�s�֫���u���s���G�D�z�O7�u��m�1��c?}nL�M������غ�z��������f��1P_��m��v|���lk����r�Z9]N���q"�5�ױ|��^t�v� ]��aHJ�^��	�5l\�!%�:�b�A7��Z�:v��k[T��4S=D�]���[Oȁ����{{{l6���3�,U��Q
8�]G�帬��H^�1���vKM���c-N����e�R E�M��,O��ITn�>X'���B$e� �Q�|ĊR��]�s�u	$���u��� z�w��	���kD$�����W:�ڵ��*�����t���mi�T�Q!
�W�=�x�=n��:o��O��qvvA�S�y�8�q�͛798z�7}Т|��O���gV���S�������MA�1�	���	D���TE�r2�0*D�
E�p/FM*��I)��Q�@��ԛ1�}��v��'#�&�gX�oȜܘ+ݛ�s�nM��� yW߷�^H
����7�րj�5�]S�b3�t�D�Ռ�����?���5~����������A_#OO��޸s��52�ϥ,�.��m�Vź��Z��e�H�T���_���|��;w�5 GG���%��������Ł�ϗ�$�I��O�	K�b�ң?�|_��������E��sa>`���ê�ͦ{s}e[�u�C��N���θ�+�r��23ޠ�>�O`��6\�����{pq�^�*��9�rpq�7n��­��m<�߿������߿��Yy ���9?7{'{�4M8�}*s���b������st�h���ߗ۷o�p~��G?x�Jl��[o������&ڼțu�:0b�*R�A:�����Z,�mZ.//q6�����.F888���z��7M}��Eu��l6ڶe�Zqzz:������*6�u]�V�Z����}��޴�j��}J��qΡ���r9�С�k Ä��y�f�T]Y�	��-��H9�HfӢ�uE�<��뚬�Fp0�G�3��E�,�g�u'�9��ֺ��m8n��� ��W`�"��U_}n�<�����()=��`�\ARu�b�@5�����:t��ia>�,g:�{M�]��D�#��o��2U�>@0`�M�L�R��:B�8���쒦IV2���N���l65y^��-�GĘ����C��7�u�|qH�>���:)��e�]�ڌ��QC@0.��L��օ@<1z��h�Z�XU%�YEa��B�ئgx�9��kW�hH�P�u-.�8#lV+�͚�zMD�7-�(P��@��*��Wdԝ��k��"v�h#1P��a}�V���xQ`T0y�KV-�z�Ū�����8���V
VB�$��ggm����5?����w���y��1mW��6MG״�9��l�ӧ?��<<�es�M�K�2����g3���8�.�H[7\�^p��w�N����999MծU�5>t=A�g5h)�=ڮ��"G������l�������Ӳ,�l6����u|���p��S��=��&۪]�����r�;��$]ښ�O��a=����2}l�Z�����m6���[�4��:}��|�T�b�mNOOx��o��W<�����=��������w�ʃ!{!���,�fM�̾��o�o�w'�?^���*Y�AbUZT���ܓN    IDATET�?tm�'���J�� Wu�ie�Xi��^D��5�w$�pb���ցD�x%8a>3�M��=Ʊ11ΈTs77̚�n�K�����;(Ķ��B̬�U~�l����n�cC�z1!�,����!�.j� ��<-��b\�}p�����y�ESA	������tvS�l�A��x�ez�7U�����N���6yfo��u�J��d�w�j���;�w�6y�m[h�7Z���E��f�eM����ʽPU��.+�B���W�;_����(��Vwſ���한��o�f�ݸ1��ixp||���������Kc��l6ݽ{�����NOO�\�5�+13Q�1b��ī��mT�n�,�x뭷p65Ä�&��׫x���(Hk�dbY�e��͆�O�r~~>�����:�Ŕ����S���޾)��g��1�u%�,��z��qS�X���)к�=F�>Ҵ-M���-Ӥ�k֯{q����n�~��b۔]�!b�	�5��8`zoH�5�0<����C_tS����`$1Y��a��5�-�RW��z�.��ζ�=�3�R��:V o{٦s�ި��*[L1DL��-$�kX�R�%M����#���p����� w۴ب��1U��3�;���,�łX���5��c��H:&�Ӵ.�)�j�6������pǤ�����g��M��)��W&y���i �@k��9���J�z�L-��J�U1�*M}��ܣk=?��g����|��R��s.�k���e�;ڮN�[��'�i�@����զtl"�b!�v��3��{�����3N>�9���}���;���Z��4�II�Ľ��>=y�_�Uj3���#.�c��̥-Cg��Q�˜�N�٩m��Bi�Ϝ�磌g�G'��4S��2�~��0�ͮ��kԍ7&U�Pׁ��u�<1�ܹ���G�����p��W8><B�ao��#O�HF��C����7����ˋ�VL�>е��T�C���\_���FI��Z�T$X�b�zb�eTD�Q%�kC1S�̚��D9��Β�J4)�*JĘ`����FUEĨ Q�	���V���ŒN�Һ�v��-&�L碪��r�ƺ`:�Y/�b�[G�FuAr��G�k�����R�h�4�t��D5��U�#&s���-vf6�"��"��\��3�f%q�\js�l�XjŬ�ܬ��;���K�ɨ8��1뎉�Hې�m^��q��q����v�7Y�B6��n6�ʲ�ks���b����7�g	٧]�uw��]��?�*��]��<W�$�6"#:rwӃ UUq���͹�\�&�ҋr��k����w���ZR����#...Fo��b��dL9�7Ֆ�����5ɼ2�N�=}�5�E�S6lH��_��_:��	�h�f#z�u�l6�Q�͚��s�����A#/��Tӹ�n��z�x ��(1M�:}��@H���\0k2��r��T[1�X�V���چ��X�X�8��t�2c,&�WR�)M�����B�5l�5���z�����'Ӱ��&{
��k��V��#Mo�������.��q����u8vb���4��L�"�u]ӵ5]S#�2G�;p=X	0wm_���
%*u����1X㈴ĘLq�
��i��8����₋�%��IkȺN�M�\"m[�&IF�u��S�r��[��g��k׬�K��a>K=�����Ԡ�>��Y�DB�@$������'_�����OL�5�\h�!lVAl9y���}�)Nj?������4�ҵB��@S�ԜG�rۉ�a�gg�|��߰٬x������O�tWto�����K=�-�؂:�I��ᗟӬ>�C]o�(�!y�7��#��LA�.H���yN����֚�|9�A�<�4ד)�{�� ���Sa���bI�<�ٌ�|��w���W_���^����6o��M����t1����l./8]y$*^��(���-2�yF"^���ω!��~�]����Uc�D��s�XH�D4@��QIii,�2�Ё�9�s�:^��X�V$��#U'`�%s���	䑪�m�UM�լJ��mG��/ۋ�.R��9��2�>7��Ġ��� �b{�U�:���;�մb��"�;�D�v�� �X���"�Y��Y�c]+F�j�1��m���a���F�"�=�EQ������i��sYQ,�z����ڍ*j�|]�<���_�9���e�֘�]ˋ%p�������������;�A_]ty��&hʠ��QTt��KF���IÓeI����X�ض�JFY�dY�GMI�W�%���G������<�5OUU�v5]׍�@�U�p|]yMY���8�U6oMi�i���Y���+����O�!�9��#��������M[P��<=;e�� �E��s`��:`�_"38v��A�b�^W$ld��WٶOz�4���ټ�xHYY�
�b�Tx;��I>���ϱB�z.�Ki��f�j���ҵ`���5l��?���c
=E,Q=b�X6�ߦ����H�3=XN��u�_�4�햳X�<�E�
_Hդ��(�Wk1
��X:�(�,+Fˌ�����O~�ӧOi}�f�b��LT�L,y,yQ�9*�xYg&Q]Had��������euq�/?��Y��3�g�,�5�I�~���)0��)_��>?��g|��_�o�;X̚�fɬܣ��j��_�C��/~�j�%_��m�@�`G�/"��Y��1F�&�8C�����˧���D����%��4W�A�8��2�|�!�D�"��߰<�P��9O�dY��U��!ec��~���y�� ՙv����{�n��c�_�6c�7����fX���dY/������o��ݻwy��w���;ܺu��2+J=z�f����������U���3�\�XV��lV�Xra��QCX��^���������Z??F�у���A�#��p�$1���hLMf2p��b���Q�_�W��!QP�H��QM^���9Y��ۜu�f�L��b����d�y�'K&�I.b2�JW���^ٴB0�"�)�N~��)�C�tmMYU�Z����QU3k��]�*s�͜u��1#��ط��?~}�f0ԛU�%d�r�]�|��c�Y��ږ�Q��W�f�Uf�jU����5��6���lfT�s�޽���/�l�ݻ�߻w�u Gu�LUz+f%BkĄ�D��$]�GP�\^^0��{V.5Zo�^�=UU�h�.�T�1z�>=���?�����o�4h�|�Z�z�M��=O�4�cl��vZmE��=�wB�� �nzy:AL��>��%Q���j�����jE�n�,/Y�V	��X|M`�<�7�+���2��1���ܚ
�5J�"5�u�=����!ڱ'��@4[K"�B�'�hVL��B������:�e;QJ��뼠�r2�h75�J�:b�p`ˎ�L���mQ0���勉�7��q���l��2�U�@LbOڶ��Ռ�#�����T�ٵ=�*F;Mc�j��ɖ4y��r��|�.�s��N��g?��䄳�?9�r�ĺ2u����9\��l�TC�^D�C_v�7ہ*����C>���'>C��e)����zY#d�u�1zbH�e-g��V,O��~Uc�ʉ�MK׮Yy��?��_��9G�ѐz��%EL�O�4�}
�<�F��<!��q���"��!u�5	XxLH�%F�@�,�-�� �ΧjQ��Q�1���t����3�������삾�rw��s�f��;�i1�n5���0v�߰�4M3j\��eYr���ַ�Ň~ȝ;wx������S�5'''<y��#'''<}�$IDbd^Udα��鹱�!����S��l"\��Ҵ�����s�ME����h�@HO�Q����'�*4>��:��#t�x�Z�HD4�&U���b�E�o���65��3��_�w�@V�bFUT	M��3��g�+	VEQfe���-���(������6_����w��	IA��-�K�f���]��B�AIsL�<Yn������9(ɒ�,
��84up�\��ǒi}�P_�Y���(1!�����ˈF���,��6�1�%��T�o����;u~����'����2zF��1ƫ�
	�mu�� �Ba-��E�et]Cy���z��Wcx���O?��Ǐ���P�8�A�T��\1J��tW�)?l�Tp;�wx}�����@�n:z؎�x�뇱��M�1�"�	1|�5��6��כ���r�Rt�b~I�;�M������a���6���k$�)�#^=�E�<g���J�M���\����V��CϘ��9g6�(���,Y.�����L[��:�+d�$1}V�zk�:�˔��6�Ib�D��A�4(W��q��A%bI��vQSM�Rg�������ᕛ7�_�Y��ҮVtю۩�	�����٘��,x��|����x�����!�͆��'�כ��i+��a��rA��1h20F�$]c:{d ���EAS.�fţ/�8y�����e�6�;3���C숱E	l��B!s�e��
�Ո˓UKpdF(r��j��X9g1��3L��&}3@DL�'�TS��JJ�9k�3A�@7�ov� A����JJGG�(iaF�,�e��Yb@b?���oۧx��9�g
�^~��n����fC����9oÜ;�����zF^7���a�If�u�W^�|�=n߾͍7!����>}������
>65��2��b��mq.�陼���e�q�&����1a�*��Ҳ}\z���ɶ
��t�-��ߢ��]��X	��q�$�g]�X�㚀!1���^�Q0�.��M�vE�>I>���l���׈��9�y�&��1cG�$ˠ���R�r���ɈJ u��yF�2��T�%�,f9�2cP�X�O��h�(+9�
K�}_f���l��|�N�1l��HJ�u�
E1��m!���9B�9���w�m �#��*���f�[%Rh�)�[���Kg�����7��w�����Y��k���άx�������N����������0ܼy8���g�<�mkNN������/��p���[am�6W�����s.//��`)B�� �)?ܘ�"��=�vR�C�7����ԎcwB�J��w������x�i/d_��,i�+��~ۺ��/;�=��{�{~�GR3���<�Ry�[6��V�`�6�O5�@:z4
y^��w�|V���M��-Ѥ~��& 7'C0Q�%7n�^�7nQO�<%����21��~���p�$M�V��h�5�Ѻ������,�Y�\'����C:�,
n�����Y-988�ެ҄�@�Oo�Q�$�#�{�=�~���{ұ����$�1E(-i1r����ʶ�r�?��'Sˏ���muM�u�[%�k�h�v�#OA`�2fW�$��X�HP:�P:a��G�u��k\!�'Ѡ�2wX�<��AN�Z�]�cj1�ơ:y+�u��H,t��(���Pa�$pb��A;\JBh�cRP#�}�qH3�y_̐�}^���~�+�kwG�7���u=ʑRox3�q�5e����7��{wg~懁�\����|�[��7��1��'D���3�e7�u?7m�]�B�D��XI�<�Ec�n��J���Df�\N�k����{'�="�:��ύq���e����Σ$#�:4B<6sxBj� 6��GZߑ�> �B*�I�#Ĉȝ�� �@��f�X!w�Xd�e�0E�Yr�a3�3��f1��t\� A!*]���:�}�5����.�t͊ns��| Đ�m�~���@^D���C�v[>��������:L�UU5� ���p�Х�S�3�/f][w��NC좏A�uU+մ���<��o�7��o���%��+������8���w��l��d��[�$˲dnC@Fd���h�Q!�4��Z@��4�Y�H��;�l+��lQdS$��*��>��{�W�����[,6�d�[\��{��s����������:3Ea����+��V��pe��$�*���6M�Ǫ�B)��#rt�<R�nx��>[�=���bI�?����G���`�e2�\.Y,}szk-��m���1m۲X��*�d��n���tQ�"���X�'ɓ���ٳ���/=�OS[j����%�"*>�inO�7��8��V+�QFf�$����c�Y s������{�?�'龒/��M��E�/]�D�:}�8�X.�ƚ⌣����^~�+7o��(�{�n'G4�5���ڹҝ�q��2v�PQ���y����-�w�,�K����R�J�㒋/b� >��3��T��v��Z�b4�=s��M^}�U�I�T5�Uloo�2��H�Ef�Hy*�1����-ٙVYgm :��m�7hi��[��� �!A"J֕�:E_T\��ʁ	ˣ9uh��꺽tr>�1�>t�!aRf���P!�+|�$��&֩O�Q�' ��������1:�I<Zi�*pc/v�`��v4�%t�U��6Fw�����E�c�>��
�g�&�;#$�EQ�sz�|��g{q|�kG���u��7"���+wS`$���Ʉ���hc*r��f�6@r ��>�9:����@T'	�x4�{߯��<���(ǔ�s�}��yR�Խ)�&b �،Q��I�Q��y/$"X�is
(��z�����fٴ�I�ת����K�M��p&�&t�=�x���m�#�Yg�T��x���!�5e�h��LG kM�mn�t�kޣ�f6_���Uv>�;�+�R��&9�J@ɺ�(ݣDq�����z��=)8(�(�Qh�O
o�|�4N���m��ku�g%)�b�7��v�g����y8���6�`�\n�j��R�a�VƳ
�� �ˣvw/���G�������oE��W��cV͌�?�1<�i�Q���NgGL�SƓ�
SJq��5���o1����8>>E)�1ާ���½C�^z�� O��4��S݀�<��M<M
k�|/����~�w�|MӰ���Ç��U��H�>Csr�À
��D���dZ��-"��c��e��e�x�����I(���ւ�&�Ef*xT�γQ&j�)>�B�&�:}�_�w��g`�g����*?EP�����Ũ1Z�)ѡ�Q84���*��U��u��	%,������� �#C�u=�t��&E>��[(�͕K/s��_���i�@�\���V�d-[eƃ�Q��'(}�>к���Ӵ�n	��V���r�EE^��$��'�a�jE�F��<�,6h2Q��튑��Tx�Ȳ��Qň���k�����OJ����]v������������#��=Gh�dh�O�=��l��K/p��7(��x�-��'ӆ��.��㼦�9:�,��� �
r��!U�nF�d��	8:�E ����ۼ~��ϗ^�1�VGp`u�!J�b�fg?���},�cE�� 0�.����%�	�Z,G�n
13��$lN���.�$	��1�����R"T�l^;�B��0�D����9�=�E)��!�t��Xaӱ]G<��iC�,�Z�3KE�6�M�~�a&�5m� �-�uEU�(��_���{ h�(�	�̡E�#}(pz�b:ً �$X����h�K��B8�+\]Q-��nUL9��<\���1h(��rdg]&J�>Z��fvtS��f��"���,�K�0:��y$�Fk���A��W��9�w=H.�H)Q�vx�����������c�AE
��cg��\W`��|ۯ��1d���sWW� �#m��s�(�ƪX���=H��#t�_�����t�������ޭy�!�u0�w bj��߭�Xkh3EU�m�〻@�n���
���g^��V>�˗������,����QZK�����/�M3k��f.�,��[���X���~[^{�TGs�:Q&[��G =�/^00R����]�ܹ�������l�����[oq��-����s����}�:y\GG3._�L��ܹs��x�o��o������1��ǜ��Fo�5�D�>�mvAaRl?������3Q��%�q�<�x��ώ�������A��/y�q�$ �g͆)���Ǒ�i��p�N$����˼��>���~��l��tL����nT�%�h¨�H��]���Q$ت!�    IDAT���ZK�t�g,΋&�s�
�����cn����I�$(��	�������C������w���s�Έw�����M�v\'7�g�$�j�(��4�(��mFcW�&�#U�f�e?�lΡ��t��j"1=�N/�E})���9�Ʉ�,��f(5�����⠦*ߴ�TŞ@�s�b,�E�&�u5M�hh�S�ȳ2�.���G�{��K��c��9�u����1%�^kF�6��!���v^��6� h��^�0�D�[���B����c!C�{T3�H}��#s�og���^i��A�1�����k͙�cHAm�ޟ��M_�Sy<�;�:Q�E1>�Q޸����sM���.�����m	N�:C�eUD��kc���7�o<J"�w�d�e$�v��܋�8�*ˊpp|�����w
�G �������?�C�]��޼Y��� �k��R��cVr�pV�>��5�����.�"G#4Պ�Ǐ����������Xr,QH#��R���n:����)z�"rC�B�*|�=o$i�����t�J���l
��0:8l�A��c�{��QA�<��8h�Fbi��l������,[�xz�*����rU�ZF�͛7��sz:��dƅ��Oڻ���uǁ�vc�w��^p.��<�êm�yG���?�����!��LS9J�H���ˎ�prr����v&ܼy������i�k[�	�CL���E�<����� ���#tabׇS8��Q�t\��6�{?c�o��yLrf<�����>�eY��|��QJWN�v`����D��<��g�1�Z6t��-�SB�ڵ����"h����ƍ�@�bQ�B��Oiac����u�u������i\gl�G0�5=�xPg�ADȳ���E�����Qx\��u:��Е�F]>m#�/�QVG�<4�9B8+~�;�f�A*���,������"Q= �MA�������ߪ;��<�FY��:��˝t��$f�b1�CY���F���mQ�>q͆�2+#�,�."�u�w��Y�ʺk�#73�U2B�m�Z�"�����o���j9�EaQ"���m���ҕ�!�6C@+����޵�Z���K�$�E�G�j�/!:h�1�`D�&`\��YU.\����;w�0��1�0�y��1"���1���K$�:����������'�'�y�7����aLy�/ے��CO�i���Mj=_�[�B���Ң:�H�{�����s�>R
$�u�Dzr������.z�7�{�5i}���{�|>����u�L��P!`MI�QAp��l	jF�j�Ν:�<~����ׂ��3.�paY���`�ym��\���s^ʳ�~wi-�c�����e���)M2.^��d2��e��:FZ��!�����f\F3���� &C�"+�vDլhR�����I�����>[�-�Zk泓/|�Cg9��ZF��ɄK�.���)B���w������D~ga��$�`�eU5� l��q��M�]��x<a:��X,9::���������+ ��M�^���3PQ4f��<���Ǒ�qڲ�k�ީ )5��1�'���(���҈�B'���X|P��<%����FcTWr���+�Gi�o�t����Q�%η��b�Z|PH��wxӤ1K �.E��&�4!X�b�������L��@b��&�,�z]�s:�E�.j9�?e�"�v8w�E����z݂5����G먣���UyL�g�}�I��EiqU̈�m��AME����V��Ѹ�W�9�ۣ�3�#�[��w^x�;��*S��sJ렻�k:r+
��'���{�6Mӟ��Ǐ{��h4:3�����t:�,�� \��q��3@+=\=PROO�~�J�{I�A�.���K��	`(�YeY��ks�9�=˪�"�@�QJ�R%�D>�ha]������'���&�,��$��v�������>�d�A9������~x�ӓ9[�����Q�)G6��E�ꆦ�c�$z���wTZ�z�ꊐ�wݤ"=Y��l(O�"���2��ֺײL �L�4��	=�{>�s������^�ҥKL&��S7B�:ڦ�Y�>�>�t���kb�m{{mjZ�ԡAw"��r��k���5�yub~�l���X�go�y����km ���ŋdY���Q/���Q�����Y�ك���O ̘��vQ�ƹ��Zr��n�x������3�{~kh[χw�X�8::���CNO�q.tѯQ&��:��d�h�Y�#%��E�b�61���T�[�4�o%��p(/��^TҴ�V�d�H�Ġ�{A;���(c��|���V�C��DmE�AD)�h|z)�D;�Ĉ��:u唏Jv�p��w������N��|'����	^�(�g��A�V���V.x	�uo&j�k��@�j� �R38F%�{q1L�<*"U!T�~QJ�6fuナ\� ��AwaU �e��Z�R!�(o��D�;g���5�5���7�m�Ci�^���~,"�d��cT�#c�_TҾ$J��.���D����+�>��ݰ���p73jn0�AS*��.�b�\�΍�e�|���I��h�?$�D�;���ӓ������dIѮaĦ���q�@�{�8�É,�8�ӳD`��ϥ�0�Coq��U^c�!S�p��'-|�&���`C��� D�D��mt6Fk������H]��{;���(�mmAS�hcQ6G)��9Y�DӇ��w'��gr����y�g�)�ϸ�O�cl3
� +��5�c��tM]S�Z��>����6#�
�wH먛��ZRU9M�p��iA	YQ��w��tBF���
��h���D�6��	"���f�yk8&���:cl����(Pb�nR�T��g�\��ߟ�'���kU��7�=/��uv���F#�˚{��������x����rA�BuC��y�Q摧�"�Q�b������x\�}������4.���*���.�j)�̓+�U�#�#"!��˃3�6�B������Ҳ����T��SA\�ֵGG{˽�����RY�}���De�5~���Yf-#�m0bt�G^S*t���8��ʊ�hU(��X�j��)�&JFi�%'�$=�L����z�u�M�h%:+�P�X<+�m;�����E0
e�Z�VDƙ!H U)%�U�P"�(gă2h���H�2�J��A�ZKP��֡PblP%�5�eZk/F0FBQ0� ^,J�,ӡm�>��Z���Ѫ��ӣ��2V�8����Ց����Z[?�,܍�dr�v��}�Mu���Fo�컂:2YvA!c"�[3�6�\p�ek:��Gwh��o�@�4<~���>ƌ�q���0Ĩ�V�>���9�ٌ�ju�T~a8mxF�睴��lP���P�~pm����I��a��a$q��F16�_�K�mʒ������OZ��l�D�(��f$@G~L/S�����M�w���{����d��$[����f��ݝ��&v�(�y^c2�9��}�ш�h�<� ��{�6���Kkr�9�{Q1kL�oK�hkk��ׯ������#<xR��0x��������-�|�2�Q��|�ֆ�V������=:�{��p^��+{>��3M���%��-t�R���u�z�g���I��'������m&*���>^�o��;o�����!��
�'�:[W��6��&F)3Ma.\�!/3&[1[���y�_�4.��yh�Z{�B+�.�������v����+���b�ֈ4���MF;�V�΍��b]v�4�,���R�UVm��.��x5*���3����o���_��Q����O�(�~�w~'�����z���۷��۷�J��}�������t��6f��R�c�ƹ�Nm�k��f`�UJ����{�L0�k� w�X�TN�h�>�,�*����*��\#�l�:d@�dNkk�C�Pʪ�����D9���s6h��Z���8��1GΙ\i��֫;T�+��*��Q=��Tv$Y�a0fi�ʴ
�m_���AV%e����t��r)�nݺ%���8��Ng�ڪ9Ɋq�> �Qd���Ն�ka�X�e{{{����������wI�(�F��szz���J)f�Y�oW��x|��ؒ,�đ�`f(�.�O�g"��?M6��w�Xd��3�9�ߔ~;����6
9λ?�`/�ֺKu@���Q�1ژNGS�N���}�o��_W4�Q�Sc3��N2�����۟Rv�q6/�F�	�������g?�R��|Ч�O�*;����"`C�+��˶��ӊ<˹|�ba�Px����b�xd���ĭ�H�{)6gw��l;�T���k��
5��Q��싷D�I4X��"�T�2�s��Ms��x|����ŋH�O���$SJ��|��z<���ϕ+W����㣏�����hm�K���!f�(W�5ň�t�h4�����x�R��|�jYc����\�x���s�}ur|��T�Tm+�r~$J���EU��AB0^���ki���Z{�6M�hT��f��*��F���fbmc��Bp&��[���=���mk�x��znL���҅������ (
;�sY6��۳���ܵE]x_Ε�lQd�z��������ʭ�n�ɤ�>�����7.2�im������ڋo��}���X?��P���M��,�q�X\�U0�h�[��º���(-
_�F�bE1c\��s����H���Y�H�@��X�\ �i��~fA+������ked$^��z�DNuΞ�m�>
5��⼘V�4�B��ʚQ�C}\Uvvv�yؒ�upppr��α������p#��TL����0S� ̛Z�(T���;��{���_����QJz�w����ۿ�ۏ�.��o�b\������-�7�#����"3�l�o�V�u��+˲�%�#�u��UJQ�%�ժo�^�6=����CUU�C��]�Uz^�^� ��� �
+��<Ŵ�a��@Z�=��E��(h۶��=L��57'�=��x�5Z"6U��^��%���15J�v��Uk�8����F����f�~Y�(�δ�Icዖ�I��kK��g|��f�=e2��)�4� ����	tc� 7e���Q\�ckk�+W�2�-K	䅉�]%�/E�Z�p���^<�|��ޅ�4����qɲ]��~�yE����bу�ƹ56�<�_���ñ�RcQX:�#�����m-��˿��_������}�փ��gJ�G��:g��*>��ӣWؾfI�u�f�b{w��w�f�4��X�������ϊsǺ�?Q/"�0F$�#1p�6���~Y��}=+���:�_����ܴ�j�Y]�MK|��y9͛OK����,��y�h ��^�\�l�e9�aݖ1uu�	����Ɍ%���;�$x�ݽmnܼ����'�����&��"0�n�H�R�՝͉�c,Yf���t�r��������a6�ك�G,���nX>>���cw�?�^�tq�T�#4{2s�}\�֞�.���i''ƴ�͛�	ʨ�6�������o-���\X�.��_�z����)��śo�)Wo�R@�}��p��������խ[�$��?�?���۷��q[����i�[�n��&��81��G�p�_v��|{�j�]��6׏.�ӫ�h�ԓ�AƩ���q+���������cK/n���T`��v�%;ń-�VK���YQ�e�L���Q�y���*7�(9����ж���8�Zoy�m�*�B�h�5tЂ<��h�WZ�v��o��.m�z�o�����t>����Z!�F{��2�����R&��y{4�O��T���O�a���_[��{�;�V�daU�em��j�7�~���P�h��L_nr!��4;/�;�NY��ʟ���j�t�Y���9���
'''����^k:�TB~�bك'�؆*	;'�2�ȟeK��	Зe�d2������O��[C~Q�����$o�sBw�ӭ>*����(3�>���u��h�B���Og��Ιυ�����|o�"�/_�j>D��Gk���}Ї������/�&t��|}���-���:��p(C��2�d���|������obm�\����w?���lxZ����Z>�w����������E��@v�.����1&>G����Z��OKe�Ά��������$���s�k�d����!t����p!"�����8�
�>�E�;ֻ��x�y�w89��M�@u��Hj�f��s��e����L&�y.Jf���?�c�֎�jI�liZ��DJ��X���/�)F�����rn"A���eL���M�����?�c� Z�Y/9�o�������7���|����}�7��称$���R�����۷o���}��Pr��n�|�p��5�����0|�ߔݺõ�b�r�ܿ~]F���|�W���C��pl ���t���N�>��ӝS٫���Ω:9��s6|��U���?s������y��ξw橺}��o����<�Gʚ�b�]���՞Blh%7Zc�A�`}�&`��k�h��k�w�F<�����-`��rN$h��$�L5}R�i8qE��QL^�P�15�NQ������������2C��tLÔ���kj���gV�ՙj�/Þ��?��he�dfY�Ot_��=�6�
8[nm�F�hm�6�茠3�����ϫ���믿��䐏��ؠ� ig�OS�𐃇�88>b{k�";�\�|��/���Ǐ1&���*�;ϔRԝZ{��t�H|��<�w^Tf�K�u�M�(�J��/�"��k�dgg�����?�0�y/8�e@�v�w�i��"g{� �/���׏�墦i<u�X,*���"����Odϊ�mF�����?�g�<ǻ���p�ĭ�4B�]���o�7�����������|7�4�`�Z�4v��4k���QOK�k�d2�{��f38==U���qۺFIl���E����p:���	�R֒�F������iZ�����~0|_YgO�ގ��O�?z��I����g�������+���%s��<�ƨ�J�C����R)2�Q�Z�c��nMQ�aUk��eC;�K?�;ϔR]A�Y��M0��)B7�L��<�{^�d2��ݻ�W6L��xs�J�F���1G_��tނ�,��������%����Z�96���4�*��E�X������|�/���������گr��>����U�B�3���̎�m�v���1<~t�������`w�W.�@fe]l�w�OM)n�Ϳ���i`o�vFg��YG���d{o��f����~�G���9M�8�ɰy�V�K�>��ݻ��ҋ\�V���u7��d�b��,+O𚂍9dy�Y ~��=o�w����ڜS�c�,J۴0P*n{8o?������4�V+NNN��&���cҧ]�γ���
���CB�y���h΂�$ӚR�%�{i۶�C���'�h1����g(,J.�c�Wa�X�Z��d��3<R{q6�^�ܮ����m���৛��ʾ4{�]�������r��ҏ�׳�LByn��+q���J�]2�c�$�`:O{_Q� k�6�Ki�a�5�!P��_.����V+����,y��^���i�i�3�жѻLಪ�/�����yD��'"}S��z�I�y-ݯ3i�n<E'%�)�����C2��6.\�7�7�������_��`�b9c����g��aC�����֭��؞��۾��9��Q�m싊���o���y�/����`��˛�g�=sJAQ�i}�,snܸ��70�PN�������o�X,��#�#vDц�4e��ʐ����#>��C2{�����or��/]�i�?�׊�d�	J������m��l)�5���ߟi���cꪔ։��e���\9
|^��M��2<uS�C��4��?+�w68��{�ɘ��^P�X�����Ƭ���Y��3�ǣޑv��Ѩ�(��Չ��RH7g��hC�EY���2�2U(�[�!s^�9���+�[b�&n��xG�2[��X	�f�F��|�t�Z)b;�4 7���;�"d�҃�"�	��7�<ͳ�\7ӥ�{m��)�ato�In�tC,�3&�oP)�w	FiA�.    IDATӾ7�߰(%�y7���h;oR�=+���Y��t�S4�y�3��m�c)�O)E7���Y���7n����_g:���ጻ����!YfP��9(-X�	ƠuL�<z��*ߡ^�ܿ�|���'�FP%����;�?��7ql����.��9[�z#}��4M�`y��5~����|�"Vû?>������?��>~�̒)�hd�@��Sa�Ay�.�?�����-9x|��l�h4�,&�W(,Zٙ����7�=o�����p���,����9t��Na����f��y�O��l:��U��c�ٌ�ry&��|<��[k��f}�.�S�EQ�Y;����4���c�t�I<�bKw��'`��G~�24MMTԳ4�w>2A�w����n��~�\�W�sjO��۷o�����!�V��^�6<ԙ�����iM�7Z��(5&�Ch�p�I`( �1*6D�]oǓ���dO{�Ҥ��KO�WaO�o��H�Q�}��[)�Wo��䱹X�m�^O0���,��Eq���ާ�__��霡�7k�N��p.6d�&��O��^Rᣏ>���j5�YΩ��Ѹ@���V�k5�讗��Ǉ8_��c��X�>�YE���t�U��F����ؤ(el�A*�\t�3 �<�T��F��OkM[�k����h�[o�xp�.o��gܿ�6����N,�<뜥��tJ2Z�@k�.62OQ�?�˟��g<f�#��P�<'�3$(��i��r�i87�\W���6���������O�<?3G� @KmS=1ߧ�|E`������t�S6g<#"=��yl�����ޡX� �@p�.�F��J89>\GJ�fT���m��bբ�� �
�VC%
Oӈ4M�
�[�L�Q���vF�90����)����,ٹ�Q�])k3/.��Pg�}O���J�Q!`�����d�ė�b�C/FDX���Drvayz���8�D�6��":	�=�Xy����XP�0�����0�;�,�g�����E)�{iC�/Ҟ�>P6��I�NW�ŧZ&"]�óܸ4�b���µt�)�lmm���͏~�#�̀��oO�u�B�Z�� �Y����s���|q�X�W��bww�</�>�is*g�>��,�"{���oq�ٟz�r7>7�8&�	����~������7?�G�<E�S������kY�jl&��S�(�w���ȩ�#���ׯ_�������cr���?�B���3�u���
�}
�S)c��E�R}TjHU9�c�4J�$@5�N�N��-e�Ζ$��|>�[�����9�a�#�L�,���<U�9���L��s��i�_k���.�l����YUUvMJk����s����s����S���i����Yn�	M���Z��nf�}��>z�b���g��}������~5b�߹2��������B����4���]�[�Xm0��j�kO#^<"�F���-1�:*yV���U�j)�:�������kc����<�ŝ��j�a� .�u ��􈭭-��'��R�5Vk��8�Hal���m��2�=H�w����
)LqH^e�Mn���� ��7����0�>�i=�d!�I}}4J�j�r ��/h��>��� �8�ٚ쓛-�Q��&4\���G�,���;�2C9�?~Ŀ{��</��?<,
l�i١�u���/��ͪ�����7�������]>:XB�^�ԒǇf^�ƉB5�,���	�v�-7a��<^=�n�r˪
 ��Ni���g_�O�JYT�G.��R�j>CG�ۓ4C��j��j��
5���|�Ο>)�n����F��j9��Rж5Yn�ti�w����?�x睿���nG<<<��m#���B>�3���sC�t4M���1���$m<��=3(�S�Q��ի�2�@�C���D�z�jǣW-A��8��*�0�,���S�4ԋ9�լ�m
<��&�B�0
�P�סu���in��]�������傼(#y�	�B�`	m�$p��un\����.{��\��C�@�\��T�GǏx��!����v��Op��K�0s-��2�C�U%˓%EQ����o�̅+���,�(Ǹ���vI�.��ӓ����]��>��	�r�xOfGhM�'�ھ�Py=�k���<!�E��W>�Q����1��h�s�����a:����@�E��<��IAr(�����@C���-J �Q�f�aœ�����Jk��y��"u���N���Zw����P����xoG�z����Bi�l�������WK7�������O���~��\���o���=�2f>.���j��^cj����5֢۞ �4C~�Zb��^P	��k3D�D�C���Z�x�}�6ӌ�s���\��e�G6�|J�*�,�X,,f�u]������"ҡ� n� V���(Sqq={��@Қ�xn���m3f�%J��Ձ�N���E^���SLE����Ÿkf�Tt(��歚Nݿm[=���½{�x��8<<�Q�=��hU�V�cMp:>'*�d*�x|h#�V!v�t��QT֩<?;�ƒ�%Fg�ҢM��nɣ�����)A��Ϣ��o3M)�	����߽�|�[����V@��ҁb�T��}�"	���"Q�B�M4����{���(���X,���u��^`o\P��`��9_�3�/m�B\�t�Wn\���q+�ݿÝ��`��j(EfKP��n"�����y���y������&�g�2�h%T�mUst��;����ŝ�����4%(KnZ%,]|V��x'x߲XԼ�����_����Wٿ��YD7�x�i��+����f4.�t���O���(�5�J��by��<�j��ß��ݼW�"��66i=ß�s����q�7�g���3���y�X�VH:x%X��"�y�T"�{�ӗY�ʾT;�����w�w�R��j]XV�f�ng6�&
�ɛ8I�c����'GqR�s�s)-���#�=@���
��k#�>����,A{�Ɉ\�OJ����ސ��Ep�6�DHN���x�ŋ�����?11}��������*bH�D%@�z.�����M��"�i�g4)Ȋ��������A+E�6<>����9	
c�و<O|��H=��aZ�1���,�Պ���>"�:�y�5
�"�4�AO^(l�vEۮ�"A;R"@z�;x�"�@��1�"(�r���+��w9\T,jG��,��UZE�a���go�c�a�~W<�bXձ��6�ۮH�K�� �G�b�QxeQ0Oy�k/�5E� �N����� l��2���ɚ�y����y�+��/�2�ܼ��*��>b1?��g���2d��ʫ����_�����^���S�?z�S-�q���-m�	W.]�՗�ί�����.��۱���)Ah]C>�c4Q�w���^fz�
[��x�wx��~��f��[�LV /�g/�t��|�;|���foo����и��ű� �5�0��^�0#���������;�NN��PZ�q�i7u�L�9�)���?�o��͹<�p�t�a�es�ߔ��<��-��=�:쬳XA���������n�h��X�쩒���X���$��|��Ai��u���kk�1z�m�A�A	��Q8g�u�IWu�G)Aa	�j��;#��^��<'���R�^a�Le>˞
��0���,)ҧ�ꏡ(
F���詀��MЗ������C�}q�TmC�^^��#��.b
��e����%`��Y�,�Ե4��j���Y��������������hM�+DJ�(�#]a��6Ɠ���5M��iWx�PZ�Fx�vh1���6*�"|�Y�"���`���~�%����:�V��h�Q�z[(�� �Ƣ�b�d4B�15�X�Ed5>�h��]L�J�Պڭ�m�����h[b�a�j����7��˯p���fww7F�f�UL�F :-��ŗ`"IX{0?)�6�[��ï�������������d>;��Š�k�< ��1Fs�����7��.�v�l9c��Ĭ:F���-uAqq����_�W�W���+��&�^@p��r/�����/��7v(&Q�6*�����T�C���8/�G�ܸ����	W/\fog	-u�6��и�v9��
�������gS��0.�@��f'BL�~��Ր��C����E�Σ�9����S@�y������y�o�3�u��:�"H�v�!�J@9	�&�p��͚�~����?����o�=��1Yݢ�Jk�k�2c�dJ�1F4�#)��#h!�yDp.����ćF��Ak,��`i��0x�o�x � 7�~'��>�ڞ�4]c	Lӿ�ņ�J��$�Vp���{�r���Çgdl6���P�ŚD����F�I�9��9Z�Bق����Q�y���Kr���LIKp��b^��(���2��5���D�5dV����P�U{���J)���L�#7��ޔk�.q��.���|M�V�m�-YG��#�炀����F��4��1P�kF�l��/q�i�Nv8||����U�����,Fi�����(�mc�⪉�������zE�j2cMs�<��CPh�c���=Ⅻ�^����J��y��&���Q)eh�Z#�}����X�<�(A�`�G�B���/���OQ�(�c����X���~�ݷ��|4���m(Fc�|L�!
��,˹v�*�x������%���K<ZTg���%�k9��|7���)�\�V���3޽JZ�|t�YՐ#P9�5��������^~�reP
��������G�G�mC����/39�Ɉݝ�}��Qd}��J��ɊŲ��ʀB�|����v�{Ӝ�Y��>;�^�y�\<�T?�ZO��͵j��u����ӂɩ\��UW葧�� J�	��ҥ����9���SA�t��
?E�Z+'(U�km�3�kl0J�lv&2`�A$j�:�����K�$Yz����9����wuW?���ְ���%��� �=;o	A� -�!�` pe�2�YX^p�	�m@/J�!��GwOO�����Uu�73#��yq�䍛uoU7��d��
�73#22"�9�������-�@���:�Օ�1�Cx���Y��QL�~Ƹ~��#-k1N��_�����Q�ũ��l�<����9�#��:��?�������C'����#b�H�KPK9�������X.��)�E�`)�
c�we��'%��s��rs��Qb����I��.m�0�l0T�0��h4�Kk˽�q�˗np��y��g����7�d���_]�J>����EL����I�=J}qcs��|�p�ڳ)�8D��'�]���gOJY���ރF�g�J�i�PVfU�j�X�P�:b0����U�=��te��J��bZ����3 �g�N_�S�&0m��\�h4��2�3JYV�;����7���J�RVc�rD�=��PE1��¸������3����u~�������rI�l�}�}>���N7א���a
�_�t�+W�����-`�\����K�ˇL���/�����+��ʷ��[��)�o}��������98�vc���/"EQ�������y���v��8��mv/^e����]���"�)}�qWb���K�
ﮏ�}w���y��������z�����ѩ�ߕ�;zdH6W�"bQUU4�Z5z4n(ԟ����s�ν؛��Z/��}a��3co�m�s�)�(��9��t��J���w6 5mk��E�D�K���H�1�`�0,+$*N�%��@�Ā3��Y�!>d��Ͼ���\w�㶼�<��C�GGG�t�<�f0�߶���&�Riׁ��`��m���FM�%�sn�s�����J�}�l�Mݲ���ݻ{�
;��xV�.]۬�	+Ч��iq ���KBlq�d<�Q8<�5���8�M�֭�%.^��d���&��$�C�E�jf��>�I��"R�c&�{�
�VL6�lo]F�"QY��n�,����QU
SR�I���RU����!��h �jD
���\��<>�2������������Z�����M|���>{g��I"Q��;��u��-��Q��5X�OKA�C%�
'a����}��6��!"W�6D"1%�p��3�ʯ�:������K������O�џ�	��G?���vl2�.js��5�?�W�^��SOq��5F�1bK6����"BԂKW��ܳ/R�D,�ٌ�{w���ko������-���&��5%�bI]�4���hƅ;�%˺�	��{b:���~�+s�	� ���t�����C��}����,JN��o�m�����$2%͓�gy���Ĭ�`�QUkQ���drG���>�_��{,�Ȅ8�ʌ���ZS8k�%���%%�cde��5{����a�M�W��6���H�'�/UU�,ND�ˎ�Xc1ƥRf��x��]ξ�o?���[�,�lv�}ܶ����{�eh7��N���b��&r���K@&�ʔm�dB����q��1���|�!��S�o��{�S�<�g�c��˲�{���3k�K99��ǄV�u���>]�[#�2�&4M�F��h�h@KP�2������4��A����ѷ�2����D\$i�<�2�UИ��'��Պqs"��1eK�l_�m�$��u�\�b�2`d@�J�6�\
�p��*B<Fc�].8����s��]��T�b:	 ��sR:>��>9-9H�YV�)kN��m<��X�X�<�����&��J'k(�u]��[�˖��&/\��g^d���t:���f�C���Sn߾���>�����m�CX[P�wo}ć����6�x�%�ַ�|�
���8%�u��α�{���m���dv��{��[?{��{��G�!˦A���1��n�ܾ=���?z�g�~�ͭ��r���f�(+�i��|U�	���?uz{l]߼9{��b�:&�,�^�`���w���=�x�DE>���:8@0ƢQ��v��_E�R%�D���Ύ���~�'�Ϩ����vt8�gM�=k�;�^i0Rc�#"FL)��J͔eM�4+M�b�|DGa�Ŵ�8����""�(J.^�e2���ܺu���^R/	D���c�i�"��!�&su��pѯ�����2�=a��\[��s���#�1������ں�p������:)+&Q����س���0'GN'z�y�
���������h�ӕV�@J����ضH(\b����рyL�\)��M��[�a8�����'+��n��8�1 ��;e�Z8V�C
/+Mwo��Ꚏ*�7K��1�+�i*�7M�~�l6��n�[�PR/�(�sx�4MK���ǶAU���D�+���9��7_��o0�G�.��쀪�N��|�g�í�e*�ý�/�u��da����Cvv�S��b��(-�G<x�[4�&��WQ-9>�r���y�m�}�����K	56շ���CmQ0�����9�� �:A}��e�6*M�1�g�)lnm�s%��m��j�]��E�@?����@z��j��E�z�iA��2ٚ�c
��A5�i<�3�^��_�����[�mˤ2�P�Ĕ�g$`բ&�1P����s|��k׮��������p<_b���X�h��b�p��.�i����7�:GӇ��nP7��2�r�bI�m�lǷs>����xT[�-U��	��<9RSũ1W$�D/�G��yj�����y��7����!���:����>˷n�����~�мȄ����,%��x�����}k�rs|h՘I�X�{�������O��l��v.�{8(Km��
�p��ڐqU�Y�$�u֡eI)d��]�<�U��2Q��M�\��G+�(J��91����
��|�lv���>�	�BI�xM{��D��:\�J��9]�w2��t�MӜ���癥˝438ι�d��Nw�0s�n���}��u&��?���w>��x��d��Y���b[\QUɠ5qUFsU8Z��)��{̎7G���e6�i�}�w�������Z���Cb�b��Sɶ���~�V�6��9�H)�v ��K��=    IDAT�󂢌-U%XI�/�7��t������;<|pH�R�$6Ɉ�J7}:���Jr��pq4>�w���$�����`�h4�(�����Ո�0��T�w~���D۶�*�*��?{t�\��loo2W��o�펊���/��4�n��0;f6;b1��6e:we���;I��E�^(�c��=	��i�R�PI�
Ԓ3�U�O�7�O$QM�1��TU���:��,.��Р0�D�cQ�?#VI K��t��3��z�J
=��!�HE.	��ǧ�j�d�N���X�Q<�E4�8�H�^Z�5�%kEmm�$��j����t���ھ.�_1���]_4��4��c�z������L�X��;�(0��e2�P���EY��D�BB�T�W�bF�������k�w�F0��11��Q�D���F�Z�4���UgQ$�rY�U�ӦiXV	��m �S�0�k;R�i��׾��?���O:}���aDR1�ު(w³(�b�Aۦ�;;;lmmqtt�b�X�Ķm;�x����\E�{��Y?��V�
�e&�_�h�#��We��t~}��1�����1�q:��y���E7����ĉ��9�>������m�z�`9;bw{�A����s����{g���;;h���뀿[M^Ʉ|�Y���xc�y�Z�A���Bo`���r�<-���$c0�uK��>;:���!���L�3�`�vL4�95!�Y[1)�0� Q�<�xz��9�-0Q-�VT� ���E\ǔ��I�o�G~ͷ'���S�J6|��U)DS�w�UG���,t�p�V��(	�&�G�g"_�nO@�k�K�jQ,F\yS���ֽd��<݌@V��dEJt�
bH�;yIo
�����&�Fl�RFULt��$�M獧���g�@��1QM��Jʚκ�cҼ��P�t�"���,M���,@S���M ���q���5ޮGU��Ԭ�^`92c�5��n~����������"�ۧ���{#Glr���QըF뽯���u�ʐ��Ȣ��E�	��_��{���l��h��kj��%�+�����v,e-�25�%�cM��5���q�Ĺ%m�2_$/�A5�m��a8�
A5p�������H
��h�Ƞ�VN�3Eߟt�d�Y3`i����]nܸ����*���F���E~����_~���x�^Ɯ�M��h֍���5?i�R=�˸��g���iO�%j0�+�6��xk~ĝ�c2�ę��#�z��E�.��{{ܽ}���}Ignӵm�l��9W��k��m0�~N�6m۲\���6)S]�ǇH��mX֋�6��i��b!�[�,ʑ�M�H�,��(�/+�(!%�4
�8*�E:%z��6�3��$4���,yf�������мc<M޳�kڦI��8��J�� �rzA#^#�J���q�"Z̟�v�IF}��tL�t�F��
���n��u��Xm�+!�)�!/Z,��t/�x��K<��M�Ĕ++練}W��9���Mn�!��_����
�I�e@L�J$6(.�-&� �&�W:��*B�#`L��e��"]Vsx����[N���n��[�������ϓ���s]β��gK����)���0�/�1X�Iy�Q���c�Z��n��E�|�>f{|��L#VU��Ԃ4U�/A*��t2J�Z�B0�	>�"cbǊxr�+�sFՈ�p���)ꔭ�Lg�<����w���/pt����{��ݻO��:��N�/�Ϭ^�~�Y�,��B飣���N2�����ѩ��l���������s������ڧ~�3y"�p8d�X��˙A:I��x�ܕ��E��ΘNۗ�K!�\*ki5�8>`~t�C[a)� �6+0mM��ђ��Bʮ�!���٧��������LA�����m�jB\"&�
�u��䶟����Ҙ�#c�M���q�BL���R�T��K����4�,��X�5.U=),QS�L2>VK
�8Q:�����
N��Oq��º�C3�C����FYU����X��;�I��<�:�b�ˠ����}��
	jL-&`5M���N�������8�>�n��A�²��&+�&�E�H�`<I���\�P�3�M,�1մ��k�twh'l�E�I�ӗڸB��x���S�IxS�t����(�2(v�7џofVK�'KD냾�����Y������������r��Fl��}F����''�ϸn������*Re��,�ъ��x�4"̌m� �ۋ/BVߗ�c�'0}����j�O6�F�xYSv���F�R�
c|xR6�����e�hV����;;;���k��|�����&�	ՠd>����z�rѰ�l�8�V�&`U�,��Z,+�g�a>�����b���J��[���j 'U�4�c�`-gg@����,DO��;k@�"��~[�5��1i�������&�D�3����%�8l!�o!�
�@�HL��F�h1��L�E�4I�^�hh�TǖΔW*��^*�
E�S�$��İ�N����Θ��Y���ghi�b���,�N.�ze(��I�H,F�Nq�{�*u8Xy��{?�IY�Ic�!z��4�jK@ X�8���s1�b
�kH��D�X��[@�O��c�u�}&��l�2}��AC�}]���L{��r
�����jNd�;��a�3U�0E2�&U��@$1	$ÞH4i�ŷ�U�FD�">���b,���B��+�gH���;�]�ݑ���%1��0�C����I�Zs��Op��Aߺ�V��y��o��|ǘ��ׯǩk���~\����i�q���y��ַx*�3j���j�Xc�a�%\d��b���e�B�sA�tzE'�N��G�APO�����?��
VI�&�
]�\��c�cc#�lU���[o��o���\�t)�������������Y��(���T�N��*v<|�p�Y8Y�z�W���;d��3v�w�W�9�������'2g��Hh��h���Q����t��<��}���_����=�ɞ@m�]b�Jg!�2݌PR�Lh �� &`b��M�8am7%��b�w�o�k���_R�S
o�t��$�� I�
�J�4D�D�'��N�f|X"�슧��$���O�7&%�k*����Đ,[\WMG5%�� ��R=\���c�`�&�!�im���&��ݦ'T�vá!�F���\������`pj1e2ê�Đ�N�Q�m�����y��;o���k����U4'a���8�l]�Q���5�+�䟙A����S߰ޘ�?v�tw]��d�1�99^%%Y3�W�I [$+��eW
7{T��>g5,��[,�.�����9Gi�� �l� /�'����xw�+C,>+Ě�=u��`�ց�Y���y��B��\g,}g�c���+���`DUV8c�1VC�qv�"�p�h���wŪ�K���Q;�]�:��=E%���Ah�8#���t��-���v��y��:�`���dBU*GG3�ۻ�|�����Y,�Õ�i8��/r��e�����Ν;ܿ�}ˠ([f��t��2C���2c�����fh��B�n������g ��������=�!�b�l+�{�;�}ј>��][�+TU��]�P����6��EA-��o�-�2o�nM��dԢ>U��@��r5=�F��d�L
u:��&9ƈ+:v%�41R��#�׮�+�����	��~��VU�eC�6����/`�`]�(�.I:B��[ �`c��h}
����m��ʤ}5��>�QbL�/�`�+Ř&OԆб����;�I��bt���A'��+�>�?�yzb����*���#�rw������YgwO�k<m��+2�H�L�QQb�ћ�`�bR}��'�I���+ �IV+10'�;�poDc���KC�I��;O�|�������y5�巜��b��cy���g�}r<���g�_;+BsV�(��o}ΥJ5!x�5��c��	M�����7����:Ř�&�2)�������S���l��v.�����`&1�E0�F5�^�7���Ƙ�~���0��T3�<Bh}b%�j'�� t���hs��9f4����n�������&}t����՗~���[�xq����|���{�{ꕯ��dbT�|��+�NUW>Wg��+�]�;:���1��:r��#�����~ˬ�j2�uα������
�>n[���xU�7g��{�U��mR��xT<1Z����)�	��XpE ���`:;��E�	��]����g�V�ڝ�'�W�0�_�Aȓ�Y�K����d���pJ��Ԩ`I7�ѐ&�2�P#fD�w�ͥ-��UI��v�%b��u��<?�k�1��u����Y�_ak�E��t�DR �m�K�S���z�fxW�s���哄���bd�)7���@}�n��ۯT���-��6������^q��?IX���%v �v��4�$�r:�#���	gA�S�$�W�����L2���OK3�B�k��}���V�# �&��9,i0EEӂ1���@S3
���x��2��c��q3�2�7"C���K�_-�À-��Ō�[;4�R�kv'����fH45�)� Ô��˸�|��h�u����#��c��,��.N4�����$��˼�`��d��Ax�jk�p��.1�0��l�mB;$ĂڍY6J�~���­Ch:_)TlWkA�I�$1B�uZ�k��0� 堢�*|�Kf�}"�_�3g[٫/�Z��!�r�Hظ������]���ǝ
g$�B�S�Nk	�j
��q�H��4���E]����;\�t����������=�/�����s3�y�g����'�����v.���ى��)�߫�jEP�Jie���Z��:��F�;���3�-988�iF���!��>/�r���vvv)˂�tJ}����ի<���:�����c{{����GB�O
q�5�v,ow�����}��Y�3y^8W�;�ugc~��
f`��/g\gP�}���U�izN��az�?�cߏ=�!�I^��ʧ<���X
�)}�#�Y��[���Y�~���)���0L�9}?���HA�z
�Pز hK �k�C66��-8n����[���g,.\����|�%�ج@*�&�RT�;�`c�.�YR��;u����u�����\nQu�M=��=�/]WO���!ee�L�eX��;�0�K�zsG<s�;�Z�s/��rx��ͯ��W��
�+,�����~�[�7�~`o_��,��a�F8��J�X ����嫴m���{\�v��}����w|�W���Wee�����@#
[h1qf�x��ח���}����޸q#�m�y��"� RkJ���j	�Ɵ��q��t��2w^�	�3�p||̃���u�dr��G����?���o������.�����Y�7����ڒ�(�r�J�]FȜ���AOX�Eǯ���?p��?�K:��b�&�����	wbS��?z�EO�B�߳b8�4(<�~�-��-�b�2�z&�K�^�������|+u��3e�ѝ�~XىH*��=�V3]U��kҎN��S���i��o]�q�ϟ��ڢ#	�Y%���$��n�,V�,�Q���zl9fs��q���!���H���%֕X;���H`<��5�˲iPM����Г,�Q���%���P�����"4U�1����s�uU+X�5���Z���5��%�	��)�%A5���#�0/'�Q^�k�>%Jb���'2����_�>���l$��_�i�@-�������K����?]��ܿ9Y�w6Mr��
<>$������D,��ߥ������7�����d2����?���q|<�M��EӴeYVQ���HlU�i[��b{���e�B��f�n,74�&��H[�i)2G�RU[M��QU��VTN�T���:����ASČ�Ѫ�fs��e��px���k��s��U9fP�����N�ݻǝ;w�L&\�|y�ӛN��t�>K�;t������ߏ�v���e��������}��{���_�c��S@����ǲggl��j}���Q��S!���>}-c��O�2I�g��u��|҈����Gx���u���y��9�><���Re��>(����@��{��k���>���a�/:�%��D��/����S�K�� e�ŕ�np��5����̨�c���S�o]�JA3]2Y���_����M�B��*��O-z��uD1x�D
p�M�Z��hLY�ƭ�_�釣f��	3���@�E�Lb���'[1�k�@�!�-�Iv�j�	,j��骫��-�O�����\�u�����Z\���~��>@̥<�����=�#V�QJ�����ژ�)۵L��Q��)�[�<���/\��'���w�r6��?�F�F����g���x��F�>�H�=
?���ѧ+��e�\�sA���������E�:�u!%nȑ��*^U�*ASC:C�U�w\�L�ٳ.�RX̑+z�z2r��-<x���6��&��pLQ�)}�����u��i9��[o�|���z���:��g�2�9��Fn��C#9�7�����~bM^M�e���+�Ē��	[�uF\�7V�I��=������$�������r'ӌ����g9�kǄ���:)������}Z��^D#���]Z���Q}K[/y�͟���S�˘a�`p���ã��ܾ���87dkwL�i��-�������z�Kw��!������wߡnTO<��GZ�u#�@aS8�,u��:eoc@R&��l�O��1�_;C��5��B��s0E�+�P�T�ͤ�Wlh0aLԐ�=1Dծ�!����h��2�N��9ۍ��>�g��_�������Ҝ�ѷnY�w�y����Ǔc:�8{�����n�m�(+bT�&�o����ʵ�?�\�����H}�\��nx�޽�nw�b[��C���zUDE<Q�3eq��|��l�������_��M�֭[�+���\}�@����s( ��X�u��ߏ/����֭[���y����:��DD��?��qm�M�����j��F�eT���P��,����h��S�C�D-֔�XB�GC����������
�;W�پĻ�!����)}`��p8<�1�����H�|>˗�� �Y����ڼ�q���g���Z�h�rD�g�����w<-⪪��+�׿&�0��^*��=f)�(�~�TI��\������|�Ӯ��J�;���߫��||$�˓��'�\��˳&�_�w��67-Plʎ]},US����o�����h��k�|q¥���R�Qmy�����!�1�ł��+|����W����x�*�shU�\.�O?�?�ɏiB��
TQ">*MT�
;�nCD�g-Zv�%��Rv�*���m[�!/^d{{���ͭ{�C��� !�H*|]PT#�	�(Y�|hS�{R�$�HO;7�L&���7(˒�tʻ������^i���c_�@__j����c�ia݄߯�;�{�f�8��eM��,K~�6�ؓ��k�4�C~���L�\��'�p?�?8�z��O_ڽ�Еû�ãoq�������j��h�r����[���h�Ϭݼy�ܺu��n���op��ݹuK�_��@�y�62����U�P_���o~��͛E�M�`n޼�_}�U{�?������~n޼i�� ������z�Bw�N/\������E�p�:���������Z������GGGᥗ^
���w�<�����h���=�;1s�F�CsT�&����#�:�(�ӝiW1ã*X���\��y�7�/�گ��y���b�Ac�2/��-�����{R{�w��Px�wvFf���5g�<x�ߵ���qL�)���`���$\*g��_t��y+P�\.QMY���'��V�	����S���~���7��-�� ��#�r�9�ڱ)�I?`�Y1ۻf����2G_��2w>�
�/��ϻ�?��!��W{Xm�g����N��bwW�    IDAT4�����#�#�[�O1(6�r��(����;���䭷ޢY(UUp�+7��K�o��l����H��1}x��������oػ� �A ��5���BU�o_��Oږ��i��!��t��6b�ٚln������K/q��U�����kNk���h�����l��:L�lm]��s_g��s����ǀ�M,�I�ڳ'��W�~�:/����ܺ�Ç�<|��Tbŧm}��^�2��斫>��]x���ni���]���Z��p����e�z
�|�"O?�����)�W�v.����u��ۣ���xn6�Q�����L�b�+e��Ԉs�w6P�!L�o�����oKR0����s�)�[G
��`�;qoq���u�������9Y�	M�������^{I ^~�u��n��@���\}�+����Ķ�9޺  ��L���y� 	����tl�) �	5Ќ���rA�����a	j�_w�E#/����͛���~�e�������a�ؿ��! �H|(�O��ݺ��2ڑa�?*b�{��{�˲�"��Ht�;Ｃ�������Q�����*�(��XЗm[ԧ��"RG�V���q5	�����V�ie����{�:	�@c�唷�~���S��;���[��S��s1�#��h%�=ku��t<쭷?Zg��]}֭�ֿ���yL��1�u\^��_�X�����e��gn_{6g�>�=)@���p�դKD4yΉb���c"��H�!gN>��i&]b��~�_��3}�x@��:���{�G>z:�:�/�b�̧kc��ܹ��]�Ե�\�x��4lo�p�ZIQ9666Mvy��wU��o�5~�����+ϲ�<�ǲ�y�����������}���6�MR����Mb�)�Ոrc�_�֯����o���t�ҕUJ�e5dkk7��+��7 �@m����ä�>�|���]��$F��f1]�8^��������o�w�"|���⒢H �(
&�	���\�t�o��5~�~�?��0������>n>��>�̶]}��`�<�:�1��<+�t^;}_w��c@4U�bS�GUÊ�W�����ln�|$���უm�}�k�ݿ����n򢭎�iƣ����LhC�3�R]e�b�����=�'���?��!$���͛�$z~FK���^{�%y����֭kr��m���y/ ��Ƽ��X.2fr<��ӳ�����/����D_~�o2�V�.����`�z^/���E]U	��K��+��m�r�	UY��~$US�c$ �F�	CY��m!�h����y�^T��j��ea$V���R�S6�����Z놮D����V���6ŊB)��.RH�"Έ�a��Ęo�����b�ۑ�'������'���B�Z;zX�U�����w���p��M��},���ى͝&�u,�SU�ѫq� j�i�v�VVˢ�Nb*��M�u]�4~e2�+g@�6�L�]' bp�ć��Q�;��|�`g�2/��Uvw�y��w1����,w������u�v���s�}�m��Ϯ�;�\U�{�r�\���5�����e}[Q$ֳm�UH83b1��NF�`�;N�
ׁ�,`N,ʲ<��}�����{�o_�G�1����Ζ�@�7bp�2���FTU�tz��d�]��K�1����*��E��
cW��'"kш5��#��ćh��I�v�-���A}�hR��q��x߅�K��&����Or͞t}�lE������-"�!����bڞ������-t>	�[�3��;�N��s'>�"�����.Z�3�#�{o�.���=�ۿ��F�S�����n<��zIeGLƻ8�}H3S�7�����������3��S�uq�+*�Ұ��.��?�{̷�_|���A��k_�j0fk�����0XW�\IQ���^���*���7ٹ��r�d>�a������w��.���7�b��Ʒ�O_c:m�ؾ�׿Qp��g���}�>����C*�E�
����|�2[[[�E�1p8=��*�޽�|����vY�ZV�zHz"��L@���u]3�1�HF�ѩHD#�}z=���#��xU-*'�d�轧��GBh1&eE���`�*bPE:�m�0���~1�l>}�ҥK����O�H��������ϗ�[�������m1jcۺi6
W��Ъ��^����v����տ3�b�x��A������W����#�o���@ �������ZJU��V�TE-m��Jdo[vؚ�u^���G�~;��33�@G�)�V�h�������j�6�+�_�儉�M�)CJ��z�CE��h�X34"v�Ī�¨1�Ɏ1&��� �1��Hcw��UF�h�NJ)��F�T�7Vŕ��B�
����/��FS1B�9QI��(�b.����c�U��{�1��J�$��9KԈj"��%�?>|��;��f0(k���]1o�{�e�����"��q����UUm�����><��������$�I�[BC�Ӂ>�^��v~mXn�@c�m�aU�@V�x�z�]g�B����|���ĸĺ���>��./�E�r�h4�|��+'4џ�2HȃK�Ԝ�zM�>y�/Z�����BL!#��d�cS��XGaEY��mp�`�T<=�7]	��q&�+�D�U$U�ǈ���U�j�&��Ŋ������CK��}g,���kJ�݂��l
s�Ɣ)fU�U>3���o�"��b�w ��j��ekg�2��$@2��Z��cm�u��^��Oh�oN_������u%��h v,r��p�w���w�������T�
��&4QM��p��S1,+ں�駟fcc�b����|�������m=�G�6�2�Lx��g���a�\�\Ԉ�ˆ����~�����m��Q�>���{�R��_cwg���-�����6�����W��K�N�-'c[�-���9��o�����'��5=�ym��}4�����0�%8���m������?3��W���̋Yc��g
���ǖ�%�,Q�:���Y̗�8t�����n�_�n�AU��h4x� �/^ؖ��-�ҍ��[ΚƔ�T��Q���F5�\�/Ն�YiŗfWd1Y.mٌb#��P|S�2nצ�%���cql�غ��3��`�C#3��c�##�����DA�v �T��0��m����hCB,�ja��0*Dba��P)*ވ��6D�J��3��łE,�(�k�Q��M*Uh�b��(xm1Q�xL4��8)�-�q=�D�U^	�Z�$��hX�c79t��=Fl7����|"Q�JFa2i�ȉ��b:���Xi�t�T��,T�:���Z��ֺ�lCx�����^�ڷW������WL�K��R׷�����~�;�	��ED��{���klZ�N�6ޕ��|�Wn��҄`���?ab<�1����?�hW�ҦbھMu>�*!�T���o����~���;�ۧ@�����3,���>��0�:�x۰�r\7�NV'�Z�? �͠���
����_Ɩ4q�B���U��� �2���d��d4���%�ii��K�6̎���b{k�j8 ����V��ʌ�l�(�#6-!$?���p� kS��������ɴY#8gp��XF)�W����s��G̎8:�&�Zr�zM��ve�>�a�g���ON���>���?�<������Z�=�qw�C�F#��qVY�,x�`��~��s<��|��lmn ��m�x��2�s��}��?����G?��G0��(����cBL&��P_Ӵ5w>�,����W���^bs��h�W�C����#�{Ɠ	M��=>��V�������;n�y@�JWR���ʲ]�`���ɐg��A5|��xBi�Q�BY���W���z��\T�9ӣ#�}�O�ٛʭ[�0ư1w���	�13��9��#(�儹�������G�����l�Lp�b5⌤JJQS�@��h@�*<���(���h�����bkk���.5bE�h2���(�����-�_�H�ث҆�mf�/�Rc��f�����Q5����8�1�oC4Xi%X+�x6��v�q�k[� ��5
�p���'�W#XREK���FBT�i	�k�cpEAT]�1�h�����)�����1���1��dzL>[ɲ(
����MB�iN��(���H�(�����<���x@�%eʧ�4���S���7��z~,�%��9,�n��e|�ò�:a�h��l*-L�Q�vP���I�K��Z�����z�1�V�ê�6�Ν;<��4��W��\�uӨ���=����,��* P���	8	��X
��Т�Q/g �*b�6��T轡��?}�M���ݹĥK0����/�ı>������Y���9�Ұd�q������3}����`��Ƣb��l��8S�6��W�����p��.�I�d8��-A-�i���m�߽�dk��y����y�L��I�;5)�k
Ga,�+hb���X��eQ`]*AU�m��&c2�1� gk����7��$���>g��{o�YYUY�7�E��Q�Ƃ4��@���������E�e =Λa@�0�a��戶�#Q$5����ޫ�����.����q�fV5�ZlJM�Hd޼Kč8���~߅v>���y��[���}R�H���Cj����Ϻ]���ϧ�>k�����c���p�Z�72�u$�X�����֏���c���Wv'$o��C�p��G����-��7����+Wv0�,}��R�m�K�����-G���4-J�O�_�am�)ʂ#]��t��PJ���q/�b	>���������>MQ�� �cL�-����}f�1�g��S�y|� �uG���Jcl��N�|t�.���w���b�]��R�Ӑ��R��/'��X~ު%�Oz�R��,P��5����L���>|�xTR%ZChm�$���,)^|�y��^�g���}k5"
���c��'''j6�G�Ь���!xΦg�m��S4vL�>4"1�I"��Y�8��ql��P���F��Ry�4)��Z&�Y�I	b�q�齂5Z[�Ŝ!�k����b)e8���^�1I��L��
�"Ď�d�QS��&��cDooF���~�1�R����-_C��J��q山*c����,ӧ,)�?/R�$	��N֪�bAb1O����w������|>�(���q��5��L$v�m=�RZ��{��ۇ{׮�ͺ���Փ���*����S��[���~���KӅ�c쒮�Wj�B��4&��Rk����#�e'�%�sw���$�a�i���}���4H�n������h������2[�ns�ib5���>&�|9�S*[�el���i2mC��I�����dl�}��aP�p�7��˽ֱc��_�_~���]�a�V2�J���ڶ5,�sl�c&��{�y~��W����l�R�y���~}pW��5Xm�YJW%�B�ǐ�g��aB���8g|$dQ�����kLF���~�Ǆ�e\!� �V���$���Q�iړ�u_�>��.�o�U�Fಜ�z٠�ؔT�АT��<Ea��-'�;4��t�l����?z��+���r��{��o�?�/�e\e��{��)�fOX!�.�ܑ����]�����]��\�5�_�썶�F%���:3}C���pŘ���[o�g����{� �|�J��y�Z����)�t�����%��]gsm�����h����,jR
4������~��?���Kl�<v�O;.ϯ���mۢ�����rQ�K��sy|�s���{>{��A_�R��g,�9��o��W^��g�ak}�_|���66��>���C����͙˔.��E$,�?�E�0;;e��7S0�L@ �@m۲����%Qʠ�,��Ƹ�{6nY�L) 1� ���t�A��kT0�0T줘mHR�������A�)k@�����rp��2lF;��,�gȃ
B�������(M�l$�\*5��5]�0$��2dKt��yã�]�o�s�=W,�;�FS6O�èIHʙꔲ:I>~ou�7�DT)�W�@"=!�tm��	Nk�LֈX�"��+���>��i$v��cR�h�"�d��y�~
PΟ���Z�f:�L���l�b$�K�D�T2�U�2�s���灐�b3�q�Z���l=�=��ؕEŃy�G��r���X߀Ã'3�(��U�����=8s|Ri�ݡ4�*+�XIL�@m�ȡΟRPy^jX����Ӷ�c�D�(M�\:��a݈�_�%����x��g)�����SG���7�r��u�z����{x��S\f�����Z)S8�����=
ED�mA"���\��~�|�����o�)0v���-^y���%�D�,z�]��	�$$��3l[[[@&E5M��p\�,��� ?����������MI`�j�DD��"���[�u�l������c~�_�����IL*�IM�g\�o�X���e,�AE!rvẋ�}��]q��1ׯ�0����U���m9;;�YM����;��֛|��m���ZML9�D�
�I�tDbJ�2�[�ܻ��ݫ�nl�QtmK0��D
M�/<z�����cP���5-���m�t���@oU�XfE2p`K�ד2}����c�����o8ހwW2em��ս�vm�/�U~���ʋ/=��x�o�I1��r��=�ܻ�b�@k(]%9��B�U��$m�b���6@@���uH�h�~�$�L`L�<��>�ڈ&�{v.E�ҽ��ܨ%��h��!F ��V3�0;�^�NK�z�(aI�QY�{Ũ@kM��sMU�Y��UI�JΦ� *�K;���ͥWb��A`J�y��HKJ$���%��m���zi.��/�����BΚ&�
D�Z��lS�\�>Hv-�]��9��$�m(J�-T0�E��Vִ֕�n��!Z{"U�M?x����x��:��e�ү����Ԡ��͛�����b�C	�AL\H�_��!�����hKf��eP103�Tbvn�j��c:�Ҷ-���d?ĵ���O����k~�7�ĵkW���:�0 �(���%�U��<Y�>ڶ�m�eve�֨4���	�O��}R�OD~^��}f���$��߱�q%/��2�<�[tM�qt�iy��*�:�X���:89��)1�H�cz���`M")A�6e&�]T���c�ꀖ<Y�$�63s��1vFU��`L�}T�5���(]v$899�n*���&�?�V�K��GW]e>�������-��Kr�R;2�~����w�XD����K��`lD�fѴܾ9;����Ӈ<��#���8;��RYJD;K�36�Y����	�*)\)pvz̷��/X[[cT� ��>�)M�55)vLώ89="����x7�=�_�P�Đ��$�ȁT�8�rx|���w(]�����W ��wl���,s���>����$8mxZ�Հo��2(*(����kVE�/��e��tP���X
+E���&�W���˯���̋/����6�-9;;���qp����I���5&eE�,��@d<Z��J�F2.�g�Z��k�L�3�z��#J��l��[�M	�Ǣ��2c�Gi��*^)d̲��#,�g�L>OԋŅ@{(���R"�\�,sŒ�R�ݘ^�h��J�Ϥ���y��R��#�@�ۜY����;��R��,9�Н�\�09x�1,�K��u&� ����H�
LH=�C+��ω,-�͘��H�A���%���)�K�9��DY:�Q�Zg��h*v��	=
^TJ����>|xT��u�vۊF���*�u�֧}}g�!��إ&�i܅�3]�"�EU��}��2�މv9Xr����g���2u]g*�����Ψ�*�y����`cc����S���vy�X�s|R�d�<,�]�-%^Vu�T�da�ՠo��w�?ia�y(�B�陼�īuΪ�!E���v-ڕ����i��,������ѣ.�r�
]�]ؠ�uM�4� <�b��{������*V	��k9����*7�^ac\H4!g1|��NV��*"@� ����~�V�����������}�ٽ/b[�Vk�*9���В��[X<M�,    IDATsF��8�8:9������\����t���+	���f(m�L&�D���Vk�V9!�-��&�LP=�H��ZZ�*JRt��Ih#8F;B�X#9Ќ�A:0d z�$��>�(�)�����k[LPH�>h�{�M�u]c�f\U,���tX������2�N�J�����q��K�����R�i�6��s٦����g�ʾ\��\�C�h4b�^x��ۿ����Z>��>��0����՚�|���!ggg��_�%B�fQ�PJQ�%�;�=�2�s���>�	fYB�{�lV�]&]��(3��țݔ�L6��~c��>�U<k�D2FDHBO��k���s�/%���(T�	1�e����k=D����
�!�#��uuX��\-��1��91$߷�D|.�O���,��]:�Pʀ���S����fx�����x<^�������8 O0���!�{҇��@� an�B�����6ڇq]�ηm1_̪���ַ�_�㣟_�*��~�c��F�I��!�����cӎ��*A�.�S�똢B�`�M$��Bk�B���g��ʸ������.N�q��w1�G��2�89��sݱ������w��z��2��W��g&�	Mӡ�FG��:/�� 채�>�*�y���I���}Q,x�)�H�<�&�e1Bk�'�>0��:|�ΒR�M� ,�g�pq=�M�1�@Ȼ.���b�DT>y���Jڮ��c�J��H��q�1d��s�%�y����/�)���Oh�\�$?�{*�	���3l�bʒ�K4~����OL۠;ێzq��?x�޿���X�1�ٌ�b���,�3��poL� $O)�Γ�q}prF�����f�`R�"����R���0�Цb����^y�����^f<���#f������c�+0�X�P��Ԣ�`��k�$����-	�Ǩ�C�$�ypvL�E�WH��)���s4O�߫Y�լ����l (�X5��Hm�H�s��P:au���)��d ���\���Y��:��u���ɪ y@e����'_�Oi.�����Y@2��.n�FG+/���� ��~�dܿ0�TU@K��[�������5B?R�c�B�R ��M����W�,����{����Q��>���������Q_:,������Xl��q���{��f��L<�nnKt�IEI���Ǚ+-h)ʼ�w]ۗ\=�����lpzz�3�).���L�6���ec�2C>l�677���㥗^�W^a�ǜ||����CX���98Q�tI��ͥJSN0�-�1��Z�����欪*Du����r#�Y.����pơ�b��
EL�D�wC�pe�[��)&u�q��K��&0CP��h��%��r��N[�3'!O�S��F*��O����=ñ�y����uJ	����r$��$GW?ؤI�8�|��1�D���i��}�����ID�d{�e���$��j�\yC@ň��|�R҅V�`��U�k3�ו�pvz�N��֞NO��3ƚ�Y�g�y��=�'-�Jb�����Q�S}7o�L7o�q�ԋ��AI=�L�!	>D)G���$�8;��오 %�C�	H�����䄔�E͇wnspp�h4��8<:�J)��)u[c�S�~�m�����3�<�̦���1��!S��]x�J���jľ�.�a��ߗ變���!ڶe��.'�Ld�����i��6����Bz�=vy�_���b_��[�@�<��rP�:��@��.ι~�]>�{�G|������g>] �6��4�C%A;Ka,I11oj�6(k�AR�@��i&��gM���&v�7���T��d�aM�i��zA�,�E��(2�ue������Zj��&���������o���D�2c�$��z����R�$�p��h�$��gQQ��(ML�#���XC1Ҙh3x\G��^J!KH��AZd�hⱅaTd1���������)un�vy~��۶���ev�m����M���Ӵ�VU���ll��t:�����9��������UU1���2�N���9�������9���@Y�,[N���H/�;��$�C+�1M�\�T�5���!B*M�µQ*c�SPK��2�ѯm������,^9Ɠ�<{Ѵ` Y�b I��H���W��(�Z-�'�$b8ߘj�2�^�4EAY��ev�ϡ�+X�,�f��H�xR���������D�QHt�H�.�XIT�c��pI"�:�$&�5�P.��M������"�����J�$ҹ��l{29�R�#J�[��O�yL]gT��k/�S����w��(�V|S��1�&��t�]B��ipe)1&e�5�+2�8�Z�v���$@
W *���I֧�֖ʍ�WUf���(��o�������}�Y������1fyc����KA�%-�U��0ПTz~��-�N���?��؞Y�rY.w�s��A�H.�̯�S��L������3��"�i��\��dw�����9>�������T� a������os|4�t�;�����A�+U�Y�͢fT�\3�k2+�B��tG�����A��L�ߚ� )0��Ѩd2{Weצ}���C�/K�1��.w��)�jV��ṡ=}�XeI�u9�c�J�.�B�&I��8kp���U~l,�p�a��jC<�u�"^Z�}X�v>g���j��	j��E�l���A,ZU1��Ç�<�LC��UÆ��nX�{X�>�~���i�~��KU�O
���Cw</m /�_��|��5�ס|<ظu]���׷7��Tw�&W����&M�pxr�$R����3��E��mhЩn�&H@�E�yO*�ULA^�R8OzĔ(�k��Q)bL(ՓP�!��+Eˊ�P����}�ߺ��A�֚�u9�3�a��ƈR�IU]���ka^g����>j֞a��r=��X[,��(���\��g��\�UP���(P:o���m�d$%�E`:�+�-F㔱>�wI"��PS��Ux���N��Y�1Z�L�ԑ��Q�BJ���4����8c�c���AQUGhӖV����%^�w�o׋B��>�%��hL|ԺU��wQ��s������w�?zp��Ͽʯ��o1�w�fZ�I%Q"����.0.
�Γ��gKfuM)��x�h4BiǼi�ǜ�f��_���)W�^�C�tX�2�vri������3}���Cv�I��1���l��/(�vZ�#(�9��~�kb̯�:I��)u]/�1�=���ǘf�%����K�x��jИ��^��������&��[���g-��Z���K�so��]We�����9��BYE�	c���	�g� �b�T����U�� ���F��>upp�|:є�q��с�DY[ۦ���Jn�f۽m���U��O�\���KV�gi&���� ��v66؜\gws����̆���}Y�˟aR_��2*�Dl��i�(�
�
RR�ń���L�
5Ei�!��g�[�vX]������{�?⭷�����dz{�4d��11��$,�?��w���\�/��Ļ�T�6�K՜���0����d�����bY^�_��<�y�2��:㇇
� ���0�/�����z��l�9����|~ڟgp�4I:�Wh�PJch��}3� _�����:��F�eY�)8�L笣g�d��2�A�F����g��� )S$a��$�r�f�-�%8Pl��QYĺig�^҅�PBt��b����F��8|����eц�ۈh��s	9j��eU5��<r�RI�F"��)��ژ�� $k�Kb�(ZDy�@C��AsY��A:��� !�4e�C�uRZ5��F?&Q *����t�Gڮ��,�WZO��b�>��?9>Y�����uk2�|tvv�nݺ��������o|#Z�tA�mT��:ejچv��Ç|�{�t��ʫ_E����5zM¡mB�'��l~F�8g�eMΜ ���{��Xf���&J)n߾͇~����:��e�(1�zͥ 	gt�>擤/��S����o���v�)KCJ��K�=�G�L�ǘ�a�{"�Tp�s�]�y�
/��I��j[�S��˙B�;��h���N���1>Y���T����J	Lv�2���+3OR�j�h4b>]d����&�H[wh���V�R��O��:66��~�W�\��m�J�A�Z�lIQ�K��#?��yd�(����]�|:#t�|�����*D�Y ��(�}>�W�y�2T�o���W��	:o������.���U~��x��u�no���Q�rR_��iU�a�,��/7��F(m���^�'�6�����A��e�ch���܋/PM*O�xx�0c1����z�]�k�r��t��_���փ�k�Xt��@�B�y����[Y��*���`p�?�[x��o����:�Z��1�u��Ou��lvJ�4KG��k������nBX�Ƙ�n��huf5��:�?SBʏ��X�eV|r�tV/��j�`�!f۽\I�Rk"BL:����%9��1\3Q8+h��&��ߡ$W(4]3mU	Y1YD+���0�(�E��*�yH!%���䌨:�&���耊1�d�$��1��Je�B�Ť6�W���c�7�R�Q�R?�H��� ")v1�n4��z�4I$ň�DItZ���Q�F���gWRRJ�N9R�)�@�:��EQ�RJ�`��6`���F1���c!Y���=|l�����R,�v][We�������#�M��������NO�)���͛	mۦ(ʏM<⵱�j���x||h�|�Mv��g����]��DaQ�����ʢ�����|��tF�����(f����e�w�L�X,|����w�_���q!K�m��檧��Rͽ��0{x4-���'v=��cT?��ˌ������w�mH�L���������K\��1/�D��'�<�W�.�Q.g
����Z^�y{��Y��N_q���1�Q=z���&k#�ɓmU�h����d'�p�j4bwg���M���I1b�e{k�kׯsew7{��`|��{i�~F���ǿ�5=z�3�6�еs�����C�y�������>�ڞߣ%�xe�	)���|�?��b� ���3}	MJ�-*����+_�*���*���6��u7$\,���q��φ�M1�2�"�{HP7�B�P~��ӏ���@��w�;Ϛ���=�}�y��w���RYn�e�>��>�|?G0��U��g��n.��9��Ԭ�hV�g�˺��dyNC�ou޽,[�j��Im�����ܝ5/݅���������_���)C}:NNN�������l�����X�0Z���Y���|���6%"!%��m��`��$%ڈ��5L2F%AG笏	�V��*{�)QP-� ���Et�f�����[��$*DD�GR��9E�,E�����:�R-�)Af�譈?NAG�t��L
!:e;�z�/Ԧ��h�{�:01F�I@2�e�Jr��Z�C,�1��ڤ�s1�co�E
��>����AW�R�q�I:oA�l�K2��Ҵ�b1��8U��Fb�֒��|�:b8DB�	�ċ�6�I*��T$�BE��`SLN}*��[��	":F��Rڥ�x\� �t��!��HL2���M�
��Sw�y������w��6��|��.����.�m��|h�G&���j��*�M��|t�6��o�M�s/|���7pE��]h�� ��X���1�o���Gw	ƕ�MM�;�r��ƣ��w��?������׹u�V�yBJ�΢�.�!�C���K$g&��T��x��d��^\�.���Up�jau��9�d0�l.w�������W'�U��LG���]�Ւ>N�>wFY�N�>S���/�X���rPk2Á�#m]s���x�}�]�P=�E�ޕ�dbFR0*J6��xv��n쳳�E<"���2��I/oQ��^��!@%�U\�v���u
��8���7x����[ob]����V���=���f4������c��Q�K�~��xOkB���#�׷��ڥ(3S�	-�"����Ĥ�*���9�yՒqh�Pt�'&ͨ1M��UD��ʡ�%r����MP��Y��)K����mP��t$��-�t�� �3<����'a�T�!����WH�l�;��Zz����������w��t�z�u�����r�
���<��KH�q�����ѣGܿ���q�-���$�]�-�"aHQ0�����^}6h!6�	��]�6�4���?-���v�)tSRH�ke��Ց4Ac�$ʞ�������"�nH�KI�Z�H����`;���`;��N����L�T�E<�v�B�Z��C����͛7;��7o����������YF3�R�r�L�Ke��t�m�Z���}-B�)�I��6Q�eT2R*�]J�������_��$c��H4��N��N�C��%%��(����T���1XM, M2�A)���D�26D	$/1��$m�^Bx��,=�����VX�'�R�(U)cJ��	�^D��C�����(�]�`'6�-@��zܾ��k�֭[�d2�����3}G����6v�S��o$ԕ�	�4m[�빤������������7��ۿ�;���L��P"XWr��>���ͭ[���{[R6���zu����$�s|�]�r���-r�>��7}��;�Y�~�����|C�u�f3���@�x�JXH��f��]N(�I��30}VŘ��1����񒲿X,��j��
�]=��.����0�(Q�}1�r��c�Zf����s�RFH(��җ0�����6�@�iY�0��[��g��W��E��#���l�<VVWJ-˙Z.�U����^�!0�1�
$v�l��W�L5��|����>�U�{'���ccc���X�M�_.�>1���-3n}C���w��7�蒔�.%*m)ʒ��9M�,eo��ˀ�+�,)1�ϗ:��"c�����ym�����F�|^x>f6�q:=#�fm}���/pew��x��rL�\JʘMG�.�*c�zŇ���/���6Ta�F�
�x���Pn,ن�v �V\>k%d��֋Ռ_J��O�I/��h���s���>�^�h�y�l~��"�*
Wa�Ba(&%����`}�J}�O���ƍ�!&�x��G��sաq������x�"g)t-:"�4��3��d�>�L i�L
t
AGҺ�`Bd+A����I	�(I��1�h|��jQ>h���n��u1.?H]���k�(#���o�{���{?=��o�M;��IXخ1�ģ��Ye۶momS��OZ�N�k����h�8��W�0A�^��A���(���l�>�N���D�2�����$��BҺ��!im,ؔ�7J�����	ګ:�dt��+���""��:"��d�j�H�jD�����dc=��1�%�-7���a����0����<�G��>����۶���h#���;j6�����GGGR������|����g�͛7���3}��ݓ��BPb��]l�J����b���,f���G�l~Ʒ����s�/��2/��_��Wi������_~������t�h��u%m�b$��'�����#&�k4u�n?��_������]<x���d�`:�����l6G�Q5���O��Z>0=U<��[,�e�b�^<	�
�&bub(˒�|����d�s���A�o8�����R�X��놅�9G�$٢��	i����%��i�[c�f�R�=(��m�msV�y�-��tߧ�WK�O��i��ӊ�|�5��|�<�sד�k�
��8g�b�ʒ���Zm��l�0�,�:fӆ{\�,���(HQ�7-՚�Yٽ~b�(
�
�vL��''��*~����u&�1g�9��#�lsT7�u5���=��v�$�,	m̦�*�G�N���V��C����e;D��"!$f���`s{��G��;x�w�}���m�4UU�������b����a!lb��Y�k�5���3{:y��9=;�l6���
�_���wx��W����_Ѕ����[lo��}�m<�zE�hpnDJR@T��������S����.�~��=F����2v�r��c�\��kw�A�]n��q�u�1��ʰQY,�ι�Fί��z�j����������3�O(�x����׾�˯�o�q�۷?���^0����sm��    IDAT��Õ5�*{�lf������Y���U���xD�^�a4YG%�(�����t*v�(U8�.�+��קg���zWD�[ԋ��h�����uR��E�I	-J�I��:�3��%CM��E"mЁS�T��̕R��:��i�ME����	�ES�H�֝E[�u�Q:c��C�����d�>�w��ƍ��t ���tW�Wڣ��SE�(ڮR�.��Sl�N��F�I��騬�$�7:��ѕe�&���]���@Yy��EQ(����Z�ԳL&�|�?����1��R:�=R���c[��h�(^=�1e[����.�2�m�˿.���՗�y-�z���y�f��?��{��{I)�I��^�"���o��7oݼyS_�~]'�nݒ��뢔:�_�D��g
�nܸ!'''҅YD���6F-�Hl}}ipP�Řӳc~��-=zȽ�w��	���r<��v	�C����� ������g8UKf`�u��o�{�23��/C��U����Ռӻ�1 ᓹ0����m�Ռ�j���`�z;�2�0��`��kX����g���y��rPt�=��)�l�_f�rИ����8������m-:���rlݓXW�9��FL&Fe�f�_�LҮR�eT���Ễ�Z����Y�(���p#p���!��5�D�Q^~�+���qmo'��R��jD�\^�,����Υ���*����瓼J}ILe�Ӱ�J�
�\A�f3�Óc�z�-�����0�N�ЃA����,��Z�2�K�
?ϙS�h���"u3�mj�7�4�C�tݜ�4G'3NN�\����~YS����[;lnoѶ_�%���i2�{P��E��T&(��ڹ�PyY-��*\�/�jyx��q��Bsf�Y�c�7�{{{���s��RJ����0���e��5�}�Y67�������N3=�sp���GG�����M�)���r��m:�2��u�s)�(�N�ֺA̩��$/]D�7m7&�p>��a�����]���C�d:%�XGm�B֊�l������(������H��;���1&km�˔�6fjִf2��Η� �@g��Y�gG7n�P����������ɭ�o��o~]�c��y-���O����h����qP����p�{o�븷�'��$����w��ٸ���' �׮��\����]������g��6����n"J)�7�P���������͛7?���)�X,���RlD'%)���(���$�o�D��}ĝ���޻o�������8�k��Qe�ۚE�bBi���v.?Q&g���
���{w�����RD[CL1냹jI�0.{��<!�A��qy�_� ��eЗ�;�hm�'�:R�e9�^�����~�iJ	���P����.g!WI*���I�ße[e���U �OlI=����+�(H0��'y���Y/��'��y���]}���V_Z�,�٢��8WR�2k�T�ƣ5l��7��D1�1QY��l]�!�^�[����9>��Y	���H)��_��:��rA�S�.����1]����J���~�o��ݻ?�������V�uF�k�;�`�B�\��|����<�Α��iO1�a�1(�����^f:��d��o0�����C9�I�h���E��mO�k��0�\� �ɛ)�Կ,�b��[�E]%nmu��Z�}��.��������[UU���q��5ڶ�?�w>� c�Q�+ƌ�&��g�n��3���w�srv���U���_���g���Z2���G���T�k��{�#��]�1��^z1��W>%E���
>mt!mn͛��jT�%��֣���6<x�+��N�y��jp�IT�Ϸ�op��?�� �������F׫�t}U�8;;���}�5d�>Y �)��g?�����7�xC2�J$��Q֤�bL�ֽ�M���1*K�QI�����p����[뛘�Q�����9;�*�0��l��*�NO	OY�Q�}̥7��!P���|��P�a���<z4������� J�����뙩)Y�W�=&*e�-ԋ����A�!?o��-�x�ؗ���x�s!C�	�P${2�~`�e�J�(҅�����h���^ �|�sQJaz�R*gy���������-Ύ�LOg�U_��nllQU!>��$^�#���\��*C&���4+��
1�",�b<-�i���RZ`:mx��i[��<IV�|���2�'rn��9��z�ؕ�>E
��(ʲ�p���<zt�ՀQ��DSX��sy��(����O�*RRH(�}�3P�&��FkGaRL�$c�E:i�@Y8��z�O�l.K��-�ۜ��E�{����AJ��b���1[��e\Ul�:�O�sl�@��d}ס5M�o|,���lll���ѣG|����3d:������!�����uR�|�+����a1Ei���C����޻��7�}���3f�:ox1�6�c�(KYU��UaݾR$��6!��� q3i�̨��iqf�']�����a��n�͛���-�߻�JYU� ���w����g��q|LpN��"u&�h�
� �����h*�-ZB0β��F�����@�+�J��q.��*�J)NN�X+6pz��-�T'''(�;v�#m�E���O����2鳢Ö%zE��w���%� ���)��y����TB���%&��5A]��w��%>�]��]~n�g�L&�e�R��%i���l/L`O._|���P���"*�%Ԝ��F�<HްVe�h4¹\�H�H�@MR`KK5���� 
��r�o��\�g<8;ʾ�"�q���5�5-Bbzr�b!�Mã���[o����%������tn쾴��S.g�SʎO"�|^m��}��^�AeW�k|hP��h�$!� ��e�TE���d}}�Q�G<XMu]G#]�)��͜z��ʻ�esͱh:��
0��Jh�Qo]��nyl�5�:��>����E�{�d��?����8;;���l�m09����{�fY��L�Y.3�m{,<")I�I���g�{f�4?�����1׼��ŌbbB���H-��I��-�f��X�UY�l�� "���Q��ff-��{�w�I]׉&�U����7y]����#�ׯ�tp�.���>�p����c}��tzH��3�N\�e���C�ܹ����{�pzzLU5vGتi��`�A�H���hă�cbJ�G�x^!�Q��NC��EuX����Q���?�<
�|j@��NB�a}t���ѻ}����|�HS�	O�ƤU<1ZF3�/Q�����R���x<N�u�\I ;m��9��Ϭ�两�\������,����O���R�g�.Fp�c)�/ט>����jR)�(O�վ�h����%ދ%g�� �]خt���:o]�i�T&�d�£���v�.����'�ː����^`�Y�]Ӭ��Nd�MSqr�`Mz:f���;�(
��1{{{���S�z�xx\S5�`��+��ٙ�a��,K�����O��_��=�Ō�}���)���%BF��P��o�nS���$t�o�\)E����8�`]IU� F��A,Fl�vM����ʵ��'�le2�"g4����d42�QB���89z���}�R�p:]a�!4���\K����I�_�1���2�ߺX��?�?��:�,ĨX.�<x��g�]gT\[$w��2�֮!0�5��)[.���ײ�i�֐��4~-�������,������l���	�gS�k�Z(��kCʸ��2]�MK��v5&�8�PRJ��PR*/|�Jeh\���'d9�9͏�<���N���!�\2��9+���-uJ�k�����yCp.�]��191��X�d�\�Z;�L��%��9�Ʉ�d�JFy� ��j��I�n�8��5z��)K���6 ��������^b\��&��D�&Zǣ��me�mj��-�|li�2�I������j�|�Iܔ�~�Y����}��q&#D�!��uBЈ)˒���Ez�
()	�1_M1�0�p��^�����:�@�gU/899����_���H����P�9�k�9Ҍ�ӓc�}�!}�!W���h"����2��dNc�o���~��~E�����g.�\��nb��`��x_�l��p6)�Ȩ�J�ɜ����	�W�GH�qu��!j�`<Bg�|o��d���=2c��s�w�p���rNc+�/h�ckAA1!�;�kZ
�wTU���@���[�D�x��:~� <���a'y���$��Ln֊���u�8:�������J�RJV����L�S�s\�zm������'(m8=�rt|B�8�T\��E�L�g��2�� �Hcc�Z��I�=�Y�j���*�R"e!6RHʀ+�@�΅:��%��zj�Ş��;::{{{ ���T	�*��2� B�	`�~�i�7�c8̑��r5c6=C�W�itk-�'5
�R�}U6���a����畗^�,K�?}p{-q��i�t�۬�I�M�ԙ�ni�;s/:}��]��8����1]V��j�M:�"2*NϷ������$��R
緛5:G����OB�O�������N�O�=���c ����ϑD�b>�SU�)��i�b���LF���|�;o��oP�%���ܽ{����/eN�S����#v&;g�������G(�2����lN�in\����1�q�n������'6�9�_:���L�����8�D�J� �)ڌ�a���8� Z(23`r�͛7�Z3�B0�s�sh�s�{��x��!�������x0����hA�I�$!Hf=߈��Ĺ��ŝ��S��~�ƹN~l#���]]� a~7JJ}�Skm
$~��}~]���hKʉb00�毢(BqrrB�0f�d�f�u#���!�̉A`��65B2��,M���R���qȤ���h!�*�#evp�ɫ�<���yjP��ʻeB;'c��e,Px6Da��%�w�P��L�}�&ZJ�U�'�%:�R�I<���Q�3�_2���]�>�`4住�嬪�=|-��6)cb]D�ClB�'��rI=O�����
���T����đ����k�pEA��5�sG��F�v$��ш���ш�j{>�Q��Ӻ�h�}� T��ު�X*�x����g,�(4Ҥc�
z]�k���ڲ��l��?�l�IEuQ!Q�(-p? 8�My8;c�sA=A@f4�ȢT�N����⫯����{&�n�w��#n���g:;ag8�����OFL�ƃ\K�.�$�!2���|z��l���c�,c|x�Ji�޹˭[���ڿƠ	T�$zEt��j�z����mÑ��T����!��L�a!*�9D��	/(�%�@
lA\�`�O,��rF��x�9?�1�FL&4�������r� %���&3C���hF<c�L‸X1/�I���,�r�w�s>K�hw���H2r)p�$���# �V��H,�� �D�$b@����}ָ�3�!S��@��Q;Bw��5���0���|�n{�!���$�bIPK�h�*�W�*g�<#�y1g:}H�^چ|�SN�����BtT���e�(��b�S[O�
e
�R�& �%�Q!��3Bt�:˩}���=_��tӃ�(���dY����D$���HU6��n�7&j!ڦ��$8�ɵ�6KBY1���<�ލ��[����-�Yt6 �o��&�I����q�h������ ���"�k����f3vw��9��)�$(R@���]`��3�ZQ�"8�$Ǧ�J�DV�Sޛ�L&��^F�U������ů�����6j<��퉝>S��j�@	UAH��&��QV8��*z�7 �l�	y!"o��C���minUUF#ƣ=�v��ptt��cM/��nӤj���\&� �H��������~��G����˲�����k;��.��W1������$v�4������Ͼ����7r|�z!������CU�h�g��Wi�o����ۿ`>�!�g0�����,�GX.��eI�u����h{��t<��5�����y���W�\9`�J?�֯�K�])������֦_L�9Q��4�"]M��ԡahr�a��8W�G�4�lg�f��{���U�9���W%���e�bV/@�)vwǘ�yd�ne��@������< ��Z��)��5���p.zdLk�T�kc�U��/�kO�5y.@i��8"F$�t�<�2jv�;�U��p���b"�il�ZЙA��R�Ň���<O��>&̥1
$R�q"uR��ֳjV4!$�J-1m�'Ĉ�ms\�ԫ�S�YZ/BXBk�R���;�p1��λ���y�|�XϷ���l'�"��2\�e�/V}��ٛ�s�9��9���l��Fu{G����kmn)H�TQI�P4v���{��2��T*SR���u=�|�X��ƞ��{���ѻ�
#Dp��"�=+df�RB����E1�v��G�m�VӀ�bU���!5e�%�.K6�N9=�1�9`<9��uP�����-�K��[N?h1֦ITV˶SJ�G�G'R���1�;�q�Y�&h"���7h�Q���d��o�
ߑ(7M���ҿ~����E�b+wU��e �/��ߙ�����r	@����C��������c��1�6Y��9?}@9��*��\[/��s��"u�M����s�!0���4qgH 2�s�R͖�'D���;�sX?����孺��;��!���!�#���_� U@�
�'R��Uę��<n$�c�ݣ#~��[��V�ـ��T�"g.T��̝qڜ����n����oeZK"�y��-HŰ0H�	Uē:���⃇�2�)��C�����*b���$%�%F*D`A8I��Z�:^U!p���T��(0*���A��o-R�����c�Xy�SW{�]&�<��B"L�.Fh��<;OA/��L4(�Ur�$'ELNgHN>���1�!��svww���[+]����0�۶%�W��3���4'�1���>��#�=���N�&q^J�W�\a>�o�/Z�p�{�/�n���: ��ɘ�k!�1D���պ�
̞`�>�/�=Y���M���>�D�;D����2u�n�)SYJ�&L7n����:�"DWR������J.g�3�=<b��u����Өk׸����f���n�2��D*R���.�B\�~m�bv�q�C"�l�1�7�C��2Y�l��Ď3*�G:GNF�e��+�/2���:c}��kj1Fc� F���>��s��l�[)�@lȆH]-)�!�������=�����L�����{Ì�ܠ��0��鮵�婔!"�\s�3"��ݻ�99:�D�o<��ݖ�$�V]�b�h��k��󰋍6�c�����XD�P9�,�RhS�3�E�+3z�`0�Xc��ݵ|��?e�w�����7<<=&�$��S�{9���fF�*qN2f�������4n;\�w�,Ө,G��sM���yQ���GȈ1)�Y�{�Uĕ�L*���E�"ϱNPVZ�LF�lE]O1�K�RI�\L�EA`����
�R8�q.2�r������n�geK\��ZVh�8�z����gܼz����h�T�� ��#�B��1zD���3�߿���C�޽�r�Ļ�]����k���w�L�h�c4�`�?���>����E"��ߵ��گ�\����;���;==�z���A����
��ړ:��F���� |BHC@��b�O9|�ڗԞ��;�ʙp��Ѝ��P"8?�2�w>F�4V�V˖\�я�pg��S�?@*[ "!RElH���p�������egw��xD8:��kB' :�#�Τ���z���э�bf�_n��>�OLj�2e:޸@rchg^��2��B7�;������4Z��t^��\!e���n��2��{�H��Oc����6*+��	�Z�-8���9<<\ӽ�"�h!�D"AK�̥E�ͺ���+MUr�{����!?�J���{RiI��*k����R��������(�!�UJ!�GI�w���`2��4(��%"8p�ipq��5Ŏ 7�|�
_�����GGxp���3]���?����P�cM�H��=�    IDAT���n�xE�Tq�o���ɇ�̻�-�Œ�p̍Wy饗�FL&��4W�V�")Y����C~��=��KY@�^�C �A#<s�Y���H5���6����bIm�i͔R��L��2a���|��_z�o|�ufƭ�>��_���B�(W������[���;��<����
�Uհ�b�m]�3��Ղ���srr�·=����C����5��m!�5�2�w0���N�[�_�H��wN�Ex��&\�)�J��ck,nd>����I�N��.�~�����w|!v�����	t�&:tBB�T�A�����}j{bL��	�BB�2	SB�]#��!Ɣzvn��]��!�=e'�.Z��$�R�0��Y��g=<e��&�`��h̕+W�}�>ժ���,Z�.�D��k�U:�ۍ��e��Ob]���m�#l�`�d�Z����u����T�.�-��w�w?��]�:%�v������וտ��9��Z�X/��k�s�fZ����~5u�VU�b���Wc14H��_t���!il�Ķ�Je%dj`�W�~�:M���w�t:%��r�D�D��[R�.�'�6I��TyW���D@(�(�D��A�;��˯��3�p��!7���rq� W��8?=����4u��+�1�����������sL���e��Q���[�r�`�Y�)_���>�xƭ�������M�1�eXBT!q>�\U�u�x<��7�ÿz����⋘�%ϳ͜��� ����|�o�zĭwn��G�����`4d�J�@��������J/8:����ý{�x��!�yb[�PR&�h�B�и �������o�g��n�,���)�����#������_{�[��_A�@��� �4HA��פ��5:ӌT��9�{W0ِ��-Q
N>�ڲmj��`	�!Q\TU�^_�u�v�����ԕ�ښo}�oB�]��l=�W�9�R�u����-�-��sP�ր֤L�חL�U@MgS���2�H��1z���O1t�ڗ؞��[,�x�J�[�d�B���E7�ʄ��.�'b��%��s0���	���$i�Ve����墂��b4���g��}��%�ѐHj��Z���i#X�kZMδ�zo[I��2��i��Mꮬ�N������m�GR���jM �9|��u?myW���c���x���,��z���1�����S��;�Lf���z���1Bi�ƒy����P��%X�6��hLQ(!	�b���Eƈ��$(J��:�s�������k�ٌ��QK����r����߈����Fӧ��z�I�� ���_��^c�`���r5%�$":�w��SN�ψ.�O�|��-��w8<�x������7i���${�=�����0��x���woS�#E�ɖ�����<��g1e�����7���7��������?�:�u2"�@L�m!�i�L6��3Wy��7y��78ؿ��ܾ�6 *R6�*�����+<��WPz���Y��o�M���3�F��V
��6D!�A u�x�
Wo�ȵg_�@����F#��(oȲ���.��(r_���HzM����AʰY穛����:��/�3�"x�ώ�!bׄ���s�O��W�Xc��*��u��sY�o��]pĺ�#�D�}~w���n��7:���,�(����6@�؎A@(ك�D�w"����E�#j|X���a���G�S�C�'��9��P!(1�{�BJ����#{��׷6��ðvH:G��,"H�ሽ�k#\ erbh(˄1��6��nk�\v���LW��ȑ�#�-5u�nFD��EI��庝e���e�ēX�p�6jO���ڈsv��KY�����A8}�sk�{��*�n�O1�I�g8פF�Lᚤk}��+B ����x�͂I��A`2��/8�M�5�
��(�:�mf����HH:�&�_��8�5f6l��TЄvSsM$7��!���䭂�PJs��*�kN�Θ�N�Ww�yx�Ã�P�h����jQ��FF�_�kO#�EI��:{�Ƀ/��c��9�����������?��]��������8�B��H�(����X�\A��������A���w?��)v)kO�z8$O�"wv��wߢiQUMҝ���f�NNg
Q���� /2��9Z)�,#xP�h8�ȇX/�JB�$U.�w<�l1�G�lW ��mCŀA> x�=8�瞧\Έ��*�*P6�c���e�J%]�G��5���y�����.VQ��6�0m�O�܇�tkS��^�\(����1Ɣi������3�jB�!��R3��-R̤���<���?�?��O���+�R���e���4������j�r�RZ'-�NU�&�~��&V@ˎ=U�\���v�%A$��PIZ�5�����&+��; �8���2M��ʵN�G��n5{/k��;�}��s��Ɋ�H����}j"I�ä�a�j��!��/�[���b�.Cv1&N�~)�"�;�����6e\�"����Ν;��x��g���4���3�s���>�T.�]�wL����>���������>$)ѕN<B��nQ$�b������Ae)�!Yw�^�ʲ��:3�ImBH��&�� ��wB Ed^V�,'8:;�t6�iB$���b��p���$�k�Z��{O��Ɣ����-o}VB�;ɻ��I�`�eX<&����ٔ�����6��}Ϋ�(�d����>É9 3a�г{�%n޼��sh��46�E�x��`1���ѝ{���_��1]���`=VW�y��}�`�[/+��z~������-��9�7<����o�����v
$�dgr����)�,/�^0_�P&������cr��U�`r������hYq6]@��@�Vx-��N�.Ғ�w��y>����旿�%y������b�Kդl���.�:���k7��9�iq�����x�`�Z2��������֞w���_�;���]VuEVYFӤ�%�b<�p��Unܸ�����կ���Ͻ�p�qxe�����V3�R8�BT.dĻ�;��:5~�!]�֮)�֙�6��>im�@�{ t�C���u��.��e�������>Qs�9�:\��{C?�fah��HL�*�t,]0�g�iD�"6um
�����j�T0��� O��?{"��j]�s9Ep>z��QH��A����8��(�E�ڢh�l�ƝgKf�����}�$ӻL&�����,�+�!�QjHJ�z۪2�-�s�Zo��.ӷ���8]SDb��Қ̨��iA�En1b��`P�)q�rBQ�F��d���j�X�i_҆u��7�R&���p�^��uv/e(?^r��e}m���؏����?����M��M]˛n�� ���qHi���̴�w*�����[7�w#D�m`�/u�$���rU����w��9�fMC����v�I)%Zl�Mg���i��������CJI�$AIVJb��2���i�����F`C�ɑ\�Nvp%ӳ�Um��$b�sD�L����Ղ(���,�*GsAm��d�g��R����?{�-��ʟ��C����O�ۿ�[>8���4IUF	B��w�ի׹�ʳ���<{�r1D�{�7�{��^x��_���&F�C��@��!#�)��y�y�կs���64��,8��dʉ�(����'/,1��u(��)��[������W����LN������D;2�Ny���w��ZK����x�eȇ#�!"����g'�������q{m�,ؿ��}E����Y��,�J
��w]�����C$:����������b n�5�������i��-���C�R�*�-�K����#�'o�^�h*�(D\;-���!D���@�x9��B����_�1�D$�@���℻YN���s|������������x�x��;M]R�UXwe���EX�Iڟ��c]��=ן�J)��J
�4dENn2|41R55��$J H����qC�9}��uqx�����9��x�~�:�Ɉ,�Ę�SG�/m\� �>��!��E�>ٹwc��ߕ����9��f��
��0�nC�%�<C�5���q�u�y��y����"����J����j[�^g�c��GR�����Š���\F��T���L�04,WV����5���3�v���!r�`MRJ������Tu@G�S(C��b`~��;��z��.y� �5|>�˧����\�k��&�n<��|ͽ{�����G�߿�(˚�jh|R�@hL> ��q����u���%7���}��p���ܸ�?{� ���{���)�]�j��g^���9w���W���4h-[8�!D��Q&.��(��Ӗ?/�_^V����_��=|�6�|�@��B�3CD��<�V��lJD'꫱���L��A��~�<��V��.�-�'��n�e�,x��]t�.�/��J�����k������[��o�ɤDH%���k��я~�T��Ȟ�髚+"��EAĐ��ZA
�]Kbk�[��µD���'k!"	�sOF���h��s�j�o�x�����s��Y,KWS�U�4U"�\��&�`��,C)�`4m��M�[4�z�i�n$}�ņ�9l]3�(�K�LF#�Z,�d4�v�ȱ�>6M�&�����E�q���9����}�\��0� �+������r�.R�\�*u�_��u���c}'���k+w���%�&�� S��V���µgO\g
A���L��A���(|�px_�뚥�(�ϧ��۬�vA`g����}(A�w�g��甍�llt��Ѐ4�)(��;=!,O8��M�h�9���wyNe�H���+�-.�Qx�8Z�yx^��Ś,����p����C��`�f�l��L��QJ�1%	���J~����7��_3;?&�
�cq�������d~6���y����׾J�<����89:N�6F|��4D�� ���T�^|�?���y��w��f8QV�$�%E9-�xޖ��ylD�{D��Q��*lY��d4��j���$H�9R�hr��8�s�΂I�S��9������H��ҙ����i������]�8v��u�����u��e𕋙�K_�A�bh)�D� �U��Z
IPR
���R*ɤЯya��˿��ŏ��/7U�S���)2}AHQ�c�QDA�!D�Iʑkl���^k�u�.()pw�12E5K���)����W���=�����n�\`/EaA`L�p(�~�()l:e/frB�(�����s(18��&�w!A&�#%"�V��i��(@K��
-����[,TU�sn-�V׏�jO�uYî��{鵍��Ŏ��ǡ����vI�r����u��~8��l��A�ׄdj�%�Y�]I�����I�Q��J�nJ��9���!�+V��Ya�%מ���4͚���%�si@�yY?{��w��(|ʸD��5e�����^�
����3:[�%�����ūe
\+�pT�(}��5�l�K4�[�0�K�ǣ��h7�S&��^�M6��	��g��������;w�cw�">�4M���Q�&7�����;_Q���������q<����z#Ā

�2DTT�����,=�p��n0��?��?}����6�H#��k�TD�Jj1�ֱ􉛲�4��M]!�G�$/3F��B������f�'b�� IXJMҠ��B>���|k�ɞcwO�џ<Hl;�k-��!`]�K���8:�ʶ�ww��n�����\Ƙ�|b���wY�.����(��h�
�C����S��̞h�ԶNٽ�VQ pi�ƶ'���=w�9^��:\����������[bg)�"��>~x��x�`�q��3�	��ٛש��:[2�mCpĹM'U�	�w��~�i�JY�N��{]7QzD��:ӧ�a4`�%�e4��,	��(������lFh9�V�!F�њ�>���:���bЋ�z@�$�-��n�J�� ���i}��Q�sS����uI><Ew�!D��0��q5Fzr�6�P/��S��/"MU�Ɗ�1�>��V����od-^ꕧZ.��\�ju��ޢ��6�,�kb�����TW�o,%O�e���d����>68۰�M�e�29>"d�!�Т9<G�S��y�:�gXh�sc4�h7Y��������]>��`A��DR5�5��p��-�L �%Kp��^$�d���AX0;u����
�
��b��IE�"������� ͐ݽ]�S��3&;{|������]�y��N%T��T
h$G&'�L�J�J	�J�F�Nv\�W-�MIaB8P�Lf������9�k���C�ȇ,�%��]�Ԟǁ��NT�v��>V����`�7Y��z��3��ه]t�c�;�n]�	��˪�� �����-���)cZ먢���XU�(%kQ6'O:n�ڗ۞8� ��1FA$��)7'.����.?�%Ȕ�=�{�=Q�I�	1�K��6C(����ŭ�����7��7��1���ӣ����`�)Z���
����t�����u�|� ppp��k�о��r�!�ј���6�u�b6Gg�"��;�gw��Yܻ���(�+>:�s��ݵ�v��ԕ�����l�'�.K�}�sc����MRlH@?/뎫���/�eY~,��]VnY�V�.���w�^bDӠ�F��5��d@�2�����`?�1�����Y�is�H&�d³
5"�(,Z��=�b�=���qk�ZC�L����������ن�G�޲'��{�#±ZN�)��J&٘���E	�Ai�򎲶(Q0P���t��Zy���<{�G�;?y�����ǈ��/:�oU-��U���܀�+f�#�� �BD� n��,�MI�a�*,��*�d#��l*�
0BcИ�V+8*ϸs�.Y�QN ��s���}�޹�u E$3���[�wIV�%��.���k�R�&`P"�D�u�k��',�g)��=��2�C�6�(�H�R�,Ǟ{��(i��~l#G?��R��ہn��w�)]0��襱����w�)���|�� :�����]2�;�~��e�_ �n� :8q��&�gY"�њLD��VRZP�������~����O5��ڗʞ��T �S!2��ǰp]��9"@�D�Dۇl1S��6JK�.Q���j������*��_��W�
��3N����}����M�HZ��v��|�����Xmuõk�x���y�7�˓F��������c��%�n����#Ƥ��̍���_��Պ��������5�=�u]�컒rw�Qv<r�.d�>.��4��uY��(1���,�,��yX��e$��!��<Ϲ��Vg��9?Ƅ���1��Q�\;U[�shR���cd``!B�ȭ`��ߪT�Z��uR�h���!��A
��
-FC�IFÌ<�,����Yׁ:�[�����w-�sY?�ݧ�cAGr#�(�@+�tA)�'��I��̀I6b'+0Ab��AU	4o��!�E��C�%=7n� V�z��v�l�ݻ����v�"��[����/؝I� ��[[�����,D��� :3� ��(��ِ���ͦ�|!<�Gx��c+�O��g�����W_������������Z˝���|��I��u�ٽ��#�_A�֝�B�~���`$����2Fv&c|ԞԨ�<QD�V(�m�4!9��e��)v�'[��ܔw�������=w���q�6�J�-��u]?R����9u}E���("��>����Һ�r�J�bBD�1AX���ڷ~��|�G�	p��/|j_z�T��Jʳ��� �XDi�@o1(��l���2s1�25��o��h�n�pas��	�T�W�����~x��O��w��htH����]BsnJ��|�(��e�p�A��FG�"h�Ŝ�#j&X7��,����������c:9Z���j��ko�91X~�_���Q��|t��[�'�L�.{{���M>8�aS�L��`4(�Rt-k}�6_�R=z7���"��Is�����F��E�923    IDAT��a��}"S�3NΎp��DIUUH��T��\\t����b�ɠo��1k�f�b�YӬH)ט�>���]2� 	a�d�TPާ\����.;���+��L��>��3�R���f8,��&��K�JA-�2eHQ!U3 �į�d��k��פ.�4JR���Q��s��m���Q�^��Mb]pr�a�ƴ9c<�"c6?E��h4$<��8˚$#dMN&Z
��1��2)22�/���+��2�p���W��F��#��+��E݀@�0Z`�@���9�7w�B[�젅&�	�J�5-�Z"�Lu�~�Q�aA,-f�!W%�mL0����Ƃ*dM���iSsH����
�q���˺ϡ?�y��g������\Sw8�{��BF<BEv�y�+�\}v�`��w�l8b��ϲZrzr��{���w�ِ�%.�Zi�p�q���K��[����|t���������o~��vd�{��݆7n������Fh2�ϩ��9��x���P7'K��x������9 y�*L�b�W��jB�qYC�A,MI:qa���nQ��<UX|c�9�҄�D:�S��Aw�� X*��i!u]SU�:��֮��4Y!��1M�\hvی�D�w�k��U�v��#�������{}|_�XҳWkk-VX\+'���`�@{7'���$�r�L]=X�b0j��"E�Rx?�<��;����})�ɜ���2
DPA!�"&K
�պ��I,M� a�l�Ǘ��t~�B�X�ns������ZK�+T���d���]��%?��O0&��H�mp�rx��׾�7o^���!���|�������p��}����p�����l�6����stt�l�@J�.�Y���Ų�xmkC��z*�oG��Z��9���� �m�*�׻W�������E�:����-�~\y�m�AĔ5�ϧ����;>>��ÇX[���CYm03�g�����MfX�6��:|��V�*8B��hR��#ovM{��3'M�0���4y��ޟ��'L�Ӥmy� 	��᧿��B|�o-���1�=��2�����߈�����l;j#��<u��m�j���V�M��\[+�9E�>X琤�R�ܤ쉫+NOO�N���9�o�f>�o���,ţ|r_��`A& ����K���>���|�{�s��}��!U�� �@J����(P�	USR-�9;�����?��)�ߝn��ҟZW-rcȔ��Vܽ��Wy����وJ|��ort���`h��Z�)��1�N��he�-���˔�`������6ӿ[�- j�EB�J$JI�4D�xj���u��Z��mw㷿gte��-�\7�
�1$R��֦.�|���ϊ&�Ͷ3دh [N��t������0��	�bww�3V�eY󕯼��h,��yQ�Ri%�R���Nc=-���g�J�� Hݺ1����7��:�3�ݜ�v�g�  @)����i�dQ����Op��k�(<�/O��j�*�%�-�	$��>3��v��M�9�ވL 3� $쵀����i��������	����y?g-�p��#� M�`����F\I)���?�W�ݼ�c�蓎C����k+TU�{����ﰿ����s��9L}�� ����X�vv�������]�R�����C~��1<�X��˗Y]]mnސ�a�댛뺤(�MA����O.�>���	�/���S�p�9DS��pOR�}�c�puͤ��Z#��p���}PN/x��H����pt�ϣ��2���.����)i#�ik��*�ڢ�	B������nۻ�plx 
BZ�����5�W�:���h�r�lRQ��Cʲ����0����XWRW%Q��R�ѓ���<��K���O�8sp�ǃ���#u���6��IW�����Z]Bb]՝A������r���p#�p8D�U�4F��\< )Rx�18Sa���y��+�(�y���n�b>�#��T����.
?��צ��>d,Ǫm��£�D	��,���z������7^CĖ�9i�Y��*/*am�kCʣC޻�BL�B"�"J�$��V�ID?��#AY��{�%�b����q��W��M��O��n�٣�=J;"�P�#|P�.S�_��{���7��N4�*���I��c&�!*2�P��l-�鏮�]�+�څR�m�.|m���Сut���Ű�!�|A�9!�ɹӴ��/�n�Y�X,j[��ח���p���������`0�,k���)˒�����W�Z�����qB�}?��sc�'���O�������b�}9>����H�,f��%�ً�l����Xw[�H��^�BI8�� x��$	:ߐ	�#�5Rx����R�q���W^���+X[����-Y/�Ҷ<dooo׮��/�@��x��{{{L��N��-�89�t�C���5���Y���0n�m4�l�2���i��k'���,��l��$nM����i��^t�ߓ�	��{��ߦ�O9<�G)	ޒ�9�p̷~ɀ�!Hw���4�}C����Ǐ��ˊn�,�l<�p�5oj��`m�1%��Ԧ`:�������!��״���ԅk
��)�?a�M�ע}��������.yp����Ģ���7o������9���������
�Ǜ�� ,9:�FɈ^?�dIg��Dw�4��x��MP���Bx���.���oY]]����<xp?,^$S7�U���00�3¡U�	�]����h����Wōb�b|������|F9έd��t���s��w��}҉T1�%�T�\������B�����&/�>ZG��=�:bg�����l���y��"�s��%Dg�&>3�z�5�u5�G���Ѓ��Ak���ۚ<ː��L�@i��e{����Z'��_�)�_+<k�4M�� l�R!�h���0�
����d;cʲX\
-e����~Y��n��k����&�	���
����g�g��ё�L����F^:Q�z\:�+k�a�#�/�w���r�,�� ٠e���p�AVJ��ټ<e�Z��l4�[�;�B�׸z*�H�H��ш(�(˜$������������C66W���g���3�������e>�G�[��(��#����l�SI�0)k�t:�$�D�0[�Z[�ő\>:�ǡ��^J)ZT�S��|��Ok,�
=��]ݿ5B ![�k�̡4�������H�g�)2���Y_��=��pM"�r��^Gm�(B�A��£A�T�u֕8_amIY�p�0�g���P�9u-:�x��΢��8��찰[ �$/N�s�=<s5ݢ��t�Iӌ�h�$I������&:D#�GuH�1�4�H��a��h@��U[$Ƒj����>��t|�/���q�����	Y/���R�z)e�?��|�Z�
P1�&SY8��Ԥq��2�m�����X];ǅ�A���%���C2�IJ9?"�,YoH:ai�JŊ(�w�҂~��f�Dc*��7����(���7�@�����=��#���^��hfӊ�k{-�"���h%I҈HKr���(x�?	uW�H�k �"�_0l���4�n����Py!:ZBK%i3����5ݳc��l]Ҭ��)�<�\#fA�|l/�
���d7oE����@�mO2��������I�1�����a0��?�w���?�7�@J%�?U�����+�|GR�U�g�z�ϻ�����~r8焋��	�����^;V�=k�\�=����c1[.����v/�i�l
*�5����`D)f����cl�o��7��u�y�wl?z��!zK�0���!:R	���p|r�`�#Mz��c�8���Q�5EQ���z=&�IW��� Z�(Uw��{�@/�!�F<��(�$a}}���-z��P/�(._;�󷼂]F'Ϣ{�{�%;ۀ���t�a��q΄V��x	R;�ڰT�6+��O�kF�DhW.���]��7�� �X�\�?	�(_S�I<�U ��B8�j ʡ��69y1k��,���Y�5�O\��2H�(�)Yo�J"�bwߦv%��,�(jKE\�x�^x���M�$��
��ίG���H�\�t�˄βGH��)�����"��;��5E9eZ�C[Ζ� HQU�z>-B��#�'���k;6�'�
t�$��XW�d�d|�/~�S=�a��%ta�E�#._����\�r/"� �f��;h����R�,�x���'K&�}n�>J�X�or���Aµ�����(&������dDD$:
h��p���\Acp��eLxk�!�z��by��z�E�vQ�=+�m�s���R\�����ͭ�W�u�֓$a���Ÿ)�H�p��.z��M{��\ӑpg�ݟ�tY�sJ);���xZ)�9:<A*����ß�ٿ���&k�k8�y����|�����y.�2�x\���NƫZ��*��y/�/�{<�cC�$�H�{�Cs������ܾw�\�]}T;����27�)���KE����4���b��d��T3F�>[�׈#���ڵ+�e���;�*��K�$I@h��G'Gd��,���$I�|̙#�t�܎%��
MܗpMK���-��$���b�z=��{KQ��,�����E���#}X[���^z��Wd�\5��%΅8*c�MF����~��qO/<��+A����f�ǟ�N!��E�bm��AZ����Y%]�^`�����Bx��g,x���Z���эi�j�oQ!@i�w5:��y>�xC��A`a<�~�˗�r��u��~��*��)��y��:!�����9�PQD�#Ԓ�H)�ܕM��7|)C0��iLU��"CHRTd��ȃMt�/,Z��s��N����炝H/I�.��zNGr��o�����h��G�$��`��/��*?����À&'}t���T�Li��V�R�,���S	�e6�p��ۤ����&�%��fl��1�%L��G������;4�}S<c �|>�4��`d�MXT�3���`��8��>��ܙ4����	�'�
��3�罳�-����P����8f���M]��g���B�ݽp:�m�����p����$�e����U�慗^������޿����E����l����'T�%k�ON���f�p��o���ّ���������8�� ���|B|\����y��&�m��l�p
-�
0��:�o':J��)5ei��=�ш^���ã=�6���~HQ�Y]q|b�N�E�x|�(.�
{>�vm���SJ��=��RW�i1ĝ�_�<�b1�ڬ-�<�ǎA�HR,��Hwj�e��PB�z^���/�����f���l�c���
(h�w�E��ؐ�!�,P+�v#�@���x� �g�>�pq�R�A�~4�_���_��x����	��U���(=B��Ƙ
c+�(%I�"�����-U��-G�$�X<��^�|6�Z�"M��DQ��|�#U�4MYYY�r�[^T���yM��*�D��'ME	TEG�B@)��u�#��7� )ΦAJ�Ғ���Ee1u]1�N��dYFU5|�S��pm�?�L��o�z�	��H�{=I#tB:��b�!N��g)�����c�jfv(���o�k��X[���
��#Bb�R�q!=RA�UH7�X�� ),G����M�^����*����Wz��x�T�y�uQhѱ<ϙN��u�Vqb�Ž�H��w���{\�pCגn��)��Ej
��s�2��}m0X�\b�����9��.E�U�.[��������i��M�|ip�m�T�<���SǱJ��������o��K/����XҊ���ƍ�z=����r�
����]�u]+))CI���[�[o��%��/d<W�W�W"�8a�qRD�*�,�cP���^�����G�u]s��e��~C`?�����4M?���J��O���2qj=#QAҴ�wtF
�����]h��Q�h4"N4U9�~�cv�k�����~IQ�qƲ��M�Fx'������3��9���\<�۷owh��񄕕������_kݥ3�E_Pg��7��9ٴ��ޓei�bmN�)t-;��0!'���!�x����*&�6���>��g.�s�>lϣo#�AW�5)*єEN&EG�|��V��!��w U��-�=���H���a4�ĺ�JP�K����>\���eN�X[gZ�@QU5UU�kT,�O�j���>�R�����.r"E����Ue���e�
��������}�����+_y9�9ͥ����
��/��n�]��BX`���c��L���2����3T��~kmC���������X�<���a�W�K�ʃWbʺ�zE������c�X��:!JRfSà��&�	i��%	��q8�^�kV��^3�`��]+e���eN:L��qrN/Yc��}���?!����_�7ڢ�'�B1�b��.8hqc
�kx�H9VVW�(�g�4^�?R�4ee�����:�'3��)�+����g�Bт�!�[�����,K⸇֊�*O)w�E�֚���Ά(̹a^L���ڊ%���`0 `41��-W��W�!�i0���NY���c�$ass�[�lnn�2ڠ,K�޽K�$lmm���#��9�� �����ϟ���<�y����w����Ue:�<����>��6�����R3��.���(k!���j\��[o�u�c�_�/��x1l��.rRJ��!��{!�Ctj�g=����p���*eYvR�4�U��SѐjC=�lo��@D][��7d}}��QG���G��,u]��:
�#��xb��H�&��7����t��YAQZ���7���[ᵫ̎ /%R��Izy���B���e�}k�ܒ����/�h;v�N�[~�?No'�4MI���F9�������v�פ���@h�FQ�Pck�
��BL)�����q���C���gg��'���/֗9o��k�����V.��p|<���)%�Y�|>'�Ť:�,g�\�φ�c��*7�%*��%���.�э��sM1�	|�Ó�o��,��g8Ҵ�Z�"beu��h��|ʠ��7G���(퉵���3�X����h-�g'���?��0�!R��Sa=�C$<�/r��98xȍ7�<_ya�A�`�D��Q��	��#/
��#/B������67���!/K�
��F*�$UQT��{�a4X�_��&�^�m���t����;�YƬ�hP��e��cNM+��L����;w�<\����j�vk���v�P*�R������0Y���z�M��������
��x̵k�XYY����{��Q_�����׿NY�ܽ�����,���{ܾ}��lֵ��c�w�9��\8�R�ⱃ���g=>��#����(�9'�t���>�Z�\~��ڶ��<���ڂ�I\��c�p=��cyH/�v`}/jՎ�l�����q��9VW *lUr��<�WPy@��-�4%�"VWG� s6�6��v����z����!�������X�"��-a�Cv\k	�ϬtR*�q��vZ�;��v��E���,ӳZ��X����+�jS+I�$D͝`�A���l��V�'��h�Pm��2V�p�!N���uЃ7�0��]-#�tqv>��}�t�d�?��%%��-m��f���6�Xou��s@���&��3��L��j�v�U��B(�X��u
![���"�T��M|��Zy�%���p&��,�B�H�n#�~�CE�աɋ�8θp�*k�[���*
����
c
L='�)�������_{�e���]��<P�Q@[#�p8R*��J�DxI"�ق�b�g>+y����%��ӿ~!�H��TL*��(ͨJͬ�QQD�E(o�r�:_{�޽q���Cjc���'%�� qD����~�+|���y��5����c�ݽ�/�s�ܹ��GO?�˭�v�߷T��(�⮋����K�\өq�u}rr�xr@�e"�)q�q��Z�|>i�C�1��x���Q������p���z�%;��Zs��9��kkkݜ����ŋy�׸t���ܥ�-k̋P�~��_%���w�yYS[h+:�Ҍ��Ka��3!�!����e������+��@��{JJ�Fz�!�    IDAT�{�kZh�����c��<�>eY�]��J�i� ���>
^bNڮ���dx#�d逵�67G�R��!�uf2p����F��3�i����e}�!i�����pttDY�$IF�$Ե�"�Zr��-Ue����C��Xۺ;�SEA�&��hbA\>Mv���RH6"�� g�zZ�x��
=����E9 �M)�w�)�C[�k�@�7ކ�)��)���v��E�v��:�v��`Q�dԠ{B@��=X���<u(���R���EԡގP.�S3 䂪�Y_�`}e��ׯ�#RM��!�7{ё�E���+�ٴ�'d(R�u�s`}�ݮ��6"�.�~���"k+*Sb�'�R�b���׿�������g�lz�|>�N�x�E���	�ϭ��g|�O@I&������ܹs'x�	���x�w
SC�N*� c+�g�d�`�;�X6��Ylr~m�ee�ޅ�T��NҌ�L�����4����.���}����<z�<�69��A���k���:���&�뛬�mP�5E1gw������?�1�*B������D��A5)0����ϝ�E�ϟ�d�t:%�SVWW��stt�TS;t$I�^��
 ��1�O(�^�h�JU$qF�FL'��N����s��9^x�&�	{{{L�S�1dY��/��w���R����|pg��/�e�yAkVVV��w�y��n9�a��B΄RR���������������/d<�zw�Z���.Fh'b�E)^
�&����1g�7�2����jUP�;���YV�N����>���.L���*[[�����)�6�p�2�M����	�X�,�ܔ
7[QT�e��G���<x��������'�s�$aee)%��PH���[�!���W�D����}ʘ:���E\���!t��8�����X�7y���BȝQ�6�^�cl~_iI�e�#}(V��(a2�
'�Kdѫ`� !��#}c�,�`�9����ؠ�E"t��-Ri��o��A�#E���g�������O<�X6ŞpOR���"HVV���7�䅫W��S�,[��pO�:�d�T����ĲD��
)u���'�"�~�l��l8�A�{����F�1��i6o���ˊ�����]�_;��)��/w���<|p����S��#��6YY���7�/}�Ud/a:=$M��}�������Q�BH��Y0zd��R�%��	�	�h����1DB�瞻w-�l�Qo����YJiJF�b��T���jDl1N�Im=�2�G+���-._�y�c�y>&���qJ6�&}��h���j
��>�����׼��;��:j���S5��Bt
�6�m���pQ��-�~���z!TJS��$I1��(Jf�)�露���{TU�����\c�CɈ��sD��L�ۖ|��Qy�wԓ6`8���	��.{��
R�e��W(���7o��H���q��^�=
!��H%Ơ��
����2���k���DJh�X0�}��]��=�}�����$鐦��i��5>i{7�nИw����H��b��367.p��UVeuL]嬯�S����f�&����Ƶ=�1��U�(q3�����`g��,���*���7��q�"[v�7�4��c�E����/��j�Ek��i(w�vN>��h��U6��SzM�P.dAl!���@��+�� �B����}ֻ��N_*B[�
"I,.\���9�R!�-w%q"�����k}#
���e��G�!�
���]?�}�g7�yE����˺�Ը\2��ڵk|�+�p��y�j�mK8��L��k�m��k��N�nz���m��YxHʈU�E�DIL�H�>�����E�aHe9�������W.l���`�5׮_a2�g:>�*J��D:c�_ޡ�����X�(�G���������h)0U��B��t:�,k�h~�d<g���$JgX#��!��~�w��Z��n�z���&�����u�ԜL��Uh#��"d
u����c�pD:ec}�nUR�S0A|��2��r2�b�GE1eY����O~�c~���SU����i��\���e��5a.˒�|��w��҂{mm�_|��xʝ;w ������A�M��$I�1O��ʾ(J�
?��666�R0��h��x����8fss�8�I8��=���tH�ݻG�\�~�<��ƍܸq��vm�]���1���766��o��eǿ��\E_m���v�:@�@�RI�r"���=�[H����8[�곎���}��]�:�eMU��<��y��@r|R3��p�,;�����\�r���5��)���[��r�w��9���ܽ����}N��R��X]]Ek���.'''$I�e����J4����*���->����=^���O>���w�����+�˿п����Z�F:�
�X(�������</B�֫���@4�7G@��V�L��;�s{f�p�$����*��ƣ�`�ӝ�%.��is�������Q# ��g48T����
_׃��3�c{{�|:Ai�|�\W�i)�.X	}�l���i�K�M^P�j!���DЅ'1^���ț�v��SCu�g���w皮m�O]��p�&/����?o�ƛ�s���m���>���Ջ\ؼB��ump6(r��)�uă!��~����o�����G��\;�xf�`:�3�嘍!�d{g��}��T��e���H��*���)^&��7޻��`�H������?���gQ�B+*�8>s��
Q�����xj�+�tD�`�lBR;�`o�����;��m���YY��e�uIU���no��`��v�B78O���H��TY�M'�/��� �K���8Nq�5�^AQ,l��:�&M-i1:+�V���y�3l�ᬵ$I�����C��@����=N�˂��u�(���9�Yjk�D�&;�3k;E��я���S�������H�sBi/�PBJi�.<8E�mbiE���K)�!b��z�4-s,�g<O{7��<�D���;�,KI{0��u�����F}�^�ʵ�3�N�˒���]8O������׿�-{G�$�ek뛬��1��893�Y[�h���[�Y���K�e�/�B[�"2/P�Ӧ��b!��=�����}�Gl=�
��m�h��"؄���{iz�$�eKhLӚ�h�q(!2�x�bmMU�H)�W��s�7�7m��\�E݈�G�%�?�aX�-��|Z���'��%tԇeN���oݺ���#�8��s��Y�^T�Y�	�7�\
%�:>p`A
�p ��&Dg)�2'�ׇ֤i�S�e�d2�,�ywjۄ�r��4�-P"�ރ�TE����M���6FԦ+��xop�RW)��u�DhE]��������.����gS�xE�:ؓEX8V���CƓ�y�P8g"�������W��[>�����VV�ܾͭ[��̦H����3�Lx�h�������T6�c#"G��CV��,��	4��䓒[�n������?�Z���j�zm�"$������{�庵ܷ�a�h��s�$a6����o�����$	�����j���eMk��q�z�eeYrtt�|>��_�Z�I�0:�s2�t����ۦ�lmmq2S�y�w:88`ww�?��?������g?����.���B:�]�p+�l��/�?���E_m�L����9Q�8V�>ʍ���F��DG�<�i�cpQ�	��e����`�P���sDh�Z'I�U���N#�	 Q*A�cBJ���j����Rtxd8�_^�M��y�wv�ȁ���d����ܻY��"�J�[�_cw�psJ��q�ҋ\�t�G0�?�dg����M67C+���ܻw#������k��1�s|r���Z��"�S�ӥ��S��Y�m�kreCFr�1P�_���&Uh[C�C��d�MVd��|H}BӋe��Z1O+��OA� C&��|�><yq��ƺ���I< R�T�GD�,`j��b�^�#6�]ccm�)��cU��4R%���c�$l�X!B¡���%�[ba�eN9�G�>��H�^<'�%B���S(J!�¢�EKA�<G'cD�%C&�l0D�����-�Z��Y�׶ЯT�����H�P��v�pB`e�P���H!Hc�)r�|LgX;d|,�	����9��l���A����`��B� pr"B�^���+����r�zN;FIƴ8��H�r�2#B \N,���)uY���^�э�Z���M��'�~�uQz���s�QMP�` $��}~��cNv��Ͼ�o~����$!���%Η8�k�7�y������_���Q��}�V�z�kN�czf��dʃ_�7���g?��ܕ�B��З�K�Jcs�4�H� I2�x�w���=���>'''�'B@�G_D������� �qK7�AtH���:�^Hp1r�����#}�-��`��&ZW7�8,��eG�,I�P� ���ׂ���4�ac�!<��
Q�'Ix%��$�Mf�	u=��_AG�a6-H� ��)�+�p
8B��`�'�F+8�u����35�Tp�Σ�$f6�09�Q"���P�N&��"�bp���\8w��sx`0u J��yI�qIQ3!R#�Y�)2� E��;?N�'�5����_���я~�I�޿_���E_��;m�y!�x�W�[��y��Y��
�۟����a}-��JRX�����w��������"J��C�:��k�X0�������Ehlmm�ꫯrt����i�t:����loo3���hD�$lll0��L&݃��W��z���e,�-O0�?�W��/H{����AkL0�n=c���X��$���U.]�ĵ+�Q*ؑ@���������{�j⤼k�=��FKh�0u@�A%8')�c<eY!�"K��C����A7f-�8d��U�)���p��s�a��G�P ��� u
T"I����Hc� �h�k(~]��@zZO@���X,"�'�8L���ru�{�N��ZŌ�#և#�sN�w(�YE�k󳞌�2�rHx�Rz�j��;7����o8�"Q�%���5Ζ�C*�������������%����Uf�O��O�͛�(����n_�����K�c�R�RAY8�u�S圌UY�_��� ?���
\�5v�D�T�M��+���Ռ�*��>)^��-Fh�6�[�:�D* �
�-��V�I�`�
g�BL�1E9�*U]�l�=)4Λ`g�O;�V��F���c�ܹ�p8ll^���
NNN8::��իH	q��c�ֲ�xo�L���P�U������Z�S����0���oZ�WF�QE�M��':�_�/�x��#��JL�ｗކ�+*��v�mզOg�C�k�i]z�rw�Σ�Y*�"�x|���3���ˬ��o\��>��`u��x��ct�cw����;��Q�
V���[k+\�|���-�s������n��޶��� ��a5ݴ!����=�W�l�v�ǭU���j	���������b#L�j����A4-��[H8O��|d����ۺ���E9���T�	�m�k
i��Y[nՋ�M��R�(�J!��?0���d���>��P�B���I��R�$��X�	�����I�/]��ڧ޼gc�����6�]�h���A4���*1¢��a�����@^�������2�8��
��"��rw�*X4"��� \�
!BKLـ�{B��V!��Mr����{���/��M�^��)����ȝ�ߡ͚������O�̇+��"dDGo���|p��7�)BJ�g���]���������h�XOY�sgkL-�#�3��wnq�w�Z�e}�S���J$D�	�����{�K�8�RD*9��Ԧ��΃@u����A�-=�m�89��!�2�V��'�^�w��8��K��ҋ(5U�1�ƒ	kPJ൦��࣮J�8B)��hN][��5��'��TU�3��P��JE�klm�u�q5���AG�Z��f2ws����$x���EenQ2�ʕ+!�c���l�e��r>X"9�!�C)���D����U�EZ{]
YW��*�s���e�VE���3��\��{v���HN�"M���������o8?�����V�׸�R
Q�������.��qtt�W(-��bv�<���f3����`����k�G�8�"��޽��Qh�dY����Y�[O"з����;����4?��?a�Ҏ�3RH)�|������;���>B�< �q�R�5'�)�*q�P�-n�D	2��Ea��z��������=�$j+�k�����}*k�+�s0诒d}��*np��j7$SHLT�E�fߟr���=,l~�X2�>���$�)�Z���DR!��U5UQa�G�4��p��iS�36l�w8b�p�" *a��8A"p$�uH,J���օbNhjkR��y�7���]���g�c��e:>��WDk��Z�|N�,C�Z�6�u�,�����!&��:��U𜌢Z�]�0t�`"��KZ�4E�R��Q�,�b�>j��Z��mv���Jΰ��ƹ(�J)��!�E��`	~�����2�rh���P�8��0��\й,<�8�i�"�u��WW��RjSrr�d@7��$�J"EP𛺤ȃ�6�����c����4~�g=:RX[c]��H5�3�XF8�I�OӔ��5z���T���u�]�v�S��(�Nk�ׯ_g8\��������ˠ_�sNHD^?r�?���s��]�_�/��X1lxo����ށw8����[ŧ���0�^����mW�4��n����$Iё�*s�}��e��䐣������>�"1V����!��`����d�ݻ����X���#N���'�F�΋��r�����{97��� �g�E���S/4K�x�����޷��l|��llm���m6�%�f��W�d2~�Vo]�����1��cY�eY6�����lk�[/qޅD����N�m^�0�����9�{�N(+H��N1UAU���\Y?���*[�xW1�3�}�No,^�<�gi�x����Q9��:���$�ܮ]�ֹu^z�%F�!�*�{���7?@��Jǚ4ӤYL�hL�֠T[ny�M�ƅ��&� pE��;�u��!����|�B�Ƃ�2���X#�2���Ο?O����p�i�R=��S���G�C[�Ra���!�$R1+�Оs�x���\ݕ���uU��yn�nh���K���y������siKyP�1�k$�������Q,��L`G�"�r�k?$�!d#l*�X��R;��}�rY`���8g�Lf8<Q��T���4�#޷Tp�P�s�*u�J~��!�Bk�X1�0Gp��a��$q���.%G���tʅ�h�%�akѴ�ei���̦ަln��_&�2���!�E/�{����[�ȸ:��ϻZ���i��U�E�H�z|����g5�nˈXˇ;��O�֗T�H��)�Ȉ(N0u��7GQNy��>��y�/����pm���&��)����bw�$�$qȷ}�hֲ�x��js�����c�ݻ���4Mê�1m�ܜsO}�/?��|Z�H_;�{��EkW�9����u6ϥ>dg�7n|Н�`$l���T��1e���æ�rݤi��p��o4^�vUz�ex��B{L%D� �$q�f��H1B
� "�z��mq��6�G�ń��-D���AC�5*8k��c���<]|�����PT�._y���/����&��	o���<|EN]�И����*��d$֡ �B�����(��Ix0��z���Fk����2��`�(����VV�HӬSOJ�9],|�����є�ߴd֖�F0�.����f�u�>ȶI�-EE�s���R���˧�r=��tu���,��B��s8�R^��HJ���=PJSzYڨ���D�t$��l�1�,]�U�aU��Z�bzα<��=,
��p�J���$�2�@�8jP��؎"��I�9�Y&��2���P�7]&Ѫ���P���2M�\eQ���O�����    IDAT���Ԇ�BE�^�Q[��d�ݣ�h���!�-�s�����k���sOe�ɋ���Do>�˷�*y�u�����������]�IQ����E-�wz7�`]&�����~]V.�����KHIk8�M)!����	�]o=BJ��y���7���ܿ��/_�W^�ҕk�C�
�#�*��!!�Uak��d��考�Cd�:i=[ې�����8>>fuu��ܵ(�2b����Z����(X��I�0���9�Ej���H����[��j泄,��d_ꪤ2QST+�dY��/6~��T�Y��l<�hb�N�f�=�I����� �Y�G�*�:�?����tF�KA:<c����8PY��4Ր̽���3�_�-{�M��i�D�pT��NJk��u.\�ʅ�5�Iƃ�:�����fK�$Ǚ�f��g�%#"�2kA
A�
��閙���6#-���as(�&� X���K�q_�L��������\�P�����Wsw35�_��T�zEJ�k���8=;f<��i	;��%�=$&��F�L!���Llq�������e8��*\�K�
��z��(�uU�F�����Fߎh_��!MB3g��"c�R�&��_��s�h��$�H��_Wh��z9�i%ƾ� ��s�#��T��wl�*Ꝺ6�i|`��o8}���"6-o�M�GB�zs����(W�}���ZKD8x�o��ggԭ�e%#14Ik7J[����A����F4��$;^�������%��7�&R/J�+�TiL��{�0�r�F�F�	�˪�����j8xu����'��ƛ��h}��MRoÙ���b58������E��_����gj�k���sE���q�j��TDt8��CY�޽�_�1I�(�0 ��]���Ʉ"MS�J��Ņ�('g�{p�������aww��tJhjvv��7Xq�JY��'�X��O��h8::�6nݺ�b����:mF����6F��1}���Ί��<}�^��8ŤX��R���p���,+R�C]z�y���6k�5,b��?ˌMчˑR1���0����!�u]����x�99=b�\�\�h���^)kOU���h4aR�t�4��Q�'��WH�iGμ��6J\>Ƹ���>��Yk�rK�;��cLPW�D/��5!:GU��Fr���O�0*uS��y�&���ɹ���Ȓ²�9==��|I�-(AK�۩"dYF�4����K�}{�y6Zs���3X�D^"aP�Fw[qb#�"�C$��/�����|>���ʑ�%������R��鴏���$����1�k�HB���Ɛ���7�xc��Iz�I*� �@Q��k]�Ջ�U��a1G1��������O[����.i�����3�l�b��Nz�Q+����ELr�TB��E��X�{^�=�T�D�\�9˻�ڐ8B��>��!G�f +�x��o��?����ۿ�?���NE6u ���0���$����A�AU��9�I<��ݻ߾P��}-�LN��i�&�� 0b��(���0�M� mp�O�1��*:C����buI�n̼��X�sB�r)�wi0%�UD��-�FŚX.�X�	wr>������L&�f3��������H�h�4�r1g�8g�� ��Î�S���y�Z=ٻ�`�&��S���v1����]���C�`�4��q��}����/_����p��o��S�l������*�������w��DQ�u:�&b�a{{���{���?����px�"˱VX�k�Rb`�Z��Y�	��-f)u��Q�Ν�����VG�"�G5R�%*�&6�U�x:��+><���o0��&����������K��xL�˧}���N"��I�[5/�u�|4�mEȲ�,P9�3n��g~�Bb�Ν�L�...cs��f�Z`D��g���E���)�#vw����,��`�Y�
����`�� ks�/P��1_&�k-����] &�IOXH��*��ϵ�0s�>�<�=�z����8��2x!� ����E&[�lmj����`u���צ������z�]thX�}'ǚ���.=�>$bmR��\F/��ϡS万`��@�o"�vi��:��E3���];_v⾲y��V7u�s4u�K���S�����O�ۿɽ{��w�GY,E���9e]��#�|����;;ЄN^-I�9�R� e���pĨm�Vڬ�e���ֶ���_ݥ��I~j{�K�mmm1�88�K��0�Z-�:�A��՝|�Q�8�IفT�8	�ߔ��������m�?\��bϞ�5Fc��IPE��FU�����d}q��i��j��{?,T��cJO �����b�����|b�O��\-�,P]2���h\���2�,'�i�1�TAhj|]��e"X�����^F!E�5k��!fo���9��2�1|ݘ���y��H��6�(��qy��M�����> y��U���S>��C�5�Q�%��Q戡�)rG�Y|������c3�s9M8??������Z椴Ѡ--I�T'�:u�J�g	[�����1�0�&�'pn\akmH�s��6��1���S��Ӫi����݄�\�-�g��}dk���[��1r���w?z�Ç��u���� ��˳�^�&'��� ���򐲊�z�~rNc�����*ߪ��~�"��h����E���37�T=����>'��~��V����Sr�t�o3z9Z�QP]a�z���?���7�q�Ǿ����Z��^u�_�UU��kqy�G��>�{�d#v�n2۾�[o�`]��~��_qrz�[o����{+�R��I���J}�&����4Ep���R��)�g-�ṷ���2��s�dY����܄
�2�)�O���d��D6���,��C��*D�چ?�{��o_}�����}��Y��Aϐ���i"Ĩ���vn��:���U��u8�LY�E�J�YBS��K5m�.����^�ΰۊ5��MZ�t+-'�q�Ybh�c:�my�4z,I��� U"�敽�#��(�X!AlZ�s��鰜���fD�e�����ڶa3�U�b��5'ƥjHqX��E0Zy\"��N!rz��s���ɸH��1�!�����Ua<����$��hR��������YT�Ծ�	5j�@����l�ɇ�)�kmJ���{@c-�Cr؞ކ�޿���m�5���|�bQc�8�������F
5�"�$��S��)'G'���;����T�yn������	���&�-b��V+Bp6�(�LFc\fPm���Ū�,kn��:ǯ�����T8m�g�=JQ�֑e0�ʠ�;�*�r=m�^���������Ē��6�k���y�?�%�9���_e��ĸv´K�>����f��G�߯/-���I�Ŏ*�Q{1�/�s.�	-ԧ���tZP;y�""qMk4�VLg����������&U+��	�4MCY�}֤s�D��h�!/:�t�eh�����,F,��͕�o��:�ҝ��c�*���g-�Q��朝�%�WǛ�T�*A|1��h�yc�v9���GGx��}#�\�>1�bLH��h�4���u������������t��~�����j��N����z �1��)�D?�^h�bM��9�X��7�/���:�V�t�&�ۑ@;�в��g|F��q��k��"��k,�,�9����(OSG���]�G�<��6Q7t���Ʉ��m��xRP. ʍ�=�g��i|�3��nN��'�
ʺ��!�Fd�4�ȊU����prVS5���і3�f�,s��`]�E%�{n��i��^��N���t�~
-���g��^�|�^�=E�k�8g:�2�LZ'�����rNӔT�_'���l���=f�m���lIU՜��pq���R���D�!��4�r�����������X��Y�-��ç>z��iˡC��1v�i���4���9|O�0�����A�n�fi�2�}������`K�Mj������u��f�����Nx�i����K�/fݤ�j1�ĸ�uϲ�Xe�8$��$Bu����+.3�
��F�]�nȍ0�nq�`��I)z��ɰ�`�����6��7i;��Ј0�'};w�u�	x��|_�d	���9182;�����������{rxx���uT��i�U��\��D�ЪV�������1a_�wƞ��+K(\��[pѪS�(�����M���a<O��*:|"����%�*Gz��cl�N�`p�]H�U��~9�`�z]UM4�1U;~@Y�pN/��_�:g�q���'���w>��F��j@H���
�s�b��T>2��:�@Gm�e��J*.���`gk�ӣcV��q��֘���"����HSVI�c�3*�c�mHU��boo��(�ǣ��D9:>��	H����s����F�[�Qf[�:���u���dY{�����(�:�W���6a`��1W��l|�*���o���os��>��}��Pΰ�����;�ܿI����9��X��Y.眜�2�� ��l<b2as����a1_�������8:>e4�0�n���o�Z��֭���)׍��#�tU�=M�^��I�E�L���c#��'miQX/�X����:F��=à]_��+W�b6+�t��^/���c����\2B i|���`����j����A�n�~�����9��sv����C��n���K���9;;�В�'j�%�D���y��S���o3AI���x�����4M_`ש/ucbwm��L�˅�.���S���|ʃ���J�7����W�"j����y��7�J����1}"��N_�@�c�&��VET:2��e�(��һ�s��%�rլ�{��,6�;�iYόe8��n�?��4mg�!jr��t�i�:�����d��aV���_Ԇ�Ʈ��v�P.��e��y�q��E�����m+}2$"!�7��y�=�2�7�N4���<��s^y啄��}�|�5����8?9�p�î�|<��<�f�&����ck�1*�����4JR���l�b^��H&�c����2�Hd�loo3���&T�S̏s�z\g10m;��t?k�d� &�����c"pzzʧ�~ʍ�XqL�[��H��튐�U��PWy>�(<���V�"�!2�looc2a�UY�������>����nJ��bLh��q�i�ez#M�m3T,b��ω����˟�*R�FV�z��KP7h7һO�Fq��W����ٝWM�0x��� �@@/E��	������7M�#p��=�������������G4��r�r��^���s�>���N�_������HQ��������`B�������h����C��`��Y��������u����KwOuϠ�TU�0��+�DL�2޻q���%�M$��Tc�Ce$~*�֫�m_T�Jl*�,N_zG �[�jT-TԈؐ�k'�_�+һ_��=�#g"������Lb���iA������1��i���V�4����`Z�!��EZ�-�i$l+<����Cl;��s�i<�����0�ڞ�:Ƙc_Rvx]_�6a�ԆЦA5�DIn������GTָ�>�m�:ӟ�l6��A?�����W8#_R��0Z㌧Y�m����R�:��l�+�^��믃��?���^P�D�z|r�r���"��S�RMkgyb��s�a�x;��)n��9~�hf��ެ�E�,IJ'�iSD��'Y�UUE��d�`>_��_��������wf4��������8�Q�5�ɹ�w�����IJu`~v���G�D��Ŋ���G4��9��>�7�S:,T�Oc\b;��m`�b��^�]֞'�M��TXs�B?�4�}`�Tn�E����v�-o��"�_y�p��uI#>B�4�����e��@ދ�]�c�i����c.V+2W���~�F-gN�4�[5%#�|4�����ƍ�N[g�:N&#)-��#������>h"�6.��Y��ݏè�p��uR��Q��k){Ʋi��9F���};�Y�*ĸ2bVx]a`|�c
.^����;c�髍ё�ob�@FD4���}O���������s�����e[�aL�'��֮HumD�����������P�
=ۼD�>�m�vm��k��6gb/���0�������P�4���q�����4D|c͢�^�$ ��x��J&����{<M�e����9�W?�Ï>����������-vvvx���.W������!���Lfۨ"�\�|������Sמ��)}�^��1;�3�����6\RGY.�V���b���?�=.�$�!���u�,��t���	=�1����jU�8��jŗw��T%��2��5��[os���+|��(V�U?�؞mQd#&ň��4e���!�G'����Z��1�ęƦ�����W������v����Y�y�a���!�}��9{�J'":`���G5tYߒn��#�L�١|d�+�y�o�X�c>��'�(���N��F\{���ØV�CM��� &K�٘�2�/�X!�`4�����KCţ˰c>���.Ҽ.�3���1}�҆�	�����᲌�Y�Tvs����JU��>��\.�hGp�����39}۾�y�b�oauo��is��MY1N3�^�G2I��I�H�>���(O��^N�_��i�Ä́(�j��s@]=���YF>m��2�3���A�e��TU�)��G�Sƹ��(�\O�k"RU����]w�Wo�}��0v��h�����Rc���]�mM�*�q�MlFn�(7h\����qt�«#�r|P�
�qN�8����Ҁb��U���~�����U����|A�q�:6�9yh�����{_B11Gp�Lw���8qT͈�S��E�qc���?d<��ζ�|�޻���T��?���l���>O�ٚ�(k����(˒y]�}s�7f7���+|���|��g���<�����u������P�S�m�'_��ݏ���)u��{�����l�'���Ԉ����`" S�QĸD�'%�ɩM���9���޾�b^bl����P����)�{�67��g���/������?��r����9���|��f�n�����C&���~��� 	�b���Bye�&Lw0�Ġ��^��j�B�*�Dm5E�::������r{=-��I����Ϛ�j����^���a�4��t�|�
�[�/ɰhm��z����N� ������e7�=1�Ք8M�\r�6�Ԛ.sqUA1Q圭��O��l�E�N!\{���؀����Q��^i��
W�+B�&5��(+��?<Y�c���5�pb�pNaGԥ�.V�Te�J�d�f�pqv�a;֋Cʪ5�D�����m9�wo��G��[i���5�^����0�Ƭb�=Lt"��J`�R:�k8r �MD�W�� &�J'������*��)�#9E��m8| (HletB�rhq��I��E |�  ��vM8A��)nI�Gy֓z&,b@0D ��(1᪌ &i������t�0*����JN�>�ͷ朊}��w͆�䄏[߇]Z$qߥAŵ*[[[�����l6��4�����bӓ$�q��9�����e@r���{�������^����o����O(lRI0��j����N���M���/�h�hS|3��}?�N���_������6�޾�̓vv��~倽�'''|�ŗ	�8��n���::�)�^�L�4�#��B�A�}*ˈ`�
�v�=�ھ~�\�z9��}?|���~/;+�����q��5|i����-��>F%S�L�#b�)3�\,��ݴg'g�&�Q�h8#���D����3�` I��|҃+(H���Hh�Xc��Φ�G���9�˨����YKh&Wo�}v̀k�c�f��+�0��.5\.�]
$E�������FWfɚT�P�+�8�ڀq	�d�������,P��'N��4Q�t��N�a��x�R��� �Ι��ޣ��d�P�ȇ�����{�p��~+]癴�xu�`2\6�co͸u�^y�������{�����!�}�E��N
��d&�t��A�d�_�>:,n�/��۫R�y��4�b����=��o���%�A�    IDAT�G���p_WM>��3���|�rV�
I�Ay�X��Y҇c,J��'z��
^\��4MC�U����5a�|�_5x���=jCR���>+uyu����w�L������=iR2<����{�o�IOAT�(�QSˊ�k8�k�6�3;}���L'"���1���RŘˎP7x<�����FD#N��ƚ�K$4X�����W5�b���V5h��J���	K2_��^��^ds�VZ|��B�k��+�S�;B�QR䍎�?����l�����Z���@�^��f��"3�Pb�a�[vg�>��9��S�~�Ï_!�s'�A���I���X��>˲��t�R���;��w~����6�u�i�b�[Lc�m��@S�d�e������������*�5Tu�u��M��0}�M8�C�[z?�DIҜ�>6k-2��8�kO]�,�Kʲd:M����ϗw?㓏���Ç�:`M�1	C:_.����h4��H��D1��SʦS'H�^>j�V}t�9m��c�������t�ۢH��j�(��0E����U��{��l�yl����R�o8��!h1�%� ��K��|L���]�g����hM.Q� b�1�1��nVI¦ӇHO.��fEQ"F����$j�5cHd�⒟��ӈ�R���*�}�>� ݂t7_��&>f��!JΡ F����I_,�JJ��$�ISVT���D7@��`���|JrGѐecn����ɛo�f6��fNS��f�Gºk��~7��4�fg�~���rJ�k�,�h|�Ӕι6�k������.��$1��NP]y@�l����F#[d�A ��
[����N'hU�%�O�'F�?'���o��c$�L�d��9*�pZ$U�Z���>������!��Ox���s��O����9>�G�elMv��a$'�G,V�t����,<h��BL�Fg����X0$^�.�����3d��{�����[�Ӕ]�y��e{������w�.ߟ:p���w��o���Qc���(��]۟�=���C'Nѐa�c��D�-��qc�ߤ"O�{rz��qs�i��C�$��a4���
���k�T$K`n�o`�.W j���ҿ�H_��cΣ��7!`���S1��	m�"�fkUi��#bɊ��h��%,"4gyR/(Ya0�`3G�a���o��7�џ��;��Qk
g�)���y��6�B�v��"��6#˛i��:w���܍I������Z��f��k�1�N�Ӕ5>(��+O��XuT���sm1����6������՜�B�S�f������d�5��R��H�_�e����$|��]V����|���x��Œ�������������x�>xL���Y1����y���̗+���4��ڂ0�ku3�Dvxͧi�+qQ��k���cCxA��x�^^���Q���?��5���%e-�2�#}i���@B�^5�уj��\|u=ε���swf��(15��*�ڑ��Y���t�?顈��T��;ru4
�1�jػ�*?��@l��قH�1��󞾤�4��Z1<��?�B��.��jO�����)�ټd6�����t:m9���窍��F#f���,��w44�).7��#C>ʰy��##f�}�|L^�	V�
k���l+��%L�Ӷ���6ښuz�����ue���c %���)���0Ѧ<��x<5�!�f���c�������1Xê	��SV�4�4Բ��^{�O>���914D_�:6%��雉&��%ǯ�>�=��jQ�l��M$�����	��ǜ��p��=B�GI(�KV��*z���ǆ�ɩc��9�o��ݞ������֌����|yD�=�EL��Z'i:a�1M}KJ�?��H!׵}kl8����믻{��?d��i��{�/��C������F0֦j�����?�\�7i������5��	��Mcc���"y�H����PcA-!�{	�8�h�o�;;;�y�MN�/P2l>C�P�3�Ծ!4��b�`3�CV�)}d�'�4H��g�5�~i�1(���uZ�����>���7o�d2���j��0d�ш�(zps���(�F�J0IM!D�Q�씦ID�M�5���G��2�u�?�����-��:��o�=�I��K���ؤhQ��Ib��d�����K��%�u��Δ�*�Ϝ�]��#�9's��hރ8��
w���/>g>����a}|pz�G�9�[��B7�>���6i�fd�D�֭���K��9��6�"G5p��>����q1?f�8�i�w	P�b4X��Np��&x�:�Q��ط^g2������[�n����P-*�T�<K����a���tJ����k�k�6�k�ܣL�?Jm2|}Y��t���\��n���b���b�QT�d��z��������Y���{.�Ϙ�X��Q��s�w�i����T���*�4̐'���IڢVf��,�yU�3��u��9jr��r�����NL�80XG�ΐ��)RhI|^!HlSI!�F/��81}��;�.R8�MSr��^�Zˢ��b������7�`�X "�f��-��� �U���	wՈJ:m������A9�8g:��'��{����o~��X!�)��lE���z?���ͳt��H��g���MU'<��� �R�Mc�0M�}�6�Ir�:���rvv�x<f{k�FW��h+�8$��U��ǧ�/`<j鷼 �x��7h��DD�N�\�牠�T�Vz��*�:ùTT2������cDb�:���"����(eKW�qqq�h4b<��s��/EQ��̤ȹ�W4ՂW�~��C�����;�Ai��!���,F2��P��d9�h�+r����Oy�w����.�~��i�}��%3"��7��r� /2�s,�K��a2�є��o���8
/�P`���6�tL����<?/j/�\=�X�HUG����Yx�'�ߣJC�RH���M%Հ���!PU�шpnd.;5�90�F��;;�Z/.�*0~m��;��FM�S��1C���Q�*X�#M���d
��H(PM)L�9j"Zg�=֮1�A�s��Ⱦ;7UE}"��1@�$ǃ%D�
>�I�+O+ד�c ���4�Q�B�TƩj�e`2�$�SV&-Tc�em$%�������jj�1�&�z�'�|�/������є/;��4��}�l0}�u�M)6��o �������38=9O�![�rA"�jA^��.�����K���xe'��+�<�W����yxxLY�lo�r2��d��*l��A���/�ě�9S��bLd4cd>?#F�2��������4$gOk�@'�mLj��BĎ"�+AXGT%�@f�I�8=�9��t�<Z�8���ON��~��Dt��d��vm_�]�ܽ���ng���
���!�jko���bqq���HY���
92"��Ĉ+�;W~1s.o#Sk��r��}�D�w���b�QgBPT=���Gf���.� ��D�uf�1��)��TbhpbPIE ��!�>`2�8/��i�e��%��;�� �Tu@LҀ�@M�l�bO�>�+Fi�M�eY�R��c���8�O?������K/���8��g�/{��ED���{��#�n2�F����9��޽����z;�!yF5_B,g	U[l�f�����_����ې�T�"�	��TeHT%���t6�Xt����o*���y/׷=!�L���,K���HӔ�u�d��e���5����]mhؘ�����i�4��jA�@̦����]f-��kV��#՞�vm/�׷]U�1\�e�p;ϳ͞@�Y�X��1�A�TU}����ON��?{f�/�(6�m�bl#"�����L381D�k��✏>|���}k_.�W+��QbML��;�o�R�C̞�Da���e]�Tu/�m3�3��&���j��0T�Gu]3�����{���9���a��������g6���#b���]�}����\RUu]����O���S �˫�rw��� �qA�\�4�@�T,.��O�WDٮrD�d���>�z/�ʲl�w-���ޝq4>0�888�9��E*�0�~�~�!����[=�v}K��H����ΰZ����g���G��%w�~Ip��k��9::i��5M��*�
`�!�P.�|�f���<MN����d�x<���L�I]c��c$gwwc`U^�喦IrV1�)�l�Ř��X�\�ָ�F�awk�r� ����M���9a���).˒�bѷW792�	�k{{\�4�޽��⣿zO�>����yHS�g0VԊ1��)��{��w����z�c���=��W�FFmQ\�DH���N[�,I���L�,��pbhV�|�q���C>��"7�/K���'ڔ�M�����(�jY��S#X$Eq�U]᫚&�ӗK�UU���!�oW&�e�{��a4����*w��q�rY����o��EU���X$|�J�z��p���e�"�-ւ(�� !��^7�>ǫk�?�u�W�Ɠe������ۯR�%���#��Ƭ�ˏ��w�e~r��"bD��Lr�o�U��y�l��Eç��\R�O(�r~|ȯ�����X2�pn�b�"G��ܥs���4	g��"�o�m�c�t�у�Dk��L�,U]�\�S�Y�D�Xk�&G5j��E#B���qD�4U���A#�g��k)�N��f�v����k�8��ʲ�����qxm��U�c_�{gO�?o����~�b0F�5��&���n޼��ō�)ҟ�=��w�������)�-�<ʺl��1�5�%���5�bI��3?t<�x�o�ۭ"6��ǋG�9,��W���8ɋ�X��M]VU�Dz��\8�E�C�V+���\<M㙟�T��P55�npy�"�F�bZL`*� z�K��*��>Pi�f�RU�,�X��e�ȋ0��y,��Y�q)�g���dY�V�n��B�W�$����6�Ʉ���s��O9?����b�%��CįR��u�Z��zYQ5�De�8C%#����/>~���C��h��̦	b@µE-�l����}� ���Quiq�7�|�;�����cV�c���L��V%e�b<)���Q�d2�ڌ�+U��TR�dY�u�H$���
2��Z�=�1_��>p��.?��_��_������Š�9L�1�u�x5��ڮ�쉩�+
q������:&�K�cH�"W�5���S��oϞ�X��k��Z� �HTU���|�ѝL=b��G������:$3HV��Ħ�g0i��M�n��ih�y��o���%b��X���w sC���W`\DB�$s��ƈ� ���Ȃ4�4�@R�h5�h CTPb*&�*�T�8 �4uE��T�+`MFf�����p�����E#6kٸ��9HQ�<Ot:�ł�GGܿ���!�Zsc�(�E4]G�,����t9��H�o"M���fd.c����(9;:dw��l�x��t:�Ν׸��Ërp�6qB�b�6#����c���x�s�h�Ay��7�ۿ��|��'���s��U���kϲ\`,WgL�c�[3D�ղ�,=1���8'+F[$�-�Q^P�9���9��;����bvp��;�����Ǘ_|�~�#�#�f�Nߵ��ܷu�$L��w���'ڷ�1K�y#��c��2��o�[�N�ט�?{f��v�:�b���*�X��7:��|Sш¦�}І�dy�Ү��Z��XMU�Q#<j�t)�0Kǟe�d:����m��2w�0߾j[�+-�#�Z+�#��k��P<!`l�o�<y�J��u���I)
�!�DJ�V5�¤pX��@]�I�t�\���U�ˮ|�Ҹ]�9�}�z���)���dY���>�W4�N��P����9�t�Sa+w�Y>�19���h��d�l6�ƍ�e���)[�F������wU%�e����.Oc�Bh��=Ս1���͛7����;�&PW��Δ�����7g<.�
G��M)�-��	�%�fx��N��bB�;l+?hPʺag�s�/jƣ���h��rō��kQ�k�f쫜��c_Okݤ�Z����c�ƈ���Bhv�>���GnϮ��\�&�Fk��Թli�� ��4*D�Z��0��n
n�U��S 27�p��h9PhkNr�VI��AD%(fc�G{,�����X�i�@;�]a����nL��v��k�1�y5o�,����t��
:'�;��HL�A#�2�A".��?��Zub]�2�D��q3�����	�⮃��n;��x]{w�Q�z d�fL�H0�&V�|L'�r��9��.+�嗼�ڏ���f[�ᢺ��k�1�@�R��&E�@�b��''�l���MB��������bl8�4~������t:��{wy��O�h*��7�M�Z�@�'9����>� d�\��_-ɳ1�2�8�|�v~l��y�f#���!8�h*"ڻ���N"���=`���c2��뺯�"�7����2��Z|��0����ވ�Ez��L�#���YY�U8kɍ�=���>��|�/��ⵢ��:,[z�W��1�JQ3������ʠ�x4cȓhyb.,�^�~{�=ɋn�	��(O�����/ُ# �t����ߴO�� R�} 3Bp���E`���Q��&XS�e��UxW����?�y�{��5��OĞ���{S䙫�1*>Zc��[b#q-���UX�a�eh�^v������.��[*i�H���ገQ0���V�&��ld�1;Ƣ^9�H��!�n;,���E����988`6�Q�k��,���L��~�mn޼�;�ï�ׯ���ҴE�`ggg�6�,�ma�e4�A"�/IIB1��\I<b4U���k�:M�}�1B�5>4L�#|�F��������`2���$��U��Q�o,1
D�c�T�h�(��`\�ƫFa2%�ؤIAfZ̆���hDY�,�ˁ��z���i��4Mr>��#�Yv������o2��uXG9�e9�*B����},Յp���gv��E���K2.�2hC ?j	��ݴaz���u��/�Jr��].�����I�52t\$����!JE�%�����?g�H���h���Ísꎣi�6ř����-N�N��S7%M�B`kkь�?��w�}����_n�\��'PV�1�,3��cb�+���Bւ���K��ڳ�͋("�!�,��|�޻�f3�g�̶o0��߿��=��%U��E�t��6�x����o/��yJKR뀸Q�~z��,k�j���Q�1��.)˚����_��8=;&9Ǯ'��a���x��]!O*���Zi���x�i �<C�Xk]�qbȂr�!F~�_�������OĞ��3��7�I"�1���E�T��=�${����m�B�N�l�L�pi/n���f}�YqI���rT"Q"Q�zNY/�}�ƒ��SV��ƹ���h��|� �EU�V�jA�G�N�Y.�NJ�+֦������"b�1pcg�<��f�X���i<(�3v�ʀ�a4v���INP�K|(���
Vobrh�}/��M���O@TT�s_���rt|�'}���vw�x��g��z$ɲ;��9�^[|��-2kk6YlvOw�C�%B"��a ��[�#�A����y P�<$j��iABJ�fi�Iq��j��fuwUu-��ofv�=Gf����UDdFd�/��%=�����=�,���ob����loo��u��޽��l����x�Z�qU�ށ\��h�����֢1fޖ��*E�r���>{��t�<O��!�������-�d]:��xɕ�=ǵN"�u�:bb��u<�����t��2�܎Sd��I �@4��j�U=��dǵg�*��tQ�Fg��f�?�"@Ϟ=�t6�phaB>L�� ���SXAVa���H]U� �AQL��_$�'*��s1���Q�ʢ�?Z� I-zY��J�O�0@N�1B�D�"v�	���w�q����CiP-k� h�	�z�]0��5��@9�FS(����� "`w�)>��
U��ܹ���h4�[�-�R�4�p8��=�y���~}~��ԲIm;�v��j���i�����柟eOD�    IDATB���rV���^
k�n����BT�bTUk�s�5�P
���lx��A���Y������ z  2��Pa,�)�O��	x$����&��d콟W#��*w�2����X�9P�
Fl��	9!����e	@��C�Z�n�����F;�L�_�V����PI��=,�1�e)����
�H8���3T3f��k*(��H���D���~��;����7�	�����!�=|���;��U�髯��誥����4 M�
�bŬB�B1��5��0������a�;��$�F�3uol� !�ab	A�6�k�I�=��pi��u��Z�� e$V�������1�.��s�6��x��9��)� ��|�s���e�䝄��'Q
@��a��"�"�,S��͛W��v���W�z/!8%�* D���(����m��������
ۖ�*�8Lq��w���һqR#Ԇ>�b�<ϑe(|T�߸��~�����;��t4; ��\=<�H���$I��iӓ�����|.�=�L��o�7n��H����^�\�=�=���;�ֻ����|@ݲ�52$��X�D�u�PS�x�������b�B|�?�s����B����y�$"F�H���3(	�� �`!^�� �����E�S���ܓjc��U����	Q��!��7� �Z���Q�T�^�7n��t:�{�F��"��hpG�kD+aԎqQ���2�<��n���d���~`�k�錾�z�*U��V�B�D�(s��{�XΫ[�������úz��W�p+颵D��AF��`r�JE�;�o�w����.b9Äj#�(j� I�y�d�=vvv�OZ��s�!�j	�,���E== �L&��X[[C�� �3��>���.{I�!1)����d
�dpFPU� ��B����AljA�3���*�:��	����g���� ��>G����p�]�k�
H��
��U���A~��c ���4��i{~�6��Dh�Pfn:�� � iB���I[lT5������1F|��g��f�y�fc����u��\�H�q�ڕ�"9Q�(��T�bϕ�1��_��\9���'�1�5�� �����g�U�HI�`�=�u�I3�:|���"�<:�+�$I%Yr���4�줉ʫ
-΃�>ŋ��X��D �ß�uv�"���XW�Ɗp�7���W��7�o�c�����7Z�+�v���4=�Z��m�/�~��q�1l�s�w}�[JD��p�U�M���d2�͛�P`2.����|���
����A�A]#r�Ź�q���n��|���`!�����)�ky�Eч6�#Me1ڟtt!w� � �}����X��펡	o��%�(s�&4���RK�4�i�@u��$I���������N��أy��a���뻼�Yu}~.ڨ���q��w�ߟ5�q�y��H<��,?�X�Ԍ��M V�9��9�z=$���g���!�4�T�4}eP\]���������������w��>@������.�{�ۿO��v��kU���p,�u$t]����q��[���)qD����S3�xv0b�x|S��vt�\�
!>/.�-b��x���,��v�B��ԤU�DX��a�����h�V���b|_Ǹ����o��Eh`�~�Wu��A��w�Qp�kG,���i,����݊Dn������PE28*A����=�TM;2s���|Z�r�Q����K
��*n�婳[e4.m�1�)���&|׺H�̊[[�uo��s,���풂��L���cgf�S��f�Zs���O?@٦��n�´��@���wtA�3?����i0�3�f1��)�L����N�
��x.61�� �C��$�a�۽`�K�Y!����D�Y��8�p�Ԫ�@�>t��Պ4��Zԅ��5�.Q�������;�����q�V⊄��ەK��g�R�4��o~� mf�ciߗ�3��`8�������sW����g�$�~y.$�Dishq#�ڻZz�P6����?��iM^'��>U�)�������VK�>����Ͼs�G銼�d�+y���n|J�k���|<fn% �"������ ��
�K|���WB�q(����"Y��e-�hM��Sm5w��@1w�&���%�>�q(N�_,�ڗs���^m�_�1d��F�Y� hjd̞E6F�����E�<�K���R�İT����eK?�t�*�r���)��w�X�m�&B�d�5#2}����ü/�m�ZZ)�>���35�_�֮�9����Oj�2'K�Y1	ͨ���Y����c����u����U۽�jl��܁��|'\C�UDJ���DpD(b�/���[�����q ~�HJ�_�I�6H&jjf�p�dBI-S�q��*�l�H8�����ڍL��H#p���o�OX^M�x��4V4�_'*tvWI�"�Y-hXT��"���?�&�]w�ͿMb���չ�+�C� � ���۝&�m62Q��wd|g�����Z�jL��͛�$�q���J9�eV�����d��{*a�bЁ�O�e����l�2{�bu��2�P;�z�݌a����ݿ���q�m�SH��� �n�C[���f�F�Jg���h4���*�𱱣�Ш�H��	��U�;A�0�c��W�B�������MqX�մ��!���D?*m�0�`�`YMa$E��g=� ���9:���W-�%��%�����1����6�+��L�W�%jf/Vu�0�u���s*��
��
�w5�F���v�e=����{Y�수��,�5*a_�j����*�j*lU[��P+,س鴪�9��y�?^��p�Z��>f �E\�r�"��Xq(�Z�k��}e>��Bɮ�V:�k���T�"E���8M%�M:E�i�􅲯B�ǰ�*=�Z��O���Hl8"��� \V��:%.y�����t�Z��_�g���V>/��W'��9�C�����Sc:�.��O�_��������ާ�9�ִO�_ZiѸ�	!ı�h��_��\�?���Y��I��W��G��}�e�h���[�������b�lQ��o����R&���E���Y��u��;�#/F4O&�7J|LݽD�:��\U3*]f����0�*�W���P��*���}��{ c�X%|��P n��1T�W����k{��֓��|�?*�{�Z[lO��k{�׿1�g�%��
�+Z�_,�Ԥ�Z� ���^I)k��g��(y:kƭ�N�ؠ�O]�j��j��HK�GөzGǗ�������B�X90����܁w���`{i&a,+;f>j�h����d'��%W�Qk��9�L�W�' Ai�gq�F� ͧ%�����f�u�o9.��)A�ny�_��<l��w(Y��4}A�^���h��ύ�6�"��`.��~یl�Kk�D:ퟤ���5q��l�e�:pF�� i;.�A��/�3�SEu�*5�^���5cC��~dO�^��S��#����֒$"�*�qP�7�o������yW���WM?��o�rMcu>�tJ��.-����x>dp��|���?�Ό�z�fَ��9p�+�̓��DPή=mO�����\�7	�FF��M�Ց�Tf{��RKE��:Z����<{k�����o�{{�B{.���vߞqU	�in�P190!΢miL-�O9j�a7h����1�}��z&L1�IF�)V�#�)����!��4v�Y�Wn�P#��P���%���.(���VCϕ�J6�=�T�%d�*�+�f����e�=k��Kj��צ.�92�6����
���a9�d����Cz2.�@^�QoP����)P�<+'��xE�'��=Md�;.K�E���x���l�HEt��p�!��O34"�:΀7M�sqlD������y���d�XN+�I��%�u�<�qve$q�RRi�/��4�ģ�o��XkF	�E56R`Vh�+d�K�-�t�s�S�6���mK������jE<r˳���C�,���\��P�Ilf�;�. ��g�zo,�eTE3"7��Q�Zьm��n�����P!P���a׶��G��3�B&��rK\������}�������GF#�����{\��V�D�Zp�/+m_E�[X���Xִd>��,��8呹	��l�K95�~���ңV��sqC-�H��fh�~����C��r-�����̕H.js6��S>[;��"�(hmB��%<�M��u���+D>����
�=�Ѐ�˱���,�����0� �o��D�	X���}+�$IIIk8�SW>0{X�%����_���˷M[ �}��S9�&S�I�������9�����sN���|��*!�4b�a���L=_9^��$��ys��q��b/( ^�և�>��d;�����d�E�T{V��Q=�r:��l"�Ft[Ă������9��Tg��/�����'����!�Yt����!�YMG2����p�´[���QDJ�AM|J^�1o�}�ƃ| 1'�!�7��G�7|/�X�C$L/��j?F~��ώ�'�IY�gã�R�"�d�d�ꆠ�:Z�ĝL��?�}zS�ëq� X���λ�VZ>-�g��Op}�S<��	Ƚ��611�LB-�K��v7}��탿��1�qq#�۝��]��*y�rF1Dg̽%�ʲ|�Tj�@����z�\
�~z��66$@Ʊ�DՒG�_(SB�d\�`2c�.0�=|f߳����W�^�j��[L��#g�"���t+�X0���˚� A��3u��L���|�j����C!�&�t�D>,�Z�t�������)��I=��C@��ǥ;��5�}:�}�[�h��B�.2�.�AR�y�!n�.��.\�X!=g2�8+�ThO�Rj�:�¢1k(0<���B���E�H��2�!-%BχŀZ�S�h�W�>�Y9��_���$�i��o,�=L�y�Il� m��8d=F@'�|HR�`	9��P��{��8�srѥd��t���\�ċ�� ~X��ݝ�3˔0�-�͘/�J��O����x��ƴ]��[_��G���v�t!lUP�I�2�u�/D Ք���L��(E�LG�7����bZ�\���ȴW5�,�\[pر����qد.���y��O���f?l�o=�~E���}�F�����>)�uS�e�>�����sڨ:TH�_��m����E�$:i�]~Ft�zҸ��p6a�I���Z���:u_��,����h	�A~sbR�U���~9o��E�uN�g�������&��d$R�4E+�9R���Xȇ$�/��W[�^wMY ���DY��aG�}~�����}̓�>Қ��o�tn��'6�.��`q@��4�@t����<��J�f�rMو�����1 e����Y|���z��{7�옾�Z�o�����:G~jK�6����TM���f������f�LF@�D&lX�j�1�3��Q��NJc��+1
�EL(�Xj�4���_l��C2H�-v.�������x(6���N� CJ� �\0�Y~j*����v��`�n�����3NRlWR-����������T������Ժ���WeP�DH����$۵��K7]�h���9�5۠�܊�����i��[/��.?�S�0���j�~a�FY�	<�Y�kGƠ�?��+5��@|��`�ge��`,VN9�3���$O����_�����q�Q��0I��Y�_&R'��K�>zF�
Y�T��i`G=�ĥ\�`����~�x�Yd��i]e��� vB*5�$;ﻩ����\��$\a\�� ��4g�Rj�V��\#�%%�@��|�P#)��q������8�W-����q�p$,�"����%�$�/�#w�Q�!���>���G���ĕ�C�~��'� ��޴#�&p� �zg���S#\e���!
��s:۱Hi���DT2R�������0��1���0d���ԋ5|e�2tvn����������������d����L��Z��2��1nf��CK�hp�f	;$�K��^�W�9VQ�1��r�u3�u�;��S��(&��	je��A��/_��Ӗ�Ц;�eP��U�[��b�A�d���1�����5	<��g-ԕ ����_�x�&���&hu�чe��]Ģ�?즽w��:�����]!� ��7�֎g��wGPe�M�����8��׬>��f�P��G��(����Z��k0�_��Lw�����'��w������ܸ
�gh��sUceLM�f�M�5G�g��ݙ3=�!���Rm��v�K�׿V���%~0�VPQ������P1��f^�,��� $hf����,{MkۂA�?B�y�X5�9׆�T^��}���SAy!c��Ie�������,��K'�6LY��2�z�+��Eمϟ��Ѿ��<	Q�����A8�1'�+��j{h������2��K���C_�(:o����������=,~���X�o�/i��~��ۧ��sW�a�`�@��M�qF�u'+)郎J��	��n�;l�Q������7��P{�:�H�-�Le�]���?����zo���@#����x����X���GM�4+����99��PX3O]���P|�Z
V&�n�e��Hӵ������.�ҡ�`E0+�i��0�}hq�.�
������0�L���n���/󾦫Kv��]��;���c���ZON����ޘ�������)�Sa�S������O��8s����_��/��������D&��v�[��v��{���|e!HN�vWx��3�P�lwq}�v5��V�N���-�T1����7�w���SߚF��{[%�̰x'B,^�G���N��UZ �����A��q���^��
�)�Y�6���Ͻ� [�������zݰ��	t0�QP$�W�l�lu�W������f(�)�Oo,>E�!I�����!��g�bH=2+ǚ׳�Jg���sC�e��0�)G��2����� ��6K�ڭ�P��;���@�2��%���p���~9��?tn7�Z����m4q��ˇi�\F���PzׯT|�\�J����K ���p^�H��͕����t��Yā>�qk��d�K��&SX���Я5����
��x>ێN���3�!
�Iy��oA�M>A!���:_L�w��}��8���H'�
r��=T��U��B9#)o���:��'>�;�)������z��Ҥ��!ɆA;K�WT~V� �VӀ��u奔T�[PwY\���ڏ73���A8,������i�!>?��r����n��g��̼Y�� ���qbuZ%���4�){�?T�@gQ�4|¿ո��`���c[V��4���i�s�������o��/�,�WN3��C���F8#(�l)�*��U��_u�5nZ��o�c�Du�&�[�z��O�/���}ă�ݏ�}y�>�?����u.ՕR,�1���N��Mν� .n�SqG���d�(�M�$����#^���<<A���͇��n��M������$�����x),����"L$�V�g���&�Uj�؋@N�U����������܌H�s�/����\�E�����moΞ�˓��:xm�WG�83���Y|�H����;M�:JU��r3Ҙ&�@$��Ÿ�y�a����2�:�4����%Ȓ-� ����tb�00��
�+��!�ib@���{i����ܬ�,H͇�j;XM���I5�?����@�tq0�U��Nx��i䕿g;'f������;�&/�֫Yx��DG5�t�I�p�;������e��"l�}�]�b|[O*|2��&׬Xo�"d�H-�����o[\YBv�|�o�7,�(�sh#2�T~�ڎ���3Ko��,�IH	cr�C=\n̩h4����Dگ�x�����-�'�"���k_�ٽ���"S�k�zW�6��ab۵����fK.�I-o���X7�)ŷ����U�-��Z>�v�|M7Fh(�U��tj\ﳒA!be�APt{�/~x��Av���=�^�X���XL,DG�'���G6�8q-�̧����@�m�0y�^K��������EG�uM�~����w�3a%�������ƛ������LO�g��n���n@*'�Sv�V�I8�]���.&NǞ���ã"��/��ؐQ$$k��s���c/���(x��J�յ�Ⱋz3l�G�RO�j�Wb�(�#��X���%A����o�&��s�b�>Z/�.�h�_��W�g�Gy哒!a0�R����7�g ���� �0�@�,�n�"tg���������)�+��5r<T#��ߔXɵ)0?Bo�F^�-�`0<�@�a1b���ƣ���i�D�#>g�1-�膷��j���.$�-4�����}�Á��{��Y��N���[kC9�퓓�	gj��FZztZ쌼���2����G��̗���\l_ϣ�߷��'d���Dh��m��0M��T}�5�#J*i�J�w��Yp�%����k�5��9^\�O��U�rt����rKK޹�Pm���&<�(v��+t�2<cJ�Oƴ}���9fg������4��j���ʚu$nG�
��џ�O���u�aJ��
��v+�O�GQ�����TVU-H��)d��֤��*�n���̳k�*�T�Z���.�5�x#E�4�c���L���I�|�*�/[H���C��G���^�*H�'ͻ���U�)LC��iz�q1C��o=�e�o�}2y|�3=�M��U�QT�����ݲ�L7��\M=�zmXw�c�I;Vj�P^4��e�3�S��/�Ic��`:���_���h�~sq������u�ϲ3/����v�<�?�NED�+?Zߌ�s �N+D�I��(�wPD��-+�$|	Y�g�$6+��.?�Z����t�3`��<h�Fru�E�K�qÚK{w鞭v��
xF�v	���"���P�D��pJ�Е鉜i�r��g��&��Ʌ������pe����'�w1�A�X�JAV8 ��4̬�����O5��_�89�?P���w�c(��f*�3��^I^���L�{M���
ΜO����n��oϪ�c��^��Om�?[we�v�6�������3r�w�\���l�}F����z��׿��_6,�����oq��-N�O��	���&j�S�\�Q��N[��X�j�xवc�<|���UИg���]=Y�s��`Bx�56���l;n��κ\�9��d}�/�'8 z��MNO����k���$B��u�qiC@��%����1)�F�~M���A�����@�����`z_Cn;]�wI·��?I�`\7�������E����d��gK�����1;TnG��r<���J���H��Ժ���y׽��j{�H��(Cfd���o�K���;^��9M�@�CS�����>�~n�q�����S蔒2&V���1���^�e�H׍rĵ`^����M��1�������z��E@Δ�-/0c��d�P�7EM�����w\\�h���&�����g�@{�ȧ�5�}����:��4��Sf����f�.�+�(�X~�/	��_�Ǆ��lJ'Q�4��18±<��+�_���	��<H���qo#����?MŃ۟!��7G�ɟn����ݽu��	"��m�cO���[�!/|�����6�;�
������y-��T�v���z7�ĳ�;��G��CPx(`�*!��yY~e>B��	��l�����{�H�@Ҽm���r�'n>�;nő����0"�F,��@��򗑨�Xh����Q�T�kZ�f�Q�Ol�����I@ȃھ���$�{� Ʒb�n�M;;��@���xOk�3����z ��o:��u�a�O��1��d�1gk��v�J���|���2�  hen��86�sJ}"\[.�+sL���}]�T���$J�+�3\:S����{�*�	z"�8�|fA�2K��.��긶����ո�3�M��5�e�x�|OƝ$K9Q���.J���F�6��6®0�>�
�؏ �{Q����q�oh���!M��2�'y��t ��V���Zy������򢍛����Vv��L�� �{.�3�7��� g�1y|��|g+W
7��	���xh*�s��0���T�w}� (rm��ӏ�b��")��k����JT��p	�H�����8 S�9Z'��B� �j>�DCN��J�#Lp�HlS�$*�D�'i�� ���#q	�$��W��G�ogfE��w�t=���yI���dbb�DS�c��9g�˰��n9޷c%����fb�(�w��\9����n؛��s��zF(LV�.}r���^��^�n{��vݴTX��jB��P�gee�e�@My�m;�ω���)��xy %�������)}�JO��?e�`ᡰz�,�D�VZU���o�Nd~e7��F�V��	�./j��ܲw�W�դ�����񅄈k|�*bb�+\T?�˟@E)�\y��h1�EB��'ؾ|Y{ۓ A���Ɠ���wϽ2�F{����aƶ��iɘtm�E���s_�&�_�A5/[������o�h��hp��ϹJ\S���7�";���ʡ�ӝL����ʙT�����L6R�I��r���l�?bA[̘gY�
Y�7@=s�P��Dl��ׇZ��W���K��!�=2�&1��G��6����h(�?��\�c+��R*9��)#�H YU��y���>��E_;���  ��f�j�e���Yョ�ޡt�x�_=|�r�b�
�7���T|'����G�
8�E�,^-��\����
.n�ӷ�5�A���z_!zSO�宩�f�I'":��������H*S� 0E���?�}��E��_?�U���7�W/�Vqf,b��L�4є`	M"�/,|n��	�/**��f�ṷ}w=��,�+fS����ᗛ���K1��"B	�ݎ��5Yw0��L'����:���k���`ᯮ6�4�W�s��X^��Nط�ѥ�^T��vPSp�<� ��iU%�����g�MFu��4��]cg�-���iZ`�K�B8h��`�����u�&CJ��a�q���x���b�q�$�F��]QE���F�A��T�́��2��F��F{��i��l���/}�H�&x�@+0i���s5(�us2?3r��@F�B(G�o�=Ώ��E*��'���Q��SǷ	�����Z(�X#�"6����y����S�IE~J*ݤk�O�t&0w.��O���(ͱ��0��6W.�A>�����J&��lM�6[v\\_{up��F&�A��@��ꭞ�,#�M�� �W���e������c���Ǥ���3�H��j��Bz���NҬ��v߾g?�:�N�l�W�U.���jp�59���
QMѶ��*�%��x�cn�u���"j�<L���гhtY�w*��$*�B�Ԑ�RiԬ�(x���hh(���vu��͏���rۀ�|��_���%�<V�JI�L��7_|O6s����mЗ��;1L���������㿖�{t�>�,5��?D	�{��Y�E����RM��� 5 ��܍�E&��M���UC�!j���d_z�_����ƣ��`d/�\ݭ�_7�v�q*���Yt��C=ӌ~w<Ɵa٣5��5!3�Dj�A�J⧃͢�5��8ס���yՓ�X�$$Tl��#"��r
�?v��5=�c��0� 0��!�"�ՖI���í��)FS�&#��CC���YR�r��-������H�\!�r�9�+|W;���h�2�j�^���ү�̨55S3��x2!�y>f�B�~�@�A2�,���0"�h��	�����IB��@Q�v]�rGH5��eZ٤�5�����\�����E[���2�j�|�A�k�R˰k��0u�3�A*�r��}����+�߁���3m�-���_�OW6t�����7lR\6�gw
b�q2�tJn�]*�X�G��;��=<R��~:;s��q��D@�8h_��10��1��y�Vl��.Q^ۖ/���uo��s��מ��T	��xV53c��)x�e�W�V��A�� �j;�[�h�7�(xo����5LEVk;��u�}�����<���HI�
�Ї�^�@xq�C��d��8/K��*q��=L�pkqk��g��g�Bo�C�k�B���Y���G�����/3D�\��v��}�cTs�"�my52�M�@�T����Ǽ�܁-�ʋdݐ����=2��v	?x��g%�ӯ�_�\�5��#��gU�j)�ȋA(�yS�g�l* !_�]H� �i��S�qs�,��Od������e-�;cFY����'�2�j�޾w�x���7��\騿��ԁ���V?�.n\�s�Z	MJ������5�I����>8��B���w����7��IOg�O�pG+���A��J�U�I����`*!��'�G��Y�p�0[�[G�*˅�}������4���1���N{����
_�Q�q�`�V����"U`*��g���wm�����o<�nٱ/in�&{���_P���&�Ʈ��P"��bg��(xڔ�B\FU�s�m~�����n���I�'��n��|��#U�<�>��T�-K�3��Д������SB
��<����2-����Z.���0cY�hZ��7�m[���X�K����͐�iu��铍$~Ԥ�Q���衆�M�S	(Dܾ^޶6�0U�^%�����'���n�=�0=N�l��T��\L���$l�����bM^<��ʥ_�#@!��&�(���8[�ވ;��PV:�1}�Ye"��K.�Sx�8=��
�<��tC���4��İ�j�$�B�|��	}u,A�����O��mc�B�T]��;s��$8(e��Z��j?d�q��6ӌp�#��\1?`l�^#��yÅd��Q�ح��Q��R)�g<M�@�ϵ(y�����s7�N&�q-jY�~e*�,@!
�*"$�I!�/�z5D9���f�ņ�l�Ww���68jڝ��0�K����*�Y5�O㨕*{�� -<�&��dX�^fs�:�Q�����_��&Fe�fğ�J��ۺ�I+�rp�^�܉�s=e;G�����`.�
w����J��q͵:t,l�P9�>-ڄ��	����7y�o"L�j[:���ow�s�\������HR����K�#&�K`N![^�C��LȘ��,؀v�%2$7>U5�������d��gP����Uu�6aF��J^� u18�����^�uTDxX�b�/�U}y(� ��uh�.��if��J��1P�T	��CG�ۤ�����*���M�%�Df10��E�����l��d#���5�������
c{�<5zW	����Z۝�iB�#�X�H���	--���|�����a���0o{�$SYm�kk��Jo�%�����
��Ad1�d'�{ƿ��g�L�����}�@���	 ����P\��pȎ�k�Nmuz�|��N���wnd�l�5��-���D0�%�L �T$�J
1F�%�����&���mGx �ƚ�հ*TJ��a��%?��SW	��檜�Y���3�!=�^�_����9�Ʀ�R/ɊO�vU�v��Y���K�߰Ʊ����E?iW����֠�%S�%P��Qa2����#a���#��uA����_���[�{{�Y���I�Gc�0p��۵�KX�嘼1�j����M�n��rYrl�����C�� iZ�*�o"��s3Ɯ����C]�������Y.�����=~��������h��h}���P���r���&>B���D�A�?ov=� &r
�o�!=(s|�g���,���ɀ)��A�jր���xr�Kޗr�!����~�u2�-˘�����y��g��66S�>jq���SaIY� (��:%m۪ʔJR�G9�X$b�ԩ~�K�Z`���[*<���W�D�-j
���^vĆ�!��>o�Jph�Ḛ`@��,H}��@�?��9E@'����g�+���HMU�.�)�5c����hC�<:ں�b߽i"��q��3\�h�����{��Ǖ���#�� \�~ؐ��U���zv�V��~�A�{�_w��NrM��&C~gn�C+Q���b�)[1�HD�G�G�΂���0���c{[ۢ��m�X��Ȏ҅��bP �Hi�Sy
�;9��"�W~�	S�
���m������A+j����sL��}\��D������{k5 yxx�&�?��o0���ݧsl�X��
���&Ao� �Y����7���:���,��M:*���פ�Gs��GA~f�Fm�1^'�42��yq����d��Θ k����5������[��,資�&FfZ[�=]Y�X�*�=#�r]�5pM����-�y�嘟�������w[���ލ?Å�I�>��(�hJi���3�+EjU�ɨ���'J��%uѦ��Z空�����n���eu/-{�դ#�5q���7��w�/,.fD3�`P(E@�����ݽ���3��_מ��k?;1���VW�2�ĕI~�p�2EAO�~2	od�?���'��N�+��܆r2�48 �~� A�%H��1��1�L��T�֗a4q��~�r�v|�o��4!T�tU��GP˛1_�؞ߞ�w3U���ԣ穀<Ec�"��/	���P���al�T4E�����ݴ���ܘ�5�1Y��+!z�:���ɋ&:/42)�����V��3�t�Tj�*.O�F�\M��À��*���L��K�*�w&�	�[l��H�����7���W(�B��?ц����X�w+�y��#�)O���GQ�>MSCq|��GI����M���뭨;)Щc�E�	��j��[7�Vo����	��ʯ�{w���b�C,�l��E�����@�3��j�-X�~��_����!��r���3Wq:�wI��7���Ns�|I��^�}�dO����$8�r��v�̊�H���p�c��7��O�+,��Z�;����y�7LN$�K*��IHF5��|�@<?�O@�8��o�g��z f�6
�����'.���/S�Ô�l����<���;ã2����,£Eb1f�V`��T����7�)�7�2vL���+��ŏ �������xu��@���w.�`F��<�$�#�h�:U�&����M O��T�Ğ=#�̫H�LE1SI�k_���}>���H���=�g݇�u:�ɔ�
���}���,���w����B�ϻP�I�*d�y�\qX�^���to�q3�a��`{�%���z}���sWmt C4T�OT50=LR��-�\Ǐ����ͩG�?�#�J�ɦZ5A0�t��F������y4)`p��*Ԅ��{?]Yˬ���W���ge�T{�uv��g����t9����˄�5:�A�^�=�(t��beK�4�l����u�6�j�ءL@������eU*S���vX����d����OjS�S3�L�0�:O��"��=w/9���~6�CJ˭�Ic��o�`z��{ϡ�M���g�vE9���wX�1�M�!̮Pm^ٞ����L&��"c�"�t]B�j%{h�����Y"qlG�@"���o���e�Q�b%!!!FM��D/�)�9���(=�/p���+ ���ږX 4`�?�����e�g�\�i��+S�k�u����;�`�.��Awl�D�`|L�Щ5�
طBƙ;G�׾g��G�c
x7?@.�Ն�~���h:����KjKYI�/	ɠ�H��H��S�҉��d��Mj��9��
��v�Cw�JQj��w-?�ne�=U�3T��nF�	>	���@q�M�b�*�_��<GlO��>����R��iQ�6���?�N�|_����9��顦 ����R�*(�f@���Qڿ��6�έpc��D�:L|�o�P�6�|�{-�y#;��Mi�3Noyx������k�8���$��ּꜯ�w���k���B	1�#Bm	��qp�t`�e�P1d��v�P��5��	�٧z��Y�)X*��bD�|5�����3��gS����j�Xb�z29���Z����"A�����7^!��M-J���1u���4q7����&&vo��W���~,&1߇ q�u�l���ۗ'-�]_�RF���Y����H������{	��3���]�yp��lk��g�3��$�[O���OJ�w���k��x&3��q�H�,At �`�a!Fb�[J���z��ũ	|:@4G��9�OR��0΀��Ҥe,&�8s��C��^��;��@ׇ�,���D��I��@=�Yo�q�۽��ΐ��`(�sG�{��նVϗhv#u��6�.�S����sU��^��X�}�!�I�O�Ԕb$� e��YKz?�̭E�c��?妥�E"6�� @��s��%=
����#p.�� �X��ئ��\P�aE �!����]���;�i5�m�e*�������Hi�P����b�3؟iV#�ts'��7�UظѮB6��lK�����y�M҉��j�Po�������������g�r:��f��8H�H�C)5]�����z\Cߦ��*/TvD�H�V	� ���&o�������?�Q$n�5�Q0��땢�
W�o�99�[7&��`������M_�
wy]#i��}2����v��PZ�b/^�ݙt�����yt�`$��*sS8���z|��I1Q2Z��Z�VG �y����vX,#R���fX �B�ŤX�X�?�	���x�:���N������p㕈HA	��iw�d��t�
���u����_�\4�������^�	?�
�M�e�~�₎�a�ο�	��r#���?��x���x{{k%����:WDi�\����_E���5S�U�YI���/��7�L?F�8x�7t��id�Kf��]X�{�W�|#�w��Տ���B�աINT��ֳ�}�22!�Lma���~x��7�]>O|.�S�`��7_�?�?�5�z523���7VG���]dޅg����$��c���5��p�Q� ����C�a��~�i%h"���u՘�-f�z}���i� �����N�;�z�r�Է�pD� t<�8���XI��:��)��P'�	
#��F��J.�<n�FO�LN��bݢL��A�̿ ����G�Z�,U�����	�G�w��$�"�EO�C7��{3@�ۄ=%y��&��lۗ*����؎�%��]S��+c`�N�hy/�Q�?���mCٗ�)�C�&q_{�����[l��з���J)�H�d�ym�ˊ�(�
��\�&����N�)p��z_��V��~r��	�}���b4x����'J��I)�)���O#��$�\��=�m�����������m޶2I|��eϸ����gmfo��=nt��Ob��8���9�7����B�P�E�O�o���ϲ�<�ʬxQ�����g����ދ��;�������BM�kG��6�ӛ.tY~��y��}z(W1��5L^[Ȓ.��]�K����u����=v�(��p��uͻ���P�t1�ZE�!������/Q�iR��L"AwGKwC�������^�����ۛPe���M��`#�H�fW�
i%�P�����@e���3�W��t<�c�ˠ�0++X�y�����6��!�Gw�|� �J��A$a���>�v��d� ��#,,JQp��^pW Ĭ�)�����POu�Q�(w�pbޮ�ПL&�Z�(�&�����x�I@�Q���/�#c2�r?+����%A�rF�R����w�?�Tg�r_�������{���=�_a�V��������o�`��~|���p�����0�CK
,�����훷?e�*�K�Xʝ��.��E��� B��
��|���fa��#M�y@0�	�K�Y���w A B?�T���v�F<�K�$6��=�@:@�	V��o%D�o|r�ѡC�e��vww1�E�iǓVj;<=���w<�` lQA4�i�� iR���2�kά�N�"ů	�ϧy�Q�')�]{��'r��{��/�o����8e}����,C��ׯ�}�x�ė^'�k ��O"s��Q!����?��p0�z�G̬�F�b�!��捛���(�}�Rĺ��E����>?��cb�xHP���4d1Z#Djӛ1�� ��� 
*d��i��h���ܖ��/Y��� Jd�Z�^�J_gy1�O�OC���75̌$�VO��tc]t{����1
�B �� �Nr������DS��|�9���ٰ*����/�����_��{�����R���ܛe������Je����anXB��V�L�.ݤ�}�k���/'�����"��&��K7�����^f���l�|RM/���>���d��;��t�kr"b�I����Ͻ��7����6��c�i��^��ۛ�9礎H �Ci��	���pN��+A�����o�e#+�z=(V �'�@!���H�5 Cf��
�DP�i����K�C�Z��i�_`��}�O;V�^�Β ^��|�p.@��Ĕ�<u���ܔXͲ^Rh���a�;�]"�)�*�7��?�I����[��9��~�s_:7����)�YGH`�� *]�w�p���?V�S����W���N)H�3I�TJ�g����>�v���x"��>u��g�(�>92Y��U���gG�Q�^.���P'����R�͓��0V�Ƙcjͽ�[�J��������8�<D<z�>|){�� �d�<�)q:<\<�`f���wr�@��QH��
|q�;�?��F>2sC�S�ӌ�A)���p/�[� J��×��>e��$��
1T���DT26:)4kd���V�@`o�W��2ɏ��k�Ի�V��W��g��P�������vP��4���f����C2 r/;?�hP��I����1Ed�[����={��IZxo�d2��Yi�t�w����;���GH����؟������"�{�h��*Vױ_�'+�W�ui-m-��b�r�#�p��<����&�1a��~~CSt�/���ʗ:%!"����D�Jڃ��o9sx7t�p4�s�C�Z��&�{�9�4i���q�� A< q�}�$ H�$9�Oi)5#�T��Q!��M+WlV���{�>��}��
�4*Y������ �2L}�x�2T*ػi�6�֥�W�+�[���p)B~2�j�?Q&aEdX�`�ɴ?����&��I����s��ō7�Ĵ+���y��\�?��m��3� �<����X����8{�,�y�\�y�|�<�r���w�܄1�Q�݈/����')�ە��+�< �k#8 ����Ȥ����СP�#�w/F �F�>��H_�^��\ 3��Q�0 �p��H�N���'ȳM�g:'��wΏ��=���Ɣ}3�� <�T�J��t���e@B�����Q�"�(HP�(S��?��2ڔ�ZUي�D�����Z0�MgG����V5+N��~��5vww!lmmaV��Y�&g�v.<���ڤ�6�z�hU� ������/��,��;��;�i�,�2%�u Gb�s6�<���!tu�g B�����D)�{�����Y���f�CT��t6���;�B �}�[�����5	}(���q��*O�.�N������Qณ���;<
����ó޷��]�J?h"{�`�Ƈo���so6����G���g�I��$q�ϒ�F'�}�[>���r���R��|�����}��خ3��ѼDf>-)?7�z����;�=��,Ͳ�F�C��J�� �B$"�
y�� � �uI����"D*(f��U@(��(&<	^i�"$��6+�B͊Ib�*#���H�Ib�!,���Դ* �\� �Z���Q��ڷ~���ج�1KD�̤�Zk=�I��,˰s�^���{�Lo�D����?�'��]���硲E���Rʧ�F��P���]���1�J A)�s�Cu�N��h��H�E�[աýx��?�XMY�:�P�^)�%L��"�A$�.H���A	)�B�7Q^�"@��h&�'��{OeY(�*��!��@/IRff�C<�V�v}�=��s�����G�^������ɓ��f���G:W��s�s�F��Ȳ30Z�9綈����.z����k��@�b��HN"���&�1������2���N��C���T�:tx���W׈}\+�t8�`"�s�9�e-.X[�;cHi�+�b�����;� >8�(xq"�A�V!��"B�YvΒ��O�S
���>h@3k��QJi���r�:�U4~xk�׽D���y>��%���eΜ�A�g�u�&�b�Clll�V��t�;w� �{���]�L�iVLo�?�?�ү�گ�����Y�)}�lr�f��mKfa�%�HH@�P���k���Z�[A��o]"���P/2z`�(m���Q�yo?f^R�����q�w���=���e�b D��B U��Xc�R��*Q"bD�/>HHB� A�D%�+k��W� +"�	�FR313)�t��e]�˺���b���K�}f/�Om����~���-dY���0�L����Z��
E�������o~3�~���Ʃ�-�������U���c]ҮÓ����Z��A�RXA'�����f���6�� "D�s�p|�:��p����C��6ډ��$ċ��z�ZnȐH�'B���\� 9 �&�q�ИN���i��b0��H O�!fM�}`kmduPꕣ-/ū
ߊbȂe�W�o��hI�ॗ����3��bVL���I�N��:�1
��֖ ��Q�=E�� p����_�tx���>}�;���Z� �L��D���L"� @���]T�����^Glj���*�{����ѣ�� �(����v���x����:Q��*}ǭۼ�>��<*�)��ޤM��"���dfx?.�:�13����i�I��:Q�;����V�ݼq�{�(�,� C�9sÍ>f��s��eQ!� �ij��A$yֻ�on������S������H�]f�ƀ��BbK ����zi���0F�V�4�6s,G_�:���Щ}:,���I�����!e-���z�!���2�h]Oo��kq.j�I[J�<�\�&� �M�D������S��E�/�p���}!,����^�G?�Q�>s����-����j_��V�$�h�&߶3��s�_��_�8^0<�;U���p`�@���wU�6D+�*Q��(Fb�# �߹���Б��G7�u�P����Y�t���f�ZYRט�ԫӴ�a����ץ4Rjq����Mۦe"��UU+h�s��]�~8�{0�ϑ�9^{�5|򓟄��,K�z=dY�;��6��eY �4y���*���a���W���~�N��/�������rG@v3���l2�['N�����c�q�rVS=�L�&AE��)�$���CQ�0f���:���YO���,���]m���y���GᨴG��[���A���<i�`y]*�G���qT��z><H�����쿣�J"�8�����p���W�պH�"V��8LZ�|�^�m>h�i�u��u�~�w��yy)�М|�Fa���������.�3`{{���'�$��[��N�:�O�=�d��O�������+ ��#|/��F��W_��ߟwtFw��ǟ��'gI����I�M�1���ꢬ��@�A���P�S�^�`�F��u�p0����A[�jGyv}�p� m�|9���"ǘ��1�ͺ1�<I�4�x<FQx問೟�,^}�"���
�~����p��M|���&�n���pk�Iʋ��w���_}�T��S�zU��׿n�^��Q��J���Y�5��ΖU1T�9I�*ɒ���&676�@��$�,�+��l���Y���?�>��C�Ԣ�9�A��p(��~{��6-��kCD�A��Df I4�"xo��p��ŋ���ckk!�z�y�<�#�{`����0�_*Q����n}�W�W���_������Lっw`���K(|;�^e�NΊY��e���I��Ι�8��^�\�qeY@)�T^p�r ]����z=��t<�ѣG�i��������|���w��1��qǿ�$�q�A���D��t�T��/MS�Ԧ����㻿����k���ad�<yŬBUY��E�߇��wG�����ɫ�;= �_����#�P�g�;5���'/��3+���~K��D�S���p!����>qr���Š߳��P��$�;�M'��"(X��=�*=ݓ�QX���t��}ʎ����3�(p�>k�O���,���I��У/�1�����>}�}������_��!��41M.�9�#��R��z��{8{�,>�����q���:����O�<	[9��3L�%��iT��wn��	�N��?���<Ҋtx���J� �dU��
W��/�$����_*f��^B�C�~n@Ӽ׳y��T�M^���B��#�S��v���Ӎ���G{�����yW��t�5�>(b�~���j���+}O����s�~��7/��(�,K�$	N�>�4Mq��&Ο?��/�ĉ �z=�GwB����: @�|�]��Z�����v��V��3�V� ���a*
C��>#���~os��^���Ui�W�$K|pN)�$���{���F��,ଅ��������ĕ��Mz�U��;��xԤ�Q�q��G���Z�8��o>z��1���?�wl?��w����~�m�z�u��A<Z366�8u�Μ9����x饳x饗����(ב��Z��ޞ�����1�ͤ��{U1����tK�u�궹z����f�u���KL��`�����])ڝ3"٪`�[;'w_��˷.����ڀQ�0����1��?�N���#��;��?G��q�5MSlnn⥗^��/�������`���[����{�5��)��@��ۓ$�RUe��J��i�X+����
� ��}�k��o���1�L&��A~{�u�����~p���������);33܉���IY$voJi�(�f���z!�JA��^����&��8�E&�A��񷸬�q�\wIBz�N���#\!����*���8��0��m�0_zx���܌"���:y�Į����L��`�.b2.���9ݻ��r���Ǆ�1--}��k�5eZ�?� (Z^��}|��,�g��Z���o;��#/�9�bu�����f[X^�`������i�X�+����o�w��ς����P�˺O�:�q��n���s����X)8���[*C<G\ybu\4�,�=��j~�����b�7k˥v_���a9G\���2O���i�a���v���	/ƈѦ3Dc�=�b�Z/�)��$3�97Oc�X2��p9��u�=�ݞ�_�� $	��:�X���`���^�Ͷ�9L�S����g�;}����!@��߁swo����;w��w���K�� r�����ކ���wn!�����7��ڿ����� }s�G>r#��>&����'v:�}��Ib�щ�TU���$Ku���ΓىS'�k�����[��;{�����H�(�.ԄB��-� GY�c�+ R$�x�ѫ�iy��ݣH�Q�����p��I;~_L��'�-�b����v��U�О��ui�#N8���`��UR����#��d0֩MW��&KXS����H-ױٳ��X�4����q�:Z�i�����'B�4�,��]�vߵ��>^麜���O�6��y������m]>��A$pRH͵��PUJ��9"Yr��2���r�:�T"�l6��I�W�r P���>\��Ƙf��v����kκ����H��X�Д�Y7c6���hD���oږ��c������6Z��<�Q�2'ζ�^݆59�~1fBX?�e�܂<���ً�ؼ|����곤��]��n�Y1��.q �e	�666���1�q��-h�������&v�<��    IDATv^�Ω���
�{cTU��~�����>�*XW"MS���e	�1�2���&|��݅s3����W�^�z�õ����a���i��+Z�[Je}R��U�4K�,K1&U�1��z`����o��y��M�g�z.���u�>�Y�b ���y �����	��t{�<G�"<���(�������Ԋr�S�:��������-�����:�����_|�o?�Wϵ��V")\/�	��}���M�"'���'����j�����
q�5�)�q���o�]�u���uM�޳�j�����:�6n+AD�(2qR�u���*Xk�$YCļ�ͲWq�6���eu�c��Q-�uH��9o[-��QJ�Z�(j�,�:���&6u,��F!���4M�k�[%=�ǵ���^��4MQ�%��+�r�R����W�U%�M���^%�]���.�s���?��mߧ�~���ƶ�Jg��C�����F���}�6nܸ�,�p��Yl�z�?^����Ac6��UƧ>�=x���B��_�1��0Q]g��G�L�(�+���c_�/_�r��O��>�?�]G�{��o��ܻ~H�4���$�����_����Y�J�P�4�3d���i�ʻ���$�~�����y�����G`�B A 0Dh!'��Ȃ�3/���C+u��v�x$ȡv��S�����C�C��=����X�.�0����ww�q�W a��|��U�\:��~���)_�:��z��X:_�	#�����C�˽�������^���������th��D��G�������3N��2ah����{�Z��������2��%"`�8vՌ�&>��B�{����@UUK�_]�UHD��)�2��<�6̲���&�J)h��Hk�L�~Q��n�+n/�r-Q��&�^:.֯m���5�Z����`�d
o�z�s���kױ����n�����S헠uc���^�V�G�g��g,@�[��v�m���R��~s�i�$�%�~��e���1�
a6��Zcju��*��H����}{��)�Α�H��Z����PFa4�C�ll `m���eU�t~oT��N�������]�rep�ʕ������w#�c��YQ|S��|Wk��^oP�keU��ͼcDBe+�����i��=,��2��
��1X1���� ��C�jӮ GġESp�[�:v��y|8�'���k>��$�i�A�r�vB��a�')�`���^<H����O�,�@,@ K@@ I�]���(���� �

Pj�vi�������b�W2(���Z,߽���O��������ʣ����Y#MR6p������= ͏����ܨ�/J���6ɉ ���.�H� W�Wz�\��=��:�*m���*��H��9vU��][�i��/~��#�J^Y��$�L��,��i���ܼ-V3/O�(��h�����KkmC�$iHO���~�~��,K8�`�bY�$I�r��G��LTۤ�.B�e�<�ֺ���~�'��J� Sm�����jz���{��������n�����)m�3�IDP�e���y�<�e��Z�5i�ĭ�OJ)�8qb��3^#�����%��_$���J)8琦9�,C0��*��N���� h4 �n�� ;;;�o��B��{{�U��V(K����7�����?�?_��?��3W~�J��u8K� \�tI�<��Zo���`#1C����D��%ȧ��,K%5�1������&�u{�w�ڻ��n��hei�� ��H�A��U�C˳������ e=6i��P���ں}�(���G�i��ïϭ��dd�\m��uXU����u��u��:����Y�t�գ���quP9��V��^�7��J�	��*Eј�V���sr��t��a�'�֪p��N	)��2�V���:ڪu��M��HE��d��H�VդU��n�6I0Ơ,KE��O,�lV�إi�,��~o��\�d��Z'�WPS{�KhaN���sB �f�z�}h��,g(�
֖71� B�N��sq~=�*$I�$� �9�RcR������) !Ծ�����'���5��ޣ,K��(����Hh�ב������8����'c�y���m����j�|-�tF"I�Rf���9�b&�K�d�'ܐ�<���a��Y[5��K�m�m���	���}3�"�t�5�3�e��aC򫪪I>���y���w���7Bo���g���y�&n߽��(`�T�w����A�o�������_)�\��[W��ӻ�@:��PIP���3��l03'M��։V��}�W���<K��r.��i/�43 e��8�v�;��w����=�2�I� F�F3/���Q�*�Q��ㄠ��2�}|������"�>�?�|G��z�<h.7�N�h>�������7��'���Ѫ?�:��J�ڦ��b�6�����b����?P����0����^����>�ܹ��h��H�&4͹ԲIk����fR^%�"�4S�
���U��6�j�'N��l����T��6o�rEu�MҢ�U�H6"��L&�m������ �nUU�iq0`8΃K����F4�NU�V�r(60�Bb2$��V��BeKx`]	g������E9�b�43�����3i8W�*\�`t
m����MK�`a�<u+�I�Um�$�_
˪� ��su ��<�/<�C��G�1޳Z�#P% ��h9� ��i���~T(��h������Z�,� |�͘Q+A@��*��j�Z���.�����X��A�1��<�c�Q?�����ss�n嶙����gM����m3'�u��֪��c��������t�ɴ�d2���&�Ҽ���mܹ�k+y�����`��~�O�/~��~nt�C�C���I_<�������O���W�~f�+x��!ȧ}e_~��A9����:�]A������}�=��aooB\��5~}��F���aJ�B��Z��P��}�v�O\�T�'O'=G�(��0�t?8�x}��YM����S�$�e��k�LŴ��iژ�bPF|��f���Gr����|I9l�mSO�H�	b��_"k��ŋ"��<jD����qRUJ��YS�U2֮�AJ�`�[�O������گM�������?˲l�Ik<gUU͟���`���~��O�UUa:�b:�6�9�&)'N�X2oF�e5�&��H6b����`{L���n�]����Idiִ�BiT�/>��Q��D��c6�-)�JŔ/u4�IL��&��s�9�9)��Y)ds����x	2'm����$s���n�f������Q�Fǀ�,��=�R & ���ʞֵK���KY���sEQ��k�8c@2�Q��8�G�@X(�޻:�̼O���b�<��4m^ʪ�p0��j��E��e�,�1>/b�͊1��:TU�J+mS���צ^ ��_Y���Y�������Y����ǰ��N�;ބ�B�����2��5��+��g����>D;tX��"} �˗/��D��>m�R�n��}��R�7�?jg�~���y���i��F�Ėnp����ƍ박ŭ�w0�`t
cR� �a��h�m��ќQ��'0F`��U��c<n�S)��1�ALC�����SќI�RY��H�=�B���n5o��r����f�iO�q"��/�!��=�k��o|�����b�g�T4�O��`6�5���(�E$8q�h�h�����v�^u$oO���%B�$	��>Ҵ�o�6FD�B���&�<�s�Q�vvv@D�lM,�/Sl��O$h��i�6�p8���.��h&���Փ4M�RUU=���7f��p�`L=���]���X�����4M�mj���� x���`&��cL������ʲ|~�rZ�����B��&�跴��ь���Y��r�ǣ���|E����Z~\2W^� �^��c���e�2�n�:[�c�/����{Hu=>!��=�E�F�Ў�m�x�R�y��o1��DP���CL�R���ǘH�3�&��eH�UY�:���<R�ZL�$&i귪�:��$�ι)�&����xi���\��u�������9�<���	��s�u>�P�~�ߐ0V�o���
A��?h},"��A "�����O�⠈-)� �>Q�E�v�(TUiʪ�B���AC�� @���QPJ��B�i�".�(��t[�V� ��%`�"h4�U &��V�����?��~.�O�. ���Ν�鷾�.��r��+��x:�_ �M<��}g����/�ߡ�x��/^��_�rz��;����`��OhCQn�E":����r���Z��t�1͒�x�U�0OQ��Y��x��N0�0)h�@`�5�Q���	 +��	L�!XW�*-�^V+���<$� ��P���i�7�j�@[-h+�A���1�����;$f��,�1?�z�F��>Ey�7�0^?��C�e9Z5q�	fkk�1_E�,��#�&����s��lS�?����S$s1:��NTVΕ�5�iH�s��%I�y^����	3*M1��s��h������M��bT��|T��m'�8�Gu=/�}!���X��9�D��M-�M������*g����TB���OE��&+����T�t�U4�IӶ렍��,ʲ�u��'��/�[�H{ۗ/��2˶�p��+�;�2�Ib�D�67�y�a�J^$V����aE��"��W.��]z���lU�HA)��F����0�`���#��|=�����C�j�"�B�9�����_<��������ypZ��jk����ֆAP�}]��Kkh�ʲ�1	B��y"q�	�X�֋��Ԗ'�� !	B�P���&ˊ"DD���@$�a9�IZ�Ê�3��z@>t�\����xϹ��x 4��$}+R�BX�E�,�$RJQ����2O K �CL��9��'�@`""�P�EH <�aR ���zAsP�,+vD��k�l! $̐���$��I��;@"A��B">!b�U�+b��Y��_��	#d��UT��t����ݟ��y>���?�L����A�  �/_N�a��]�PN��O���*����dF��aY���a�;߳�K�,�$�Nz�0��BH����N�X�QUD�(�i�<O6cR� B����ij�ۊ^�,��A�h�icTs�Z1\�����تI�p8�p8D�e9��"����⧔�x<�p8D����d2i�^���<:����l6����� ��d>��n^��R��ͣ����s��\�:|��R����a�##�"M3��1�ჯ#���H �4C�&K�l0)H��6�B�#&dUK�.��AԘ�j�!����è�(�k3�yZ�������o㱝#��j[��8��<k �s��E�uDg�Ӹ � ��R�pE�)��lND#q��D9��s�U��¼��m�w�?S��ڼ��^ӿ�����IUU��!oT�73; ,�T)^'�+�l�JIT�j�#�I���/�H2�@��+"��M~��פO� "�+�zH�E��9�HC)��0����yP�dA�h�l]pD��5�@��H�/����L�&B^���y�l!^+dV����}W@,
�"u�w�y�uU��^o���nN�4���LJD�H@�S� �'"$@��Je-��*[��2-�����	@��J��r�tU@��HB�E�D��G�1���H $�A�AAI @������2 ���sW,AẀx�V|W@=fQB<��D��$x�����)	 1	D��f"�~�pD` 3�ibė�kbH^)eCDLM�������(2b�)E�$�'&H1Dd"H�2�� U�{K�f���Ay	��#;�wn��N7�����L���G60��ߴ �ʕ+-/�>��7��{��{�0εҼٓ�U����T��,M�D�t��̺��?���;�ub��^� M�4�$�xv�Bو�H��677[*��RSTc�!�m,"jT�����Of�[2��sE�0�����H��&f����*���P�A��2J��%�|���H���KD�Ρ�*�������D�Jկ�<w쟓�:��CzC�S:4�~B��O$ޕH��A��{("�୅���5Rc�ZCs��! I3���ے$�u����{ddfݺ�MQFR�L����ؼ���K��z�٘���Jf$!U7Ш��k�����<����F�6���~9~��s����:�k,�U��)i	��{kG�UCeA0���9X� T�bɵ��&$3�8>�Ja%�2b�,_��^ � n�w�5в���-^�V�(�c�r �����Xs��3� ���{@+e:^gS��cV	���%�@�(ux�Zz���������ܘ���P[�}fh$����C��df$�0zD$]\\�܋��{I� `�,�ٶȔ��ڳz��<"Aw7���� ia�7my`�̨��XI���ԡ��Q3��Zދp�ʵ�#	�^m�������$ #@3/f�$�H��+uiXҸJb*I���c����X� 
@���5��v���2�e$�$4��w ʁ]2�sl�"C�Z)H������&�d$W	��=�Rmm	�F�E���g��$�@l�F	� pA}>��/ R�(���W�JZ�4��\�'$I�z-�nM�[�f)K'�p'�F2�S* D1 ����ک�m%xEr���&��##/(�'��mD��v&܂hi6��2q��%6 ��-�-V��kt2E��EDTAFh��b�w�j����=i+i"�vfv'��H�+�Y�h�����>��s���m������=�����������������O����T�e�9x�ʟn�G�/ß�c�'�0���l{r���N��R�����0_G}�a���uj鬐����k$2���� ��������G'���������]��a��~z��&6<H����<ߧ�: 뚫u] �#=߽��>������S�=J�?�ൃ�^ŷ�4Tv���NN6�˕�7N2�`�۲f�^(�nΖ�S	'n��ܐh	��B
�XriZ�h�i�D�� ��2-
����ѐD�	�U)�Ī�(Kw�4YA��&W��2B-!+0�2E��.3�����s F�$��2	�18��~��Ps:�fT�L��*�#�be)d��0���`BA�a����v���PI�̤����T�

4)�L��f㍹M]H�$P�)d��L/t/���%Pf�D���%�$#��,�~��\�2QA�R�^��(QS�H+���֖u2c�֧��@�P���}D��RH �G�	�_� 
JI��!#���:=Y n���}�v���Ğ�
��d鳼1"rE`�TI�)�h-/I��l�@b�
Ҁ0�М3cf���A ��2@ �4���3��h��o3�k*�F�SP����#���f��I�+tC/���u����+�@fJ���L)�H���QIb�q$A;%WAň!%8�;A'�m��  ��J��_)�KȾU�^���NED�7	�X�k +�'�8�l����=I'���6�k
��4'�Hy �m"�A��ɜ� ��p-��M�yVk��T#���nU �������ni �B��|&F�% M�`Or��IR��%��?북_��~�ܜ��'O������8��c�>���իW�����G���N�yi�+���"�|���T��t7e�Z�l�O`�֩�@�2ġ����x9�O���qdɎ�s>AB�p�Bz�f"p�jzT��ʠݛ�>�a���M��B�h�;�6��8s�������t�?4�P�5��.�D���H+�Yk)���$��Q��3�\���H){>O�{�ہ�."=�v �Q��)$�v�9�6�	 ��F�aZ铨g��Y�3����0M�v�XB2t�8����L;��׵���Ief�gt�X)����������}vP3�sg�jdP�Q�%47[����1�B]�Y{>-S�'�  �IDATϻ� �2R�y��Պ���80:<|�gEĆ]`�#���fB�}R �IY�$.��P ��́��X[�� 2W�Q	,��8Q$Ԛ��_�֚�e���fՌ�nT��[�sR�ݥԤ8egD 1��"A�1��,)A������3,(JU�$o�>$��=2�Hj{�5�M����Ho� �a��!�*�$�9�	��-�;�/��OI�SZ	��䒉;%�ILNlEn��H�S3���]n3󝄕�		�TK�#һ)H6�n���Dx���^]j��!͈�Ɔ�J�(ak�H����"?��-3�B�h Q%��ߴ��ɖ�7� �L���r�\�]�E�B�Uٞtɥ"3P%x,�=��@��V⍓�('U��q�d�RH����+��{����Lc"E��\͆�\���U�G08����6Rq5�F�3$�L�-�&���*�+w4)���IM��t�w�ߺ#����$2�-���5�朴pG��(�� k-�k�gt�TgH3����Ӭq���f���&NOO�f�������_��o��W�^�v;��x���g}@�Ꝧi�L_���6?����/�C/+��n����M@������8��$Ǻ)uܞ�T��m;h,�����=�8�����ﰎ���x��#�Ɍ#���*/�;�΁G �R��(�`5ph;#C���PD�A-"��A�:�$W7��-��Ks�=���*)�fls�w��T�c囓M`-^n���m$�������m�k��[@��F"�|]��B2(�P�d��3�b�������ڕEY�|�wo�͙���s��O?W�g@:�4Zs�5�W������L܁E�H- �N��WI)E�Ҋ�eY���.J�p۠���!` 8+u����	��n [6�͔�kk�����( ���x5)��x#q6b�Y"e,�˺�wo���,<!yzD����~�����ȑ�9����ImP�+	; ��!'�čB3L����aߦ�Nfb/a!1H�i�:�`�"�k�)�f0/��~��Z���'f��r�S�l0�Q��s O��g����T~f�gF�0�.�k�R�\��݀�!ٔZ�^Hy��i����e���� .����f5	�������ߍ�˔�ؙ1$EH�D
L-���vR����H��B�!�s	{$/�!I5�A�.�?P h�0K��( '$nIJ�(J$�0H��n�_"4���쓐S�D�<S�U�Ud �A@��um��+���\H*"7f~����R*;;�R�LH�6������d�_|�/hȬh�$Z��R0�h ,��KDld\���v�kF��b�j�Q�eb|)Е���
V4d{Lyr�zY���� r���8��` �%w�1ǛKRb���ZaZ��5
IX+���4�P_Yï2��L{W+�Rָ����zJ��lssz���;ȯ��*�����=�w�ޭ_}����k�믾�˯��C_8]�����_���o�����������_�ի�����-��|����EU��,��Z��0�i�4����8�G�mj����A�r"Pͬ���D�ѕ �g���, ~H�t	��;i($�~�F��9�\�eCGx7� �M�i.���  G%52Iq��ݲ\oo�-3��:b�1��p�S�F#�&��*����\�y/7F�N����IO133it4�\D���)!�{�M 2%3���fZ�"��г��֊�p�EȚ絖��g���\� ;�� ��s#��0���?���[Y��; 3L���\��d��-:��.h�0)���7����D~"� `�]�R#�~a��M�|
�3 ��ncm����	����w�~���1��k�3|������ߓ� ��ไ3
��wmk��.)�q߱%�g����i��c^�<!��]&tA����[C���F��F�fƧ��<Д���_�"��(��� |�@�X  �[%6N�*�6�.�$h� �=]��,�3 �J���[#/	m�)��4�)��ĵ�Sx�^{P%�;�{�F	���m�.�ې(i�-0p� �� }���L��4dg^nL����܆�"�&����r͑կ�r�(&��y��%�;I7�o�	if����\R��D3�-+�%z� '@[4��#y��}E�ȬP���wsY��G�Ӣz��f.w�����Z Jq钭A`�{� @�=؈@9� 9e� d:k�{[@k!��� �sRՒ3
��C��Y���-�e:��<���V�/(xZ��F,c�=��Xչ�7f*)T�eڍ��L|6���ʥ*��lD�(k��������>�Э����͛�>xSk\����Zk��� �Ln�Z��,w���`!� �Oc�ئi����NNv����z��J��>׻��ś/�͗��իW�c�������} �ӟ�����nj�'������l*�_M�|�����?+�gn^H�����͆�1���Jq7�.����5���I��3�� ��@�vR��� *�VX%5��A��4)�̱��W;�+׌Ʉz֘G/+	2�F�5���ܴ�g��ˌ8����R:3c�|ۢ���)�Y�&h t�n�ì������V�$9�B��.�fU�W7��Z��P�@��:��eYwkks��9i3�k���^~'e4(�	��כ�Dg$�م�B�R�m��	If�
�Kwvyf�8%���N`lۥtr�� �EK�]223�Pb��zrL2���R˥�C�ŀ�T.���v��D~"�ԀJC�~)7�)u�J��h��%]��IFP��Ab�sr�����$]>��� 3䚀���� ��Ժ��^�|U�%8#1��B��̼7)�N���a�zuHK�c�dy�	��.�*��	W����Z �t�@k0yxfJit }�?�?l��g 0v�%ݍRKX~fBK��akB�H	)�M��Q�Z��_����B܃��F�P&ҽ�݅�ѫ�#Jos���M��R6���um�R�ko+9M�L�<��@����k}��w�����e�p��_ʬRF��MS���� ��d���q�I�vw�ֺnطO��|�u��~��N����z2 �ݨ�:�o?��D%BelH�-����C������,�M �>��0WL��^�]U���YK���sؕ��~�eZƉ�ɾ�����%�' �a��4ޞ�v����[�8��
 �6��n�?�=����˟<�����ܞ�ɓg�!߼�B_~��^��J/_~�������c<�s�AAЭ\���FI�M��fu�/	~2��8����?+4V>#����W��҉f�&���TƗƣP;$n(�ӱ5b��LI����7�HQ`V/�(R *�eu��g����dH�h&5>K��id��t�����
3��NK	��B�����
p��0W�S�߈�4�M�U H����m�� \�-�u���J����q;όZ��kD\R�IF�>y��-���Z!5��D*$:��)0� @E�3�mf�+RA���$M�}s[{i%uH�5E&��x� 3����DO�Q�" `�`�,�0�JQf�J���
q%R;�H{ �������$��0��0i&	���̔��y�����L�d�(�/#��.����.-���(�@���i��?����Z���³�x�̜N׃֨�r`g#��l�ZoKQ!}<XY`YZ��eo-�����E���a ��{���,�e9M0��Y}y�o;��'����uX+[��� \�8p]g�:>Lo0σ��;��p]��6��eYUʠy^u�G뺰��q\8ϫ��է�O�5 ,֥!.�fX�}[�ۍ?8��k?����у��:}��|�߾̇��>^qh��ǫu�a�t{ sð�_�,���3w�u/,}�����q\�����_���z��<m�������.���۫~-oa�ߟf٬3�s��f�A�����(Ĳm������ v��w��x��W?xN/_~}��ի���6� �1��?8��W�����o���nv�� `:�k��,���3񒴉�k�Of�A�_�`@R֋1��=L/�Lu��ƍQ/H���{�P�&�)�\�͸d�dC��� �������U�p?�Y$VB�LUR��AO?1�i�ש|����h��{ !r0 �v�c���4ebDv�����(����1���=]�v��,LLh�AQ$Y�7�|XVZ63Xʰ����_m�h����|5++�A�d>e�T�<3��ߊ+���d+��%�V@rgƝ�-i��ꆖ�Fz�֙(��,ꂺ"�6�`fm�0��j�)V_�դ��=f#
V���'w�hfvkV@������fV#su	�Ze�ȭ�uW�����꺟5�Z�=�N#����6�~Ts�Ojp�c2�NO�ED��:�v�SEo�>׋����o���>\w\���;}��x��+�˗_�͛/���� 8nw\����a�����_����V p~��wi���i����xr�A�<�	<�8���7�{NS_/1�a���S��ސ��Jv��ZƱ��c�����wG 8Y>�P�f�q7�=:�o�z`7��$�ۉ�2r��sYfN��;��$���fk��i��z���V纹)yz����������|�m?γgo���}�;��O?}��	h~�K���ׁ��?�^�ze���ן�>��9�����5��_�����_���Y���>���1�)����c��V��4�7c7>}��_��!�3酴�3.���XO�� %�ޘC0 TB'�vNh��7���[*�tG�^����L��>�N�>�&F��pD&�P���mY��g���,׶<s��B�+ɯK��� ��xY����\�J#'4ݑXH�\[�@�j�[3�0r=T�Z�Յ�ȴ-����P�����9�8	��3|=d��^�e���ζ�"���
��b��a��E���R�KQ)m�`�9Pb]�܋�|�2oUc�[����<�P�ڙ��� �8�pW
��K,�iXі�2�h��ke����9�$����\d5n�Ǫ�o�Lӓ��g�a��cĊ���E;?ǰߣ��5����\Ob�R�6Sm�5y9_\<���Rʙٮ����N?\��!�t O_�9�ޯ?=,��^
���k�3#o�>���#�:h�7o�����_~������a[�3'�u��x/_~͇�>\��s=�{m��7��9�`��/�!^~�/.��˗_��GV���ա/� �1��4����O^ճ�����~:n��$_��!����2]��O;��Mf�@�!qE`1+����^�]| �J����N�v�׊�V�j�½�k�rH��)��c.<JA�>V3���<�}�2r&=��x+"[]��W��*��e.�e�(�ԝ�<_m�mm�4�-��,eЪv>Ȃ6S��tW�ڗEcC)�J'�9xk�9֕��4u��a�0�˲�f�����Z���C��I�]����q�����,�L;%�%�\{?����9PV2^�Xݹ������n��2&�I �d���6��%6��X�^e�s4�~�+e_���f����,���F������v�Dggo��_�;�����<����}��>\��I���#�x��x��x��o���> ҽ[��ۡ0W/n���h+[8�+q��iC��Zc�CT.�ʗ���G�0���B����S>%=2s��P�P<5(s�b��t�iLN�g��+�Ĝ�����Z�s[�7m��c�
 eַ1�S�=���|�7�� ���0����nW[[��C�J���t_jD��Ϙ�%:��o ���M��#�u7jwW�r��"�g�%�m��ۃ��+Ǯ!��>��`��lnm���!��A� gg�����_�`��__�_�I����<���x��x����s�Q��C�?�i��ؖir��l��"���Ɓe�lM��>�q��u�6 �����ף 9[���ib���RV�y��\� ��]�W��Y�Png-ۑ�Ǝ1�4H��q�C��~ G��t���@tqq����_<�A�c ��{�ꌞ=����~��y�+ �?}���<Ԁ�P|���ݴ>���1�1�1�̠�a�'?��}��%?}�������/~L|~�����ы.>{�#ktd��/���x�� �~&����~3XzD�����������B��K��    IEND�B`�PK   T�(U��!�D�  Ԟ  /   images/cf2dd1a8-295d-437f-92b8-7fcc138ae9be.png4�uTT]Ň��z�iF���n���n���)���fH���|k�e��̜{������މRQ��zM�a��J�?c��4�<u��Ar�b^�+]޹��<�B{�������\�K�B�EБZQq��SH�y����87�����o����b_�,��9X]�'�O!_�YM�cMO�S�ր���nS�[#~'���SB{��7���	"ݚ�g��)L ŪU4y�����[h! d޽�v�YHl��T|�S�F�>,��	�Qr�4Y�@>�T`Kc򆓓3�����=<�$$$�?�dff�°Ȧm�A�\W4�^l��r��!S%u��m�=�-Uv�q���)$%�_k8���恢�u�����G�j!��A�(g��r/���n���OOO��\�H�ژW��}���!�A���b�ԟ�! �0�,~*<V�i$o���=_���YD!�rL�ӶyV6�y�Q��>�K;�MV�+v�3�0-���c'1�] %x��8��������.F�6N�6�j����N����L��z���D�u�����ဂ�Kh�#�R������۴Ϝ����Q�J�w5�'�TB�G�琄����q��|����ٞ\9�s�\Ԟ���A�AEA��s ��Z5���͟���<s�P��I�̋�ƥT3�Xq���fFZ��d�F�h錓��Y]����A��ur�bR�n�쐝(�0X<(a#���Ό��Zg30�2dq���ai֭��N�\B�p��n���M�ɴj��$"Tޥs@�a}���(�B�3�����@T䘘����gs�@?J+�&�4��@~a.��au��E6���"�s���s���-���u�n���b�g3d����L@z���L�͑�숀r�{��͇5ua��p�����52�)���~I�ό��N�x~,����TI$qɁm���>��,�4��_:��8Ej,�nT,�"�dr�3���zmj��(>�>5Z�7�}KK��,��y��U}�8�d�ݝC	?�3U�9�O��}&��̬,1�n4J�Ŧ 
`	uk���%��#Ȟg�� q3�(Q��> -q�:���Gq���9����A`��QG,.I&���Y��I@b�����]鶟W~^
��a�����O�	�镏�~��2Ţ��;��������/}���;\���-8f��v���0���������U�4�;d�U���h�OK����L�/݈_��)N�"�'��!N��sFr���i)�i9���I@�@���5�8�ۈ�|*;	ѝ`0M*hڂ�PNX������M�Is���N�����a}�������ڞ�(�����`�5���X��هl|��2v���N�feC
R靾,�X�d���b�J�>A``�����Q�F��=)f5�������kd�3?*|c�3��!��(d�(d���Y�"c��2�����W3N�+�Ӻ��􆇯�)WZ2��حwSt�n�`��
��u�&)W�a5/�#�� �xз���۴ח�_!��y�g)�n�������GC�I��qԨy?�ZS�WB�R�ꝓ$�{!X�.��:F�!nn��Pξ�Gbl$V��+����N}��N}_�P_��Ȩ66{�ZO6�W���J�GMmm_�I#��ˤ,UJ�W/b�I�YRx��~UG�u_�6���,�wan�ɔ�2jŢC��D(O���;]$!���Or3��.u9�./���=�[��u�^'-�6T��D�?�x~��H�/;;j���5�R,M��ݵ/�	2����"7�掆�G�M��}gI�j���1m�l������m�#����|��K S��JJ����tV�fqZ��f��<{�x�{�o�D.%k��76�Ag�LD1_Y0�ˋ�j�eP�8GCVqY�0�!�o��o��9��d(����YU�s]�tY�~üxB+o��U'~(<}8��zN�\�a���1
�ơ\l�_���4��N0�Z��p_-Y��Oe�m�/}��2L��6e�N������}7�|�v1�m&խC��|0��EI>�"�j�6u3�B�[��p��� ��F�G��AB��w80@�^K��;�Z�g�K��_n�$ɾ�qӭ��1i���������$HL։�� �#�,2F�F�	$�8CB@���ʧ*�q���G{j2L�UZ'A�����ۏ��=��m���Ï
�o�>�XB�����q��k��K�h��e�`�aэ�ܲ�3�` =�� �"��օ��������T�lwq��T�l�,.��h��樻,�?>�?Q1���Ԙ J�bvjD���i	�$�������Ӓy[�4y9��Ye�����
����nad���;o�(80qF��� :�c�ǁ�YN"7�ƣ���o*�ߚ��"EyQ07�=�Gb͏�dc�g�3��gB'�LJ�K������W���͚�46
&��H�Dwp�}���R��{+<����,9������݆W?>��p	�š\4BH�C�83�#�\�a(fP�8t')O�3Fn�t�����n�H;.|�uE�P*ư�v�Wn#CV}�PoΩ�	Ҫ7dm ?��"��4����yV��ʊ�$UH��S*j�lWM?Դ�l�V.���]]]�yyR�I�%3@T��<�P3��c2z�BN>8:*{%�{��8������YU���N�twƞ�u��9j�c�{�t��B�ȑ-\J�1�60��7Ev�O�rgreS�$ޤ�I�"�����SZI���B�U-�ۚW?�ʱk��l��lD_po�� ʹ�q�ܔ�~�J�NCo��8��!x�Z�,Ftϧ��̜��h�w`M�������"�uT��ONmB�����gm�Qx���L�c'�\>����Qt�7�[�\�MH6V^��Y0Cq
���a�/���F�4a���B��6�jX�پWTV��\��4Z/\���p�*�r���sѬ�$�u2>��9_D�mp�M	��P���hgc��QS�u�kӍU�;�
ի)Ra�d��ۮ^8�n����7�b�L
�jL�N��x�Q��{����5��*�>��M�����oEҠ�i�T�%#&V~�T�ږ$O�m��H,��`�z��;ޙ$=�~x��g+���ill4�-2�Wx+���ǲE��~�#m��co�E,���T�jo�v�xa�#WWW�E��;��yX���ԝD��Xo�Ir[w�ղy�g�V-Kjڶ�:�܂�Yy*c�9�T���	G�����gFI��B��+";�I���ݳ����u�I���������|Y����(�ꆎ�Xl��c�gvU����v�90�~�V��5�X]��)f� ����l����pP����rwK�U�,x�J�}Tse)N\�2L�n��7�m�&�z5ZE@6 b �dc:�/d%u��C�,���f �$'s�<O��-x>??�Ƞz1J��"q�L�/
���r�Vl�X�E�zÐ�3����@�1��e�H׶C�
�R�G����]���z��$��rgٱ�n����I��^"���,B������~�R��x�rʲ�'����.���Ѝ�#+����՞,K�A����G
��pԪX�aE����4�mH�w�o�Wݴ"~x�s��Y�Խ3Q�[[�Ve��G2��-^L	��C�i��Th��<ʜ�zl�_��B�[�+�A�������}�i�$���
d�� ���>l>���$��)muj0�lG�������i\
�������%��.�]N�c0��	��S�-(���"������hHj�i�4s��8}Sb�<���R{I�%�&66m�8!Y��������MoJ��a��Y����X�覤�X��n�Cpmu���r�m�]B��=�}.�$�U��!502 a�Z5�R�uf@�L��0*�F�q�����[�$bmqm׬`���ǳlrّWTR�sb&u�,0߀�C�C
�q���}���(��y�G���[حu�X�{3P�qzS��8�O��&$ܰ�Rb��ȗ�p`r��Dȗ!��O�{�#�?[ф��l�ޣ0�s���z:#m����*e��pl�����)ӥ����'f�|BT>�e�7�a}��w�}������ԉ���*�;��N��R rOU7���X�Z�,-�6z����2ބ�-,���̫�jq���7�iR��֦7�����_�D���[3���6���!�73�P02�������|}�u
�!v��c�[1��E����?{2ϻ3S��w~�@�f�8g��*[p
~�?���	�:g�n=����)���xj��,�p� ;�ɳ�����_����MS � -Kq�=7��Ѩ�߫y��vk�
)bl��u��y�����Yh���WL�5]��%"Tp-��7�z���,�m��W��^^�_�	N�PS�*4���U��X��m�FG�95�Ь�̐2�	/
��.0�vZ`le�-�I���y��p\Qυ�2&��0tt�1#1��i�C�(�/��ю�W���J���F�>�"�4�_��L��T����i�f#w�&��ۨ�$[ɪe�;�W�(Skӗ{QP�2�S�?ł��X�]bz�Dn��;�,�L1�~0+��h0��F�/�k��qw�,摫�Jj������P��*���o]F�2�V7ց>3_Nௗ�N��"��g()�*\�>��J�SG0���H�v!I�Eg;�I>DQ�bn�Ji��!Ku���Y�d������j���D�s�@�̡��~Ϝ�/ԭ���B��>��~��U$|�r� f��G6��`����_Z�%9�ے��Z54o�Lc��,��8F����@�ov�kڍ���}�n�7bV�]ˈ��u�I�$�_V.��*�B����/�3��aL�,�c�g�y�[��^U�?��ـ���t����6b�C~Rb\L 2���
��`zc��~p�A>�V��C��W�}1:,M��V���y�=H���B',�Qm&�V�{qWCB9�T�Y3D0����ӈ��ٖ�,�:���S9�hW�J��`�P����;�T�}��6�3<��"���,�s��X����j�*Q$E���6�(�#m��3�f�.>ॅV�>x]�z��>UT�6�c�C��Q�錉"ެ�]�I�CCLVF��"������l|$���C�_W�?dj�.<��t-�:j�g��qde���;�
�ߑRŅ
�h�T 㸓C��ڸ��>�]N5l�S��d�����˲��D�٨[��?H�h�_>���V*H��h��u��p�u9��ˇ:��fT�E����Qh�^�/v���0�H��1��=R&��h̦¨�0���ƿ�0$�/�*�)QUj�}���ivZ$gި�	/��0G9{��3�Ӎ�@�T�Ҕ�������H�F�|g� \��-�kA=xl�kh�<�],�C��6\$O�n��j���!�U� :Z� Nx���ǜ~�Q��^�4GiAJ��h�<��`$����34d��-l@�6~U�+�|�b��Η�7��/s��3�,��;=e��\��@ 0��;���H�8dRh
.��ؚ5�6�Vr�D<�n&E�%OR0E|��o��y(�q�~��d���B�xm��[�,ܤ܎CB"Ȍ��==�����gDo
�"��q��]VqrX�֎y�����Fr�?ڒb�>�[�\��*���WK�~H�Ҙ������^�{�K��px�	��V�5�
�W	CN�YVb���t=S�Ϯ�i�1���F/>�[���	��f/Oh�r��ʈ�������i��oQ�;�x���yi���o��f���L�ypှ�ǊS���[��T���u8���fAp:�����I?vTj5�V���~�T0xM����{�I6TE�me���0v�z#g�I�ʟO�GȻ�R9�Ҭ��Q�Ar��Kť-wF[@��6Q �#CQ�s�"A�a園�ȅ63�z�(�S�u� ��h������7���x#����f�,� p�Ug���7�J+L��TGD7�b˟���N14� �����:�\BQ7���C2��C��c~�����ɯ�V�Z�>�g�X	��A��4J�Am۷����Q���/���A�gӶ �a�On>�A��8������ny�WhT��w8%����IC��D��0�	<��tt�`�<�.���/\WoF���|y̭��t�d��V��]���w!O#<�o�]
4�Iuί��oP&@��l��[|U�=�C�*�z^;�Kժ� �H"m[��l����5����M�o>݇����_��� ����P��c/������Gk�0re&�+?��4�` �զǮ�+��0�ơ������[�Pl�oR�b��i��Y�Z,����Zy��tqE�F2�tvâ ���R!3�@�5^{Vt�4D��^�̭̇s�����6����W�6�k����]c��A��q'F�>��-�K�ul�F��?��C���v�R�J�ίVE�U����Y�/��s�����$@,N����`�O����Ԩ��uG췖Q;�#�SңM
������&��fK��V�=��u���`&;����/��~zSV=%ʊ�=���'E~;���͚(�e��b��~���ћ<�<��Ej����йj�c۲��ݡ/;�g`�����6��ӧ�i�h
�<^pe���$!7�`�ē'��\[3�4����5ۦ�7������[�k]gIL���l��K�v͂O�C#���!^�BN��pAB��s.���ky��y�Jf��������.Eƍ�%'�m�$���7f�}7��^�w((>O>�-�!��Wa�L6"�(���f����%i�D�$W���K��Č�z��L礊�КW�Eˣz��x�P�\%���·}᭝�8%L����~L�6����u�{=�XE���NiႏJJJ; ���7��'�����-d��x�����?��۝K�����]{>TP=oܤ��Qx����q��a�<���|[��?�ӵ��?b93Zx��T�I]��b���뺊�oaL���#2�q�E�ޅP���Ý6-26o�bF
�}�:/&C��\}Uz��3n�P܄�7)�Zt�u�e���Ĩ��]Hw�P��r�����;N'm{�g�2�/�k�Z����L�(<O��(�8�׎�mOX˭���ej3j��]��:r�.������?82X0�^Q��د%���Q+����G���x����c������탊CכUO��Ӯ�gU _i��WV>�F��l��N#V��#�W#��3��X��y*�U�KWi�7�JX����V.��\�j�bj�I��ˑww�PR,���
 ��o�|�w���\�\�E���x#F��q����<g͕��;X�`uQ��^��T��������g�C���nTO3TO��-L7�K߆^q�u����k�����z�G�n???�Ӎ^u::��aн��g�	ɎN^t�>�k�a�҂���'���U����cS#%" ٥/��*�$x�/���2�T=�۪:҉�����L�����zv,؇��:�nV����_�c�����atA�YKF2�4^l���!xN����RK�� ��V��gHA���Z��)�9�^� w�1�\�ы��[;:b�8TTV6��!���*'��eu=��h��ei�?=�1�8�K�������s&���AY�҂���F�N�� �����k_�K�]���˭�{޲�L��c¡�=��	Dzy��b̖-#�RJ0�j��z�:L՚���]:�Z��>�8����0�~�ˍZAp���kIL��D��j4������9V~��/��NWEEE��t���ԩ)ڴ�h��Ԉt�+~�=9y�ofVV��/�a�$��pIf�)�	KNA�ؽ�@�֧��u�����#~�^obC�s����U~���2O:���f�����W����w������[�˭"S{;�'��z2K\�I�z�u�ф�p��I7Fmn�x���_�U��~(����ϕ��*��U;�*�B'��i�i�E�K˱5~�ZD ��(��?�U%W�T��_������d ��gj�P�!N�D0
��&���`!|Qͯ��a���
�k7��'�"�1��!H�2��殓c0��>Iv�]��+Č]Xk]*��ciɇ��h�  0�g~�� ����J���{E�lf@�4�"���� I��4Y��=�V�F}������>5�Р=F��k�P���	Qj�ZC����� u�m:�����4��������˔&�D�q�s����G�{];	,�q��:����Q��C�Z�s��狗�&����h����CF�+���xO�l'��;MN�l��jq��<�W�!��H�Kf��ݥZ&���0qpƧ���S����a�m�;?J :��n9�p!���dj���/K7.�**O�����"F^���%95%�>�ET�t�.|@��v0���F;\�w��P"��tn�v���"Ly���s���.��%���^r�伐D;���5j.~�9���Ͻ�~�j�Ȗ�e��J� ��J�e\D*&��Q�d��-�c�о��B�� ZQ�K�I���
�4�e)�466=����
���� �+��Eժ7�1m����8��j���Pt�= ��>�`�r��e�bgʵ�kO�9�|�_�T+��&D�͟��Ω�[p�W�E,�<�K�37W��8��)ˑ�L#���lK��7�-��h���_�~~��GIôU�L�e�:�>��b��E���6@��=^�dN{]�0��O)?��'��c?�Н ��Iy}��� Иf�D��ԉCDE�7����
%pv��P]�/�X�4=^���?���K���4,�����]2T������TH�y5~���F��B��Ae�O��w+åMX��/���"48�$�E���*V|�F�'#̮Z&z������i�Q�\o5��<(x���.[{�2#��;kb� ��������!�~w��.� ##����>��%
����o)�Aw��)sx�_BL�edZp���>X�K�Z�a�Ί��G��F*))�n0}�f0�#S���fp)����^^��g^���O�?���>����_�7у�dʝ�Gqu���B��G����c�P��d>䄃ůt��Z��)*��n7#�Շ���Ǉ^L�P��/� �k���p3u�3�eK��%T���P&��ju���"�n"}��Z��J�m�IwxG�?����`�jܸ�-���pՀH0�2o�Y J�+ꏟ�S7�����U��ߥ��2}pX����Ϳg�D�N�og�t��3-�0�&�
��7��՚�&<Q������b7���E��>>�/C�	 "Q�	0A� ���������>n���y��v�s�*��QX�\��c�3��w�H6Ġa�병���=�I�����S��@_�<�|�a��D�(_f�I:�!�&���*�d(���ʞ�e���fA� �&��|��Ȳ~������a��/�% ��?>~�[��h�Ώ�Q�FYz<���F1H�؅���������9˥s�9њ>�w���8Z�Y��ϔ��i�(Z7�y�˔1>�w!#�ϛښYFyZ2��� ɔq��}^�8�JR�J�j�u�˺�d5����2]pNc��A�0�����5���>���~q�|�Z�DlJ��͛����\��_M>y�v�x�|e��-5Q��F�wA 8e���F��d��r�?�0[�3 �7/7w��s�Ոs/_�쇜�Cv��Y(b��L�}�l�+H��?F��l��G<�!��ɔ����!����N�.U�xΫ?"ՠ=�W�u9�Z���G�n:y���J�Mf���+��R�"J���(k|�|�Ǎ`$�[���ܴ&���P��sr��5�̽�����6�-q������X˾w������.��:��<TW��r���/w
��}�c9�跩�?�=�4kT/[C�:-N9�Mb�^�:����NS=�̦r2�8�ߴ<\&�a]�~+3?��;.��յp���l�ۨ��G+//'�p�n��U�DG�ǡ�fl?��
 2@t;<�/O?���ގ��/�]/�~�^<��+�*no�=��X���:�ẵ(J1�r�}�-�H<�?₷��WC�ڤ�\ ��ۘ9@.��			ٯ��M��((�s��t�����(sd������ʴ��}�E?� �W[gl7G/��qD���i�f;?Ty�P=V`�PL,,S[�(sD���}�Jo<���$ߞd�a���!�_󾢒��[�+�p'�*|(���ů6��랯�8��y�O����V�6�g����zo��aK�pU�;Ez<@��^FB�^X�������T�u �����~�W��_��R��L�i����L'��'�"����8���It-���$����\^_�Q.m�0&�:�ڢ��l6�w�LoNV�fs��"p����	�y?��|��t>�tDĵy#�� TTF�C�~�=.�X�I������d��k����3 �;�����k��̾�0�y�ҧ��7�ԗ� ������/�;��r�F�Ɂ�f<E=�C<NV��>���[?��AH��ܦ��_T#Yb���q@]	#gq���OC���0�Mg0}.���a����h�L�M�j�]�0�K7g�o��h����;���r�tI���z��[α��q�&�X��2���7���rs�yZ������(����d^���m<��e�V������c4k41��!\o�1c�W�j�m"G��0�g�7��Չ6�9\�m��-��M��Ι��q��Wˁ�4E��hd�	Sa4h|盝��J�a���|�JJ}5?l��5u�����IN�`H�����v���g��1�}l�>g�/�R�K�$V��<���,�VVE���`����ó��G� �O���N�?�N���� �)%�U�m�\�dϟ���q��N�ct����.ׇ��1)py<��l}���ە9��F(����� ���tx/�G]�謍�(V7r��Ϧ��q�u�|͎�{gs��&K�?�1"+�d-}M�f� ��I���J���Z6&}r��y���;Uzϑn�h �����Z��1fc�� t��&!��F�R5FF���9r���H �K$���E�KZ�By=�m>A�[_�MWf#���4�`�����ZZ�-�!�rDZ�᠋���_��n��O,�w�#Fi���Y�G~FٸG�Z��Α�U{�*QW��s����|��0!u|:���9k�O�λ�k>;�8H���C��"���X�ɠr���@��G��UF��H�w�<~����-�{ ?�A�ժ�|�������BD��Ԁ��&��~���G%w�dɮ����tM�^1B�jmz���}�"C���B4^�\KyLIU�$b�͏-Y��?n��DP� �$b�ڢ?���V}�G�"�0Ԙ��i�5�l%-H[y�\�l�+�_/�~q�8nf����;�;"[󳰷������ǂ�+�7���O��S��X EJ7hz�<������	�y��tx�*S�" �*�����|�����N����#��m����a�߆ B�9M�{]�O��s��Ȱ1@�y)�k'�s`� �"ʎ"�9@�R `�h9Ef)��h4�5󶀚qui������0����7'C���l�7/�.%8
w�AV0�>���� {F5�Me�`^���q�$n^��_$3w��^_�|���ֽ�V{0h:��k��׆� G��ȿD�/�]��?���n|'##s��rS ��Un_BG'3���٢�ע���ӻu څ>���ހ�C�fcL` T��L?��ձ�Eő֖ cU���IL��4��m��T	�����4�&��� �VΥ'�����!�R�a�����7���FY�g�7nI��s��ŭu�:��s�Y�,���}�'.4��Q�v4ub��<�`��1�dT;QP-�a�{���i6����Bo*���]�~1F����ޣ�^�Q����|������ӎ���G�U�w�K:�����>�/���EccQ8B��[������r���oxS^��hu�3/77�,�O��J���<d�s�XNo�T�e@U�)��]�h2�t|7
�� "��:�[q��{��b�JU�J��AW�rS�3n%�x%�-�If�В���տ��S�N]���������<H��a"3OLP �mD �Y��9�D|/#-]��"FQ}�T����8���c��^]K��T�t��B�3�Ԫa��V��2OW>O�2���f��ټ?��bܧN|^������V��Ǐ8��	�����>��۝���Y�W�����}����nX����|<xuছ�1K��������O	���t������(�"S(�����QL{�y�L���#�T��ҿ��c<�9U��y�ϱ����re��ds]�P����S�Y��6�m�C���D[�W����u��4�k��i�8i����аg�&�[.B!n�A6�������v0��P��z��^�;�̞��m�]^]� ^�&�ǁ�8���t�qkz�-y6Df#|_��n�;K1�E��&o��WI� �1��dJ��>|-�ENɐc���Q����u���}�iDV��I���礭�;Q%V���x���I����Vv�������c"��2��o��x0{�6^��[�F�7�Bar�T��U����O�AȰO��������~d�b�--����R �Ah�I��@f���z5$b���r��,���E��(�3�HqpcEj"�oxg�T�y�$���UUo���T'��ɳ�PM��j3��d[;�T-�a!S�1�0R=t�"��$j�,��
�ɦf�"Z���\K�@I,��o����[B��%�B23�q�7|��+��������v{e�Є���N��w�h�2<i�e���>�U2��� Deա���s�z-M�g̙#�+~���#�z�1��ԋ������[���B���h���?�U�!�˲)I>�3W!l�pϓ�(5�v,V[�nQk+�o�����Q���>���,"qvd|r��1+R7���W�X3G��X����;���q>5�\Jm5H�R5;�D14&���P�|Z�����&�0�&�v;l�N5(>"`9�`�I��.�NƂ>`�&?��l�7��)a������61�F�ڐ��0��0���-�ii��pr����D�u�	_�泌�3ۘ��z�����
�Dg�5g2�~Go8����&F/��"�����!������#f����OML�],z��/���$(&�CaȂ�*	n����>t�ja��M�Q�e6@-i����`L��|3����y���q�m�8�4H�)c��!j8�F�<m��7�@%7��H�-�`���5ͼm4WH*M:q���!����֕�SH\ƞ8�L�t�7_=8j$����nK�$�0s���,�~;_ޯ�Z�5L  ���;sWmN�?��1x!��>p�H��͟�V3�!$�N��t�]nCk)eh8gnm�z ����l�yҩ{E���@�wb.�8Z�fM�3'�K'���=l�Lߑ��JY��[ϐ��5���*���/�
j��Z^�X�əS���7K� Bl���IDѻ�u�n��
��K�!fg�����?���RM��I����1�e�v��X���ɻ�r=���on�g��渣i�mpX��'̫�"�b!!���RE��o��Y�9�G���U��/c��eo��H�:'���%:�'e9O�!I�����Њ���ѱ �M���'7��h������哎�!AWL�sȴA�T=!��n����!�,�Ud�{%	#��Tz)	)7�h�$�mo�5�f])ႌk*M�_Ҵ�e��e��n\�K,��|I�1C�^�5�y��
�����_�G�uW�+��<�Y[{�.on>!��s>>�ɠV�tQ��g��~�wR�B��*F�?I&�A��6]��F�JC��c��fq�����H���n����r*򫟄ﴠ }��{��}��%z�O�Bߊ���9��7�r�����"���@�#��#+U��)X������G~tB��۾��813}-�D�,����7A��N����U�'}癧�ǽsu��)a?� �������ǽ��^^�����윜�:vcҧ�'U��/���^�ٸ6�#��Zr.ߜ�H�sTBp��f�l� l���+ר��S#���k���:���2���,<_��{X&Ơ᏾�R�$�8�$5&a2Uz[�n!Ǡ�����j^��)� �C�>k�
%�ݾ��Rå�t3H�7F��k��c�íz�^�k�ۏ�Ŝ����m��&�u=ࡾ���T���'B���9��`��VB�7���+ˉU�6@�Q� ���=���7��
o3�Z������n�����X,~\p?hd�rP!1����,�\��eސ�pQn�5%�Wi��4����s�X摨v�_Ւ3iZ*�se��������Z})�~���қ�����S��k�}	b�an�P`���X���rt:�ep	{Yr��X��ͼ�&#��mw����O�f���F�აG�g1p/��,�?~��0?z�Ҍ�\Y�ci��K%c^Ҝ����F�tUNx)�����
*�dz�m��C]�d�ō�Bh�z����`]x�<��������	-�p������m��H}�3D'��X	+}i��d؇K�zɉ���὞I����`��n}��x�۹
���o�u�B�5�~��نb���tI����霻@� Dd�i2��/l�*��L��
Ƣ;aC`0�q�Wa~�j���7X))E�����W��BٿN�Ԙ����XJ�A��ÊjF��{�\�y:h�_��%I������e' S�Kp�6�&{���0���	��SZ8��/PJߕ^��\5�[ڸ@)�>�$K��o��~��(�=4�͢�wYρ�U\ErU-�1-;C�=0j?On��7���c��;���}�ҶY��BAЗy�䆄�����A�]��r���Gf���!��*�Ջ�\���(�.6������Z����[okD7rK4�����WK�AX,O�&��K� �*V��ldO(}�ER����0��½�{Щ���Y+�&z��Un�te�Z;�C����U����PeK�{5�čZЊK�+���܄���y�/Ʒ�,
�
D���C2S�02XHc���R��u��9o�E��:n�k�v_R�h��J䲃5T�3�V'�ͼ����$�ʎ�Yq�>B����A��_SF�)�rV,llӧ�������Q_1H��U4i+���nlҧ��;�#��c��c�
�J�$��^����hE�N�Guh��H����1J1(����u�3{7���WN�;��߄4�0(������vT;^��O"%V�׵�U�SG���tդr]��2W��{gV�;��g��n��*�%��A',P�r�	W|�����&3:]'u�� S��&�=��fz	��6Gon���D�U��:~�t1X8==}�l\:�w�Pl���A���b�	��V��٪�:ez���e�|`v���.�d��%+b�<l�|V�'�廬��d(�9,����v,�s�(�fm�=�Z����O�,=��i"�$��@*Q\'����PI���gMwU����239���O]	�o����U�m��kmU(��ʗ�#�l��$/�{��(�r##R��!���рo���E���K0X$GőѦ1��j��mɔ'��i8�~�����v��� <v}s�P%+�����d�Z�,l���]�Hi��������k��������Fb7�%���[�O�#�Js��*��:�l��b�4�n�eݔ�&)�h�s=/Վk�,�l�r�W<���+u�\%7oh{����L|����UJ�2���9�t��%�������\X�d��V�'ޓ���8�}��섯䋘���D����j�pO�<"��'�_b�� >y�����P��g�s����Ƌz���&�1�\j/Vl}6�|��� �*OdU�K�����^�һ9�^�����L������k���I�2��N�Xb`cJ��W�\�C��SR)��<�:w����M�61��4o��Gއ��p�(������}`7�����qM��r���o	+���U��;\ҟ��׺|\v�S�߬8߬V(�����r"���֒+�'RHx���)�U�	��=����E��l(�I�/��94��Ȑ�NPks]��rdlgg�t�|3�[tR�M�"G��Y��5+5�w��y��_|��,+��h�v3'�&{�]�8��^`��6f7���S��T�f�Iv|�"0?D�B��f��K�\_�DS��,H�U��W�=N�lڅ�>����~��YA>�O8A��z�XA��vC�#���{�*2p�p#C�Ed���������w b�XæF�����ʍ5�B���P�{(�	�K.�#�nX�;��$=�W5���iF�>h�O��	\�(_�nB��[u�c G����iT�*�����?��2����-��;w� E�;�����nŋ;www�Sܽ�w��3�L�%3���9��n6~6F��6�5�͐R��~o�'ǗZxh�,0`��������>�?tl����I�{�v'z^i��-�~*�����5}cegj��w�t��?*���1A�Ű�83�m�'w��I#�ad1a�ы5��5~w��]�߽�a�6I>�s%铃Д$���3�~����2�.Ȭ�jɤ2�;��$�I�6��DA>n>;���Ӵ��vˆ�wIq�����Z�C�>����j�N�����AT�̼��*<�0�`.���6���;>$��q��_P�9�Ȣm��ͭ�7n����\���ש��5��w�+ɚ�	DM��-�i%f�Xq4�W�_>q��%H�������N�6��0z ٯz��|�0]�CȘ~��۞?��c���� �+��)N��'����qY?���s�̲��|8�
��O���F��m���/�������n�N8��P���3�~�nFh2�v2�ʂ/����N�D�+&^��R�|ݖ	<��T�+�n&)�j��:�EM�<ƱH�<�����Z��c�k���T?׭��MX���i��̭g��-���bVLL̝���V�EyE5��G�V[�Θ����eG�mI?7�<p��m/�я?��8���� �>�L� g>�~V�?�����j,0�$Q���b��ᮊ&D�2�ڏ�ܷ|�YZ/ ]���?}���b#�{h��ˑ���N���������"�+�l��?��T"�y(��O\,f1����̈́�:���
aɗ�'�O�Y9-i�fѦ��&K���DCz���"fU�:��f��ܞ�����K;F�ьZ�L�Ҝ�բ�G����@�Yw�s�>�jJ�}+g�[�	����$��B1�|��$�5��7Ǝ|u:�]�j1f�j����y���.m2�)�>Q~�"F�%ݎ�p���OO���͕�lB'&<Tht�^4�oZ�B�_N���M_~r^^$Y(�t�tQ-4��#�<��`���^]N 5�5�}(}�I�E�ՂAt�JN��׊bZ�'v���*4��C����4}
>�xTU`���*��ւQ�PZ�k�V�S[�l�?X͈w���c�����;���10,=�N�2%_�#CYUʘ
�2(��<T���g6��c�R���M�s�0���w����ZUa��if�{�ggg�1x(��6��!I���E��Lģ&'�{Wxudk�UkU�޺��̒W��n��n|5��[6C�zTkc�\����݊m:�:�1w�%��ׄ�p�k)�J-�:��9��m�V��(�֢�'�8�?먛
"��������^��]��=��������ml�'5c-/Ӫk~wI���ԇ%��ƨ(q�'�ᱹ�=��l��O��'�H]HG���o}��V�T���M�.��p+�M}�n�A����W27*���5Uh�X�I/�Wi��=B���B����+d��2F}ʍ�O� .ҬA�f�[T|�]N��ML͋X����+����>����<�t���;�'VzOnK"�q 7�@��(�]��i�A�Π������'K���AN5I�;)�^�7�7���0'W�L����pI�6zO�	} Շ�I�VE}��T�q��w�{�e9)LwA�`u�L�P����б5�1͟H�/������32A)��d_��CW�dd/�OK��-QW���Yq�7O4K�?'�۾���wA�W��L#.����� !�^y����Q�쇸�Z���f�g>Z	�r�(åD�*m��m�Vz@H��a�&Ufj�gc�$�?�c3l7���E�mPK����pޱ10JH��Q���R�C��sΡI/4v�U�Y�@8��z�Ψ�����>v�GD7�9�S�b�V�3����EDt�e�+$��BA6����WJfPw�ŝ�q�79pT� �d�^��V���̖76����Γ��D��H� <axs���""��.h4�M�`� T����ϻV<���4y�YN���t�׋bOJq ��+�p�~M�*V����+�^ӺG#|�uP�ZVVó�70�G��㐦LPvXe!=$��xq/�z)a]=����m��EI?x	��RC�F��C�E؜m������ؼG)x'�v[���$������ɵ���TʘiJ��X��+��d/�l6�t�Ro���ΜWD�T� ��T_;,Bn���v���G��fȍiƮ	����q��b�o(�ڌD�'�v�1�&�8]~UY'sr*�V�ԺU,�wsO�����s+��G����F���֡K#+g= ��8g���X.�/͔0X���v�~%)J���b	�YH�S�D��B�	��L~�V�<�b��0ɟ����]�.L~�A����*R��#�Bq�Ԁ�к�3&�b�P�Ee�0r_�y���������o�"U�j��'#�YF�K:S��:E5�1$��e5����4���͌Q��,��9�����5�&�9��ť���w�	ܖ��D�S|`�[�i�^`���{��ʋ�ZY�բ�"�s~��s�A5��By�ߗ����[2lȠ�MI�K>��9���<���X�D��U|�����J�ƿf����&��*Z.��?W�4�T�!�PEz��n|���ŐG|Vy�@�&}M\	����W�K]	ھ��Y��!��0Ox)����S�d�r��/�KKO�4ag��8FAH�\�I��>=hsu�PK�������|��e�S@��Z����;[%�}�U	ބ<	Jn��0��B	����f�n&�;�vd&FT1oE�e������_i�*���l�-�����l�=�[��ַ���Da3�mfw[�hu��"e@�V�ş������P$��M����ҽ�M)t��ɳ��Q��S���) �h�j?s���ױa�Cx�+�bb�Pv�!2�o��b�4�;SH��(��\ ������W+������8���885�������)/�v�x�����PpcH�1*q�M�Q�*C��JV���1�A�2j ����碉�o�仼5hd+��k豟sc-e�[����~~A�<�Ċ��:]��8��e�%:s�4����+������6d�e�f>E��u��[qk);�pm��x�6
x>-g�4{z�4"�s	���|��(��
a|�f��H0�W�����{�,�� �x;:�ggg)W�����LOO�	��e�r�ГJ~>~I����,�锚�Q(2@��s�"�V�6��z�%[<��9��>N��P�RZrRX���
�L�7���2Lǻ�d�|�*\�?nOY�a�I}ϑ	*K�k��V��ϔ�+�a@(�pY �`�M�d�CN������Y��XY?�s!�߲�2N	SX<��"e\hJ�������b�֨�}�����sX(%c*i�����L�M�i4 IСHOɫ/LL�>@.c��D��!ڸow��e̬&��L����-�ǅ�H��}�e�m�͌#8�?��d���H G��
���	z+$߳�zy�#6K�=���3�v��$vvv��sGYk�����ٞO�4o(Ұi�g;����p�:�l-U�Jb�^����"�(�siBq�%�<
^�n��r�l�N�Z�$�e��t����j���<ȅ�-����.���,�!:\���9����(�o�p���*����ꗚ3����\�$s�/Nu]��d��\/!n��o�/	KW�i@2e��)�x��EmG�x�h8�X/Rh����I̤D��u ~+�O�H��0��t�/��W�4aQk�O����H�5��]��β̠x��3�!�����@�U��^
���Z&��f��I����0_#P���������	tOM繲�~VF�/��H���Ł��V1�T㇅�D�e�>�V��-JԚ���z���T�k֮�8]��͑}e0XS��F�����س��\6�~�Mx�Z%ڤU�N����6ď��T�ē���Rݼ~�q2�C#�:SDh$���l��A���[��ݩ����`�r��3rӠfD:Rq��.8`!�g�r�r5�=&�U�[$c,x��},���L���\�AA$�^�Y�뗑�\�kĊ�?��O��?�vGHfu���<�z�Y�w�>�������D!{w"��3��]�#U��`� c5~�ȁ-d1���܄4�������k���4�{��5�{xn�Fi}KW�G�.�LB�|����O�����>e�	{��MQ�Φ�ҩ����ܘ���'�Ёr����������}K�䜢Ф�_���ЎL�4�hw�`T��S����8FZ4>&^�ɹ�*Q����{8����v��*�*y5
9PX��I�,���L.�]��A�'A�\��B�g|c�0^%s�����S;��F��K���e�"�\�+�D>�Y�&�1؎��ʇ�Wڗ�?��ie��>�M%y���	�������Oeu���h�6��-�X����&ֽ3��|�>��# -��ypԈ��d�������8^��/��駬� bTC5d,���V*؉��{vYr�!T���P��J��x��=�0��Q��h-����R���`ٕ��p��e��'��m�W�=龍|n!a�����wf�N��FyQ�����B�H����#����X�v;��4rL�s���N"�q#4=S ��zj�"WO���ki���3�M?����ܝ��aM��>
'��D�ј���a������X��?�ʒO��Z2��<�D��FiմRs��O��Ef���,�OQ����>�BSE��ס:r�pd*.&p�̲%X0��΅�Ӊ�T��6>��gH�J��y�'����Yb��R�%|������!�;Ӯ�юfûg��%J�H|[�G-"Aِ�0>T0%����Ȱ����8����CAD���w8Oն��=&F�U-�����τ	�?�K��UW�i�>Bg_ۨo�k�a�
qy�;�	b˷���ST��"�fĕ��r-��vN;c�_r�{yB�.�.h����q���d�k+#��R"~9Jǰ;Z58�
���Y����f��ڀ>��&�M������|����,�c���a�9�nWE2��K���$�K�����e)�;���TF���,E��7�v�h	����{q�E���nإv٥�9HUC�vQav~�o��o���5K7�*^����!�W=�����4��#�Z�'���|�(�e�3�,X�5�&��9��p�X�G�;o`��6'�^�O�6if,��4ØOe��i��!|P��s�V?+��
7���B[�v�W��i���<�T�@����>��:!PF��=��i�k�2w��R^����V!���O�VY�s�������.�PL�gEs�h�tw^��ٶg@|ˌN�(��K����dϋ��ǁ���%�W�t������:�._��(Fqs}?w�[g�^H&f�O�[����5��%���%
���ar
�Ŭ ���g�V�3���R��"ٱqp4S �7X"�f鷯��w[��U��|8?A�[������.G]h9��E��7���c��{��^� �X�0 'Q��$���rk��[X$ٿ.�qvx(!�V�~g A]mm�����F����}�m�(C��Ԅ�ѣR�N�X�Nk�C��uB����P��p*���X�@��R��g��"[�-�����>f�B�g3i�-lUKxal�.歝�T����@�7��z��;_�I��Gq�X��S�e,��۷h�^'���,,��#ۦ,VE�_���x�ͮ�F�Bi�������
�'	� %{6�g3�%f'�;�����k�XkC�1T��O T����{==$�%a��F�_�z��]�j��LԦ3Y�	�I�%ʖM�|����޿��W�8���Ic��-K���V��Ϲ����7d4�Q?��fg����z��B�I1p>@���l��r����̖h�����˶��2��3!������w���_�η7�H��kM%�6t	��@"�W��M��Ժ�ʖ����K�n�����
���t�,	�\-}�?��sICW��}��(3�sYo��:����&
�Y5Z)�a1q5��*g�J�,)ٮ㻳dHZYx:��U��xC<Os\�Nv�/[m;P=7|=�����e���w�/�~~9�~3`5psK�����Tf��v"�쩾��!O"��2k��]��(о`��N@�b���������y�#�^���NJc�ؘX��cƒ��R��Kn�9�HhP{{{S���^A���u4��6�W����E��5,]�m��|㾤��dV?+�-��.��/Hz4AJj8�Aᡮ�I�ӯj�P������`]~'��͊d˫����s���֯�,oŖ������I*w���jc(�YߝÜ���j�}jʭ������:`��n^��oR-#�ҁ)h��j=W蹴ç�C��κ�ԇS������<��X;<,:_�c��M��څ����\VT�U�ަ*Td���fU����Rs���.��^z#�2���I7�,�Fs���0�ѩ�u&x��e���@�7=��K�\���PD\M�QYW�މ	9A��/��q=�����|����@�a�06>>�O��	��L	6��5�ft<i4�%+�t�WZJar�D����/�.�Ӏ]��a�x,��R�KR1������dvD9��{�{�b7PK|ފS���<*�&��?%}�+�nys%�2�,�(�a,z .��[���.���-q�T��8�����쁍(�U��#�Dt4���/��-V�6�-�Sf� �R�ת�(�h��yY	I�C̯d͖l[�wߐ�}U@+X ��h	FDF��{7�ws���+���鬝���[o�����?Bg����CG�|kɽgXU�٧o�V��˒���j�����2q�c�.��ոȞ�ē6�~L82 �=������,,�{�C��mr��F)Q�=8i:���@�i�`��N�[��^qBdPN�9�b��Қ��_��.o����<�
s`��t���ʕ�FZ��QY��!��y\m�;Q�!:Ȥ�Z:v����<Wb����~��笋�=n�)2�)����xl<_E��K]tj��YA�H(�V���G)�,�LQA`ˇ��R��í.Ǿ.��*$�]O��0\��*6��ۨ���*{��yif��_�F��Z?�=����B�����)�Ｒ�F��"�h�{D� >�C&�r�]�����%,'�P��f��� VnS+:Ş=ňˬ�}t5�YP������������e�<^���#�h�����+��d�?��M2EF�I��s��C~|�zD�e�"���L���wN��&@f�m`MnLf.7�W,�o���Վ���������F��~b��)%t�*l��'��U�0����0�Vt[���ew1����%J���M�0:]�}g����7Eab��hƙ�J4sN�QL:S��ʔ���}�����;���F����r�'�~g,:�5����"�V�1I�q��)�kң��Hǈ�@,����T�9���I��e2������rǽJf�X{Y� �h|'Y<`z&	EB���.ϿE#<��y{G`��M;�e�����}u$=����^�ނ�����Hk�/Ɖ��Y��f\(-�)�HB��hvw_��عU���<�ؤV ttps�n����z��s�8���ƭ�D�l���nuuӫ��'+U�C��V�D�ПN$UjQ�77��|[Q��l���2�y/3�8{�zz�¢^�g�j��a>����4��F4- ��W�6iU]�E�Zw�6���i�A�<��KI�ڰ7`.�PE�Y*jiI4����� R�A����sv8��w��$����pc���NoY����%�)�w@��Cȳ*��S��;��4�9*٦�w���a�� �296���l�����/���g�E4<(C����}^�V>����M?H$��/���]�gx��zV�z{�np��[N,��-ZNMV����L/���2{��X�����o����z�ۚZ��/9���W琧�X����sE3Je��$Hr��:2j��Va� Vt���z�'-6�R�F}� `S~� W�5�0������c�g��s���r�~tq�F���8��X�e�>���b5���]�PNY�I����F��NO����|�����#����X��`G�����p|z��g�P��O��K��,�,��+�~8�����+��ΝoW��.�x��JԮ����$rp$R�ZU��:QCO���&3�8O�b���*��m2��<qpy]��,��!�l˙�LCC����t	�%�����Vy�ݟ弌LL���?��G��	��wh<��G�qYu�!1�"K�7 �7����9(η�,*Q ܰR8c�f�l�
��_����8A�v�,Vtl�Ř��d�a��Y�o)Ɖ#Io������ 
�zd�oT@Ѯ�@֛T��ʜ!R�>V[�q28c���}�T��@��'�?�j�ff�H��K�^��'Uj�4�UUeLȎc8���t��~�3�h��'����B���0���g'i�R�oJiӌ͔T�T�	�X��(ƕ����Y��6-G��*2���-�h;2�#����.��&!�2�^\���=��{�����j�	3�HSn���<7�%�:�uZ��ύ�P��B{oDC�Y[Z�:8�vZ'\yU�9	&��de�� ������ʜ�Vd�`F�ci,#M�(-e×�#l3Ŕ~l�I�&���G�}G�gJ3�˭�Xg��]=d�v�ғ�e�T��tT�!�ML+3�B�"�`F��v�Uwqi�fz;Fo�*3;[\fԄ���-vEq����-ަE4w�_;��L�� �sbr�HVx�io%q&d��By���a 7��|`4�A�VO� =;�<U]7ܯG�]�SjkcC���T�b6�b���E �v�-�;ᚺ����,����($��-��,=��
����-k��,]�CQ��Mkm~5⢴��*�����p�i�A�s%�q �����$����;R�i��E�Y�VS$x60)n���d�`�;��{s}��{?=*��b
]>|$�8m���l/��-}��x��W��wl�/..��Y���D��#�U=�gi��Y�`��,��}��o�xa������`#G����:\��gd)�*���.��*.I5PG���7s�GV��G����� }!�)uL�����;�U����H����X}���Ł��=^����Bne����������9�u�uLB:6�ē��
�B�[���&|6���Z�6׈��R�P]��w�֩�]�%9O��~���4�g�j��®%����BSs( �~�*+x�Wed��s�֕�!�5�	@+W�t#D��?�͇n�=�{]!�����ߥ�B��B7�/B�Q�B6���'Ζ��x�d��H͖�ײ� �8U<Z*k�p�z�_ �.�Įl�|R���7X��m.w�4��8L�m�����nt��ݑ�ib�AIA�%
{qa�jjjx(�|nѩ�O0)�u���1�@�ؽÛ�
ܧ�D�@��P�?��|0m~P�y��;>;���H�4�����>DQ��޶>�I޷�^�1����]�r�������_��ƀOT�n�f� �*P�"��Xm��a��PQ|FڐrnW�����͋ڏW��#��읺Op�������_+���{�k;E�)�N�s�<��f��"�<&�sd�,Hk�<vO/T��$�(�򠜞�����y��2H�ea40�]7��	�r�)"�����"C����?̐�oI"��H��X����N�kQ����,o||\�B�\s��O{�Mv���u���4<�����GՂI��������K��Q8��[z ����B� ��7��׷-����s[�ic33j�20�8�w�w��Xq{��L��<c`pޒ�3�1�0@>��{��=W�����0ͦ/���߶.������o��E���z���<S�,�h9�8n�n�n2��c�O�+q�[��R�Z�B�S�9�BQ�v���T��e�.Ԝ�?O��z�#��F�^7�u`k���Z���U7����j�����,�!=;{�N��gz�nGeކ]}#`��:5b�Hljkc������5��|j���z��cy��(<ׯͽ*�������_��`����z�G����.�F����șs'��'Z�n�KͰcE�'H�W7tv��>��x]�0#��*~L(*P'�O}����v�%��Cb�����1v���`���j�+#��Q�~��&<�t��*�G�V�� S������Bܦt���Y�܃P��,Y�My��@��ŭL��@`���9��fۃ���^X?1� M���	�b�aqc92�߿��O�o`��QcCO��0���>�����-����R��h���������'&��>����\*��B������ǲ�o�o�F�����H�1=��MG���Y����A^]�{t�c���7���S�䊝������/��ۜ���Z�W�y��w��E�N���x�e�ic!EG�!����vz���/�Hk�AW�m�=E"\�P�����q�D��]�������?=�_/�\��a#|8V{]�ߧ�/����)�z�%��F��v��E�g���9sq'�縹�o���_�������9uey���9�2���qin:W���0�I���ˈ�ʩ! ZX�g�_����pY�� `bݪ���n�����}k�S4�8��5�6�C�X�ؼ�t�� ȐT��:���{�9#��T�9����Y�(5�)�]T�$��	����a������9XǨf��/o��'�����p�����)��"�����ҳ��xM�K8;?G"��!����Ifq�9��B"(�4�����WbD(z��P�`����%L��m�l��P�Y�S����f���`��[!o����$�{.@髻���`=;��� �VEk��vF�Ix�u�(����\[䌅X�M$y�N�u��S����z��嗶3/<��eHbX�\��U}�;]����Vw���Q9�454L|}���S)c�&��[���m2����;�ӛ��j�ܭ.�|:=�17�Ij)+]�X��y2������:f�-�F�.�5Tl�$�/� d#�aT��a���n��>��Q<z��"��S����KTD1����x;p��q�X���`�}�Ǯd��1F��/����3
!#I �/s�X?:��K��l�"����]�|��n_����+ǭ�B���d*"�]u:
�ֶ{q����4�����,�9�u�XŇ�II'��D�K����	����=�u^M;�g�\ߒ�r����=N�N;�7�;��V�^ɲ��J{J����`��'�||GǙ�j���J]�l|V�bKQb�r����`A/oI/��u��9Wh\�}�cĠ4)�j��C8W�Fo,-l����^}����u������y6�\�ް;�_p'2W��o���R��3��F�2���S�Ý.���l`j�u��O�����a��N�9�����?�P�P�6�0l�1���1X��>�?0k��2Ŗ-��,e���0U�U�hi�n=]�ۤ8�ʚIcK�֖�A�p/w�J�A��y�m��c�>���@�$׾Lābɿ��;�*�*���HH���_�/�jz�s���{�6/p�}�5����GkÍ3���t�N��F{��>Htۜ��@q/�������[�^?���<]��vݠ�c67cYO�F�T�z�-�0�L��%��:CP?�r����,��U5�������sm�s�"���B�����@>c��v0l<�H�,�nU%�Q�m�CXN;Tf"/���a��U�2�(�KFU�]C�bL��v%0L�i�|�+�
m6<^�]��4=g��u�j�D�����7���*hOM�\���-IlͲn`g8���r��p�@(�8��s����<�*[>��/,�S��䘅�{�����=�E�=-	x�}�������(�,�U	�by�g�%�b憡��Щ��
$]�1Ԡ�����rI^�@BO���#,�o�qY_ �:��]1�%���}��V]���/��1h�D�h ���92\�g\#����ttb�"Uす�gUL2S�>�`���44*�>�k>hˀ@�_*�3˙?�����Y�U���׶��..P0�("���:�^�eY� �d/J8��G�Yn�W"OOO7����?�m~�#y&���e`-Yl��"�e�J�@0%ˆ륖
^}�y�W��L������������3���������\���ja��-�V����p#I�T�t��'���G���~�W������8��e��K�O!��}2Q$��y
ټC�f��Qv-QhAmm_WϹ ~����l���xB���PY�U�����!_-K�M���O��b_��P���.b���C�\�zJ��{<Q�4,��×*�j�rwr��lk5I���l�&���hn^�T!� E�%kh �?`;�9���1H��*'(L,-#&�u�.%��)婒eB����^�5;�b=������:f��++�h6u���bq��u��q�x]�����s�wGw^����{�lC����T��Gqa:>o�~I [���[���p�6���%4�+$���=va���:s���!���"!h��m,�@�8�'?���N��z\��b�m�#O�O��;#�D�� �%� ^a�`"X�z�Ћx삳����7O�����:�B���_c;ÔQ���k��٬b{w�%����NCj����g�Xi��>����a�;�̡!qh���^���'w� �C>s��h�Y���`Y�ܳ��eE����))�x�ϐ��t��Ƭ�]��a�.�B��ߍoX��;I#����������&Iҡ��қ�.�։��j�*���S�g�Vo�Aw��Cx�Dx��Q�=�ŒZ��9�z�O���}�f����ܩ�tu*�x(ԎY	2�����!�"�pa,1�39:��
�v��͍��D!�B�������$��Ѝ����ښ�
�Eb��d������$Yф%1����@	��:]a�u���5��Yiv���3�6E$/�b��/3#�kK(o'+�)[�Y�#s�1qu�/r�D���]���dFw�s�m��Eۮ�(�(
�gͥ[����c�u����nF�bҐ��F̥�Ʒe�o2��"Z"�e�.�58�֛�LN ���њ9{�o�"?Sҥ�9ت*����åk��$���s㡤k�n��5�h�~`�4�E�'��΂�N\�C�7}��e۰2�j;/d�Mu��[��ѩ����C��a��l&<�o�nq8�Q��R��rm�x:{4T�8�.�w�u·,>#������O�sg��|�|��6{S�z���W!�̨��QH[�N��ZЮY��9%�/�}c��N��\��eL	q��ڤ��sL��/F%7&�9�#U����s�0�Kp���<��~��c}�7߻J{z�ș�0&��>�пg���P�M%o	\��_�a)�Q^Z�[�xt��`��9�+���y�j冟~FW��T��������Č^g�Yx �`OV�BVT����|� �Qc1�j�2E.G�ڽ�D�ݑ�eW+C=�u`�7OlYJ���m�\"y� �\�qOOZ�Zy4���X�V���q.��������&'J��bݥ�˝�r�$�H��a���W�h�q����}�5Ѫ;5��D`v�-�(�9S�,ҋD����8md���94a:cL5k�v#hr���	�lY�(z����$�X��zJ�}kl�mY۱FgQrRxC'�i�j�}�k�7�#1}X�-k[���$����S?����8m�c�P쳖�/�rE�hE�z0�`Qΐe�T �jq��bbu����S�pn1�y��es����ï���,��6��l�4�u�±޹<���k�	�<�"��(�8������7s ������(���,�B:�Z�V��8��ā;��/
g]�\�	�=�Z�nT���9ު��3��2E��XQ����
S]���ܨ�sP=���`�2�����Fw�!�h�6�Ro�su��4 +��cw�V��WWG��:Gc�ː�t ���˛��	���?2�n��k�ٶy$�g.����^B�F�T,�I ���6�����+Q ��G��(���odn%�Ⱥw;&�c�S�����˥�!�wq߲�t@V2���-�9�h�3���3��`nY�g�wy����m��$]��wN��X�b�_���/�-1p5�#3�8��mw�PӒ?%ٿڍ�!V$�,)��iAͩ�FW���X��	��g���r�(�"1�tvO�4�N�sH��Z�2&�bY�Ml�\p��8�A�w�>�o� *�I�"�8�_M�#������&<�����>S&�4��'������ݹ\^dbno%�!h����� 7�#]�W�L��a��P�pH��0��\�d�m[_'���Z����i�ZH�[91""�O��B' ��gA��O�=���Z�/�L�t�q�xH�������E+��j[%:��gn=�(�Z�T�Um*��:z�p��8�cpH�m�ĀY���/ұq!|]�n�T�u:c�~�(�4��1I��{�o�b"f^=�lEbH�U�7�����"�nk� �tj,P�W�x�+�������D�(U�
i���9x�q_&=&�U���j��+�p��ɅM�i��!��LW�Ѡ�N��])���f�e�@�7�І!Idp_�L'
���1�W^o��Yy��e�m���?��>j����ESR�$����Exu�,�pf���^X321]-�t'0�|��!�q̝W��9o#X���g��w�NNƖ�S�s�s����_��E��4�+�� � F��8YU�ZSS�b��Udʟ�!p'�	��B���jtk�liפ�3Y�a)��Q�ȑ���)���l�P�e#�s|1ݥv�|(���pd˭��C�ף4e)c�����jz�������ݽ��{	���2[?	����)rw��ާ ��q�%�.�ŞcCگ��R�z5�Uj��#S�u��΁Uj�MZ�#R�������\�ǡ)OO�!@G�eu^6����P>.�"��
-����R^��_��* ��h�v&��N�3�r���ڍ����{�C��^�<�k���p���2ؕ��~D4I{J�� )��aL�V�}'G���#���O�05��6����c���Q�ϙx{g�U��ࠚ[Z�� D�K�I\-Z�_�Ga���
)��"8��.\w�{"5���!R��_�6����ҭw=�N:�'=8�F���}�����\����'������	������s��D�P�SR*XQ"K�;����.�+�y�T������E�UO}����[�����[�[�O�?�
�M���d�R� T	y�+�8�j6�-�^��j�CT�H(7�������Po\��f>��[of�GBL��Mră7�.��sR�u=Wi���	�K'�Q���C�%��Yh�����,��w('���~���r���EɧO����(32�V�
]o�J6��{� ��Um�����?f���]���nұ!vTSB���P�^���s\�����}�p�"�>ܾ���m����@�g��>��P_����=V�'w�M���7���lK�X�ؙ��J?�f5��.�m�2n`�͐r���89���DK�պN�ء����~{�BOe���k���u�9d��cn��%�㖍g[�9��49�ȿKK񃻻�QQQ廤�=5~�C}��Y!Rr�h���3V�[��͎k���${^݀�Rp����([52Q�j���?T-X[��w�,�"��=���dEZ\\���0��K�i1�����I���>�Wۢ����0U�D�j3!�3�>e�l<�B%W�v�~	�D\>��ַ��Z�JϪk�@Ғ[G�i{��⒝���ԖG�Z����W��(7QK‾q�
�ȡW�.=k����QN��ƞ�Ƿ2��g&1�w�ѯX� ��:O�w
���	qފ
x�l�
Ƞz���^d�;�U��r��R�{���Ln���};����tz�j��wf3=w9}� [:;'655eEc��gffBD"�@���8�(�Ѹ\64�UЋ��ަn��u��_8_4觋�=�;�C� $HL+&P�{�KJ������6�,t���}%�#a#��\��i��@�G�����U�5��V�;���'�/��1�F��O���0~�u�]�-@�!C��M�A��=7�AUĎ���&$���H�DH��%��EJu�'E���hm��� b��n��\g�r!��2B�6��b�J%�H�X%�X�Y/iUlE1I����(�qm�A�O�\�3�b4��nUpݔ�GzؖK����� b�2 z�i����^�i�$QJ�.A�R�*��Lc���qf�[�F�j�Q�TH�A�n�U�c�C����	���)�0��P`:u���t�v	i����b�R�E�Ӓf����}X�����4�X�*JlW�.�0-��d�_d}}����#�x�	}�Qj��-g��%��o�[���C����2t��^-ځ�ǃ�-��D��4M\�ʄ	�]�ڨPkT�T���Iӈ��1�� {_��:��"M�:��R������v��=3�b4��	���rU�@��#��h��y��@;Ƕm�l��q1	T*ayyY�.ʀ��OS\ۄ�v���'
#�E�eI�0���׫���T*Ah��s�q0��!���:����B}�h�PVȃ�����l�a`����^����ԛ�\�pnFQ?����o��?����q��M;sĉ$#l�D�*ި�.j5����dr���o|���2á��Yaw�F�R�Zj`U��kgwHeH�^%
�*��j���ʏR^� ����T*�!X*[�u���������n �R)���O���[���`yyY	(���.+++DQDw�W�7)%�dk�:�e�x'1�SƮ9XV��q��0���E�\�U�LS����U$�{��#�u��Ϲ諸U�o��G�D�E�E���3�ʱ�1��$���$�^ل&�&�"@6Y8�d0�ăh�I&�c�2,�{L�"m��~UU��>O�ۗ4�T]�
� |4ϭ��s����}F֓�#Z->�+��e�֤���zY��EI��k�Z�^��0�p]�;w�G?�	��/}�K�~�"wn�&�)�i�c�ʏ�7=B�R�0(�H�L#k�?B&�c	���7�Z	��m֏��?�c,L��0A�HbI��yP�F��D�S��K鯞8A�QG�U�ya�4}�q.��aN�(��u�I�w�!�t����ȉ�8�J�G���p���40=H5A���[�6#)�	�j�1�ZI���z]ͤ2��޻Gݟ��H�n"�4U�2ɖnt/F)RJD����f*���x<ƭV�Tk���U.5�ط�!��O��.}�W?����q��]�F*��G`�T*�Iİ��^�id��\?WG!�n��O�������'>�������m���$XB>�U��	`96q�0�#66_�0>��#����kTj5Z��X�	P��.&�_������&.\��T�	'gΜ����� �kд1�uj����]\���5^z�%�߿��%�vU���l6����������ɣ�>*���0�a�!V���;C)C��+�A
��x����/�������	���p���u��Y�k �m�L%�h�1��0O���((�I�`}�{�GKV��y�3�4��#N�<�L-�j5���}~%���eBO�-􆋬�B@G����r��I����nﳶ����"��V^w�m[	Ogan11W���J�QC��2T����&v�S]~�g/�η��J�?%'��B2hu	{�c��wh��sok���e�c�� ���6�qH���N�����9���Z��NP�I3
���F˶��gϞe4�7�8?u�~]MRk�����P��y��wI��Sm#!��1
�DA��)�s'wn�18�2F׭�oY,/���ɂ����AL
� L�D���2Q�k?f��o1d��8��WU����*�7_ckg�ᨏ_�9~�87o��kIE�0}b��a��eZD���BR$/��"պ�aܼy��/�b�)�x�iC旚[��؂PJ���?��?�Fw�E}q1��JS���}��a� �a<�a�ק<<%�[���1���M���>�0J�Z��ܺu��}���0vk	�2��lp��\�r�o����B��;ɘ4M�Pi�����2���S�c�;V�IV�W�� R*��f�cǎ����o����eww����4�ƃ���vH#�(ngo�V�E��֔��:=V��4M� ȣ;=���\�É9!�c#b���_�9�u�V��a����2��I�6�iX�Q̉��p �6���t��F��82�	v���ؘ�E�WM�K�����gz��Q���̻ex!)�L0=��8h��dt�8Qw%��!z5�{w�x�w�8w��u�kN�P����y�p�{׮���!��2�0D&	�e���`��J1
9���� �˰iz>{w��̨�	�шz}� �#N?����.B*
�h4�G���cG�qC�a��!v�F�v��k��`���O���2Mj5���}<����$�%/.����-�����V�E�9�p<���3�;-^|���9�����C��0BP�}���XXX��HI!�j[T���R�$������Ǹw��/���w9~�,����I���p��9��ܾs��AhJ�~ �6��v�� ���H1<�B	��TeA
HD69]�}�fD� �b,�����W���A�94��*X��Ƶd�V�0��Fܹs��8�>��I��4�sz�Ƈ�oߧV���UfZ�R�!�l���Kc��G7>���$���l�ߺO(G���,L��a�)�r�������GW����]���uKU�ۭ��q�zD��iS��Y=��ضK�a2��K������������v�o��t9��
g_}����g+�z=�D��秋��&RT=�,�$�0T�F�������4���9d0���+�� &��D��	�_���[,--������I��n��1 ��K��,��F�US�!�>�i����:[�c���K���a���UH�'��,�y�j��e�� ���_�3�}H��� �0�"bէ+@�b`H�Ȕ�D!�4b�s���2?��x&���&�%	��1̔4U����/h�]n߹A��2�p�����$2&��B�����1�G�������.�N�I��ģ�������txU�URo���wh��BQ=�]����4���w�JBFq����I�ʢ�:�,�J�cm�8?��2Y�ۘ{�昛���'q�):`�)],�Cn��(���XY�N��ad�Wf���Tƪ�t��F�.����m3GHT�EA0���f����z������j��=��m`��,4�$��4I��$���H�È$N1��t8y�,���"���[�ܡ}0��X^�(6�1�tq�
�b���G]�$ �F��T��>�h4bgo)^9�*����%��N�K%$�Ķ�<l�!�$!����7	�1�q�51��Li�����dnn�n����6RʼH�����y9(�1a4D	�a�Ѩ�0b���[��s�c�YB�D�iILK�7n��f���-��:��~���$ID�D�1$���k�쑪�I�5���|R��xj�
X��EE=T���j�
�_�%<� RSҬU�l�A�mJ\��6!�c��׳�*��K��v��yY.����Q`�:s|�w�k�^f��݃��P`ul�Ǳ�Xf��iT�z��5�2����D%�eR�UU�!�ٕ�벾���ٗY\^�Дǜ�!����\u��J�e4��u{�j5�{�.��ַ�F�͸B ����8�1�(P�L�ƶܼ`x��/�T]N��b�)q2fo�>�/�´���R�T��eY�|�q�`����p�K?���:T�l��2��EF7�lLS��	Q��:MS�ՠ(#Q�K�$���01-A'��,�[3����<**��:�T󾑒�RI�][t����矪� �ǲ��Yẖ�����0"�b�PҘ[B
��p��۩0����`��L�ڜ���a����q�iݧ�8�A8HeB��!�z}u�۶M��Y�'���n�ĊG3X]=�������ͫխV������9??�A��@ɣ�贈a�:��`6F�7�礔�Z-�x�HF��׿2��pH�����ܼy�S��8P|�̉ͯ�ܕ�ٵ�<�����5��2U�XH�8�ÀJ�J���v,�z��(�NZv�T-<�i
Q4"�TVP�{�4lR�湕�|i��B���Klݾ����9�c�峸F��[}l���m�!�2?�Z������>O�V'�$����%G���s�4�sj�H1����{�߻����4j>�c2�P��g��kS��H���TB�|N���1++6+++�޿��8��ѣGsy�;w��.+++�;w�q�
U�6ۖK�L,K2���-s�����t:��y� �s�������n��ƧO]��u�~oĹ��z�a�H��:nN��l[}�˗/�^W�{}nݺ����HŘ�*V��ނ8���k9yZ��:�f�X3��X���F���͛ԫ1/\��n������S~����&�pY\XQ�f���쯔�P���z$���>���5VWW9v�����4}��6�v;�^����
���[ �Y�e�Z�R�Jƣ�h(f���D��&Q����N���S�n�z��F�dIν�]�����v�
A(���x������aܦ��c�����>��D��~�j�Ā�Ԛ��~������f4R�`0ȧ�i#y؀�X��:�Mm�L,JPmԱ��u�$I�����3�>��~�ߔ�����,/]�$/_�,/^�(�(�:��>�}�������[��ߺ,��w�ȗ_{]�˷ORNl�k׾��s��/|��W����߻��z����oO�3=.� �j������<	^{�?j4���������;�v��Y}��B�[�7����"��Z��'������t9�14EG��U�xAzk6ڤ��3��Y�O��6��!�Φ��bW����IF=.tw@�Z��ޫg�O7n�CWpA�0��hFГB���*	�XtΦ�N�1��Cu��8.�`4�L�rt����?K���9-�i�)� ��/Ӈ�\�"?��ʳ��u�u�i��<�@��|�~|Ys�'��5����܇�vv��L�T�6I<y�X�h4Ĕ)�2cF!�����c��2�L�p�ö��5Mϓ<���3�?I7ߓB��گ�$݅O}�i��+iB�WB���F�C����_��ѓF�����ӂ�y�'���:oQ���Mjp��U���d�b��`�w���+���(s=����"s�(vk�y�>.f�`,��F����5-B��M�T4�	C���tiL�=t]G'�tޢ,xރ�f��`�t�g13-�i��Ρξ�Y�z��2PJfY3�����,0����nPj��0m&�noH�H�p�d%�dE	�Wͅ��3m0:��=�A���:�C��&Cj�Z.SV�:�h]�g��vzu�5�_Z�h-��0J���Plڟ��	�qNd�|�2�� ���J�d0��<&��.���3m0Z�R��U=ֈ�z���U�?�ӧOO|�(��̴��n<}E��Sh�kOw ���o��Ǆ�uc�4�03���nY6f��W���M]�Ų,�޽K0����z�k��;-����Lk�l�n���{/��8I��\qt�N�q��Fy߰���}�����!�b�0±l<�x�^�4A0������Z�D��uϗO�.�tv���t���u<K��	S��)e����_�%e�Q�r�3m0�J�P��8U�$�om4zz�$�O��h��`&�z�^�����VY�i���1ד�'M��G�>z��iF��$�j]u]���ݯ�փ\�xTO�i��a��O<7�	A-+�/h�j�}�a�M�,�+�̴�茫�*�C�ȅ�ҒjZ�p1�>���6�l���~��َI�q\�$I҈2*I��*91%O6-��'yB���Q�y�s��he\��|ӆ�7��Tٲ�z���T�CZ,uLf�`tۇ*z�vQ��LL�3�Sa\��|x�DYT�� �i�LGI �j� �0�J/h�E'��q����J~��	�Cв����E�0�8cjҘ��G��?a��>�a����wp���ӥ��Q�!�3}�h����=�Q�$���B�R��Wq]�4��a�ӂ�6-������u�Hk=��6~Mݘ�|�L(�W;�e7�۶��6�b�g�x8���`&�^����j��Xf�,�7��O��&��Sa�(�L[�z�f<s���|tr��I�tY�ƓEc�Ʋ�\��i�B�ϭ�8e��E����3m0��q�����=_d��碈��է���h�vL�x�������L'���T�yQ�l8����H5����N|}���OZ�L��>j��m�Ξ�SD,˿(J�=�a&�ZM���ɢ�#�25t�u�i����I� �^����2�h��8��L�4(t>7�	a8�Uc����� yBM����Q<jd��L��ԽBOÇ�b�_���)NK�&c�78=u{i��#���&���OSY f�`t-GJ���j���H����2	�3m0�b�ia�-֏�c%�����ۍ�m�p��ɈJ�"�4������������Y����+˼x�%���Q�k�A�Z����f���n{�k���s��ܱ�<�k�{��<	f������5N��N�&��8^�z���_=}�4������������f)kmllP��B��/|�Ry̜�H)���R޾}[�axOX&�mq��}�%ʕ���u��666�p��i��o"��:�u�A.�����7���JS�x\�ԕ4�|�0�Vw���2��VJY.BGb[[[�qL��accୌ#3����H����}��$�ˉafN)�Y���E��u����V��S��8{��gΐ�db�]JyU�2Ǖ+W���G���\�t��p���oI)e�2�cY�'~)��R&��������ŋ'�q>5��W�نJ��y    IEND�B`�PK   T�(Uo�rjL  0     jsons/user_defined.json��]o�6����k����a�:�5�fg���A%B];��A���#g��Ѫ(�˕cK�!��|������O������,|Ym}1�M�����m��8�f��K�ӫ?>~��u�����N˲�'��ۻfO��i�ow�#];���'���ͦUAw�TerL�,QP�$Өad�k�g�;�i��֫�>���������1���K�Gʳ��-�w_m��r7��8�>,���&}��64ϩa��,]u�i�{h�i�<+<?�ö��@#�.�uSW$OO��`��ځ^W��c �L0\i��ڿ��w����<�M����M�iv^y�z��t��B�w���:K���\����mgT����^/�Oq��CU���������� ��@Lڑ��+brB���}��-h%�LN��䉓�L,���(5���2�Q�%�2�����k��0��0��P��͡ �I^�ah��=�����~��3ù����+��áiv����8l|�y)�R���"QҖ�&��s��z��0��G��V�8#�N�4J�p(�L#pR�и�n��f��F�0T�" �W1r���|�+
C�,���,,TNnlE�RcbJ'3��N��2B>�Jǌ�Ɯ�R2��P��`F�ƙ��9�M�2_c�H�t �_@�Q`�_0�.�2vC,_iY�fr]m���˛�C��M~�=�*?y�������^^��\	"K
^���i��d≕9�Rgh�^c�cx5L;Z��[��B_�a�$U+��,�:'3�1��L*33(.�{8@��-\ra�(������jQ1)�#W��dҀ�ݏ<V\�Pi���[F	�7Cu������ %�?t��:� �;�Qw�q��F�}��.����Zp���uw3��X�r��'����pfg�h��?���Ew��i���t4��j���a�
tLktH���a=�ɷ��ƕF2%щ���a�*-�0z��=�K?�]-St������G���{r���a۞�~��[	�ƌ���i��0S������8��y3N���$AOpFx����n%��i[���z�]!lWr|�8�c+t���J~�j��@Ι���D 5~u��J	FYۚ�'34�G��0ݯ^.��\������y� �2Q�с��S:U��d�(yjG�����N�e���]p����W D	��f�(�)U�a�[G��c�f�"
I_����/�E�j}3䕜v�к�	 (3b�m�Ps
� m:֒%�>�Y����V�ʝl+�G�`���V�����x\eh��>�Yϻ�8tB��!���z�^C�q�2Th�e������Z�~n:������PK   T�(Uf��8s:  D            ��    cirkitFile.jsonPK   T�(U��c#��. ��. /           ���:  images/46b9f12b-d0df-46aa-ac71-73c8a35b8753.pngPK   T�(Us�7+5J  dK  /           ��s�. images/6c71542d-16cb-4630-930f-71c4de5e1144.pngPK   T�(U��4�� ̻ /           ���/ images/7a4be1c8-201b-41f2-b584-263fc50cb409.pngPK   T�(U]�!��	 &	 /           ��+�1 images/98931e0d-18f3-449f-8fca-8d5f6b2df0a7.pngPK   T�(U��K� 	� /           ��W�: images/cd1eebff-8d4c-4172-8358-6f93b12ef793.pngPK   T�(U��!�D�  Ԟ  /           ���~> images/cf2dd1a8-295d-437f-92b8-7fcc138ae9be.pngPK   T�(Uo�rjL  0             ���? jsons/user_defined.jsonPK      �  #?   